* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv vccd vssd vdda1 vssa1 vdda2 vssa2 mprj2_vdd_logic1 mprj_vdd_logic1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1_uq1 vccd2_uq0 vdda1_uq0 vdda2_uq0 vssd vssd2_uq0
+ vssa1_uq0 vssa2_uq0 vssd1_uq1
XFILLER_3_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1828_A mprj_logic1\[359\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1902 net1903 vssd vssd vccd vccd net1902 sky130_fd_sc_hd__buf_6
XFILLER_41_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1913 net1914 vssd vssd vccd vccd net1913 sky130_fd_sc_hd__buf_6
XFILLER_28_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1666 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1924 mprj_logic1\[314\] vssd vssd vccd vccd net1924 sky130_fd_sc_hd__buf_6
Xwire1935 net1936 vssd vssd vccd vccd net1935 sky130_fd_sc_hd__buf_6
XFILLER_3_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1946 net1947 vssd vssd vccd vccd net1946 sky130_fd_sc_hd__buf_6
XTAP_3202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1957 net1958 vssd vssd vccd vccd net1957 sky130_fd_sc_hd__buf_6
XFILLER_19_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1968 mprj_logic1\[297\] vssd vssd vccd vccd net1968 sky130_fd_sc_hd__buf_6
XFILLER_41_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1979 net1980 vssd vssd vccd vccd net1979 sky130_fd_sc_hd__buf_6
XTAP_3235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input127_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2044_A mprj_logic1\[214\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_202 net1865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_501_ net332 net2057 vssd vssd vccd vccd net791 sky130_fd_sc_hd__and2_4
XTAP_2512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_213 net2071 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_224 mprj_logic1\[284\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 net1459 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 net2002 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_432_ net1554 net2198 net91 vssd vssd vccd vccd net550 sky130_fd_sc_hd__and3b_4
XFILLER_26_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_257 mprj_logic1\[78\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ net1702 net1365 vssd vssd vccd vccd net931 sky130_fd_sc_hd__and2_2
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input92_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_294_ net1720 net453 vssd vssd vccd vccd wb_in_enable sky130_fd_sc_hd__and2_4
XFILLER_48_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[8\]
+ sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output513_A net1143 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1144_A net502 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1409_A net1410 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] la_data_in_enable\[25\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[25\] sky130_fd_sc_hd__nand2_4
XFILLER_53_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1680_A net1681 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1778_A net1779 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__304__A net1634 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1945_A net1946 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput467 net1063 vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__buf_8
Xoutput478 net478 vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__buf_8
XFILLER_42_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput489 net489 vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__buf_8
XFILLER_9_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1209 net1210 vssd vssd vccd vccd net1209 sky130_fd_sc_hd__buf_6
XFILLER_0_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__A_N net1585 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__214__A mprj_logic1\[381\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2161_A mprj_logic1\[158\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input244_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1710 mprj_logic1\[63\] vssd vssd vccd vccd net1710 sky130_fd_sc_hd__buf_6
XFILLER_5_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1721 net1722 vssd vssd vccd vccd net1721 sky130_fd_sc_hd__buf_6
XFILLER_1_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1732 net1733 vssd vssd vccd vccd net1732 sky130_fd_sc_hd__buf_6
XFILLER_46_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1743 mprj_logic1\[454\] vssd vssd vccd vccd net1743 sky130_fd_sc_hd__buf_6
XFILLER_19_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1754 mprj_logic1\[449\] vssd vssd vccd vccd net1754 sky130_fd_sc_hd__buf_6
XTAP_3010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input411_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1765 net1766 vssd vssd vccd vccd net1765 sky130_fd_sc_hd__buf_6
XTAP_3021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1776 mprj_logic1\[438\] vssd vssd vccd vccd net1776 sky130_fd_sc_hd__buf_6
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1787 net1788 vssd vssd vccd vccd net1787 sky130_fd_sc_hd__buf_6
XFILLER_19_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1798 mprj_logic1\[425\] vssd vssd vccd vccd net1798 sky130_fd_sc_hd__buf_6
XTAP_3054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ net328 mprj_logic1\[120\] net72 vssd vssd vccd vccd net531 sky130_fd_sc_hd__and3b_4
XTAP_2397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_346_ mprj_logic1\[51\] net1344 vssd vssd vccd vccd net944 sky130_fd_sc_hd__and2_4
XFILLER_30_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_277_ net1763 net148 vssd vssd vccd vccd la_data_in_enable\[114\] sky130_fd_sc_hd__and2_4
XFILLER_31_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output463_A net1145 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1261_A net854 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1359_A net444 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1526_A net388 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1895_A net1896 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__034__A la_data_in_mprj_bar\[51\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1006 net795 vssd vssd vccd vccd net1006 sky130_fd_sc_hd__buf_6
Xwire1017 net783 vssd vssd vccd vccd net1017 sky130_fd_sc_hd__buf_6
Xwire1028 net763 vssd vssd vccd vccd net1028 sky130_fd_sc_hd__buf_6
XFILLER_38_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1039 net751 vssd vssd vccd vccd net1039 sky130_fd_sc_hd__buf_6
XFILLER_28_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1903 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__209__A mprj_logic1\[376\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_200_ mprj_logic1\[367\] net190 vssd vssd vccd vccd la_data_in_enable\[37\] sky130_fd_sc_hd__and2_4
XFILLER_51_2837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2007_A net2008 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_131_ mprj_dat_i_core_bar\[17\] vssd vssd vccd vccd net889 sky130_fd_sc_hd__clkinv_2
XFILLER_14_3393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input194_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_062_ net977 vssd vssd vccd vccd net695 sky130_fd_sc_hd__clkinv_2
XFILLER_7_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__386__A_N net296 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input361_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input459_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input55_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4010 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__598__B net1950 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1540 net362 vssd vssd vccd vccd net1540 sky130_fd_sc_hd__buf_8
XFILLER_24_1052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1551 net350 vssd vssd vccd vccd net1551 sky130_fd_sc_hd__buf_6
XFILLER_24_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1573 net31 vssd vssd vccd vccd net1573 sky130_fd_sc_hd__buf_6
XFILLER_19_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1584 net285 vssd vssd vccd vccd net1584 sky130_fd_sc_hd__buf_6
Xwire1595 net273 vssd vssd vccd vccd net1595 sky130_fd_sc_hd__buf_6
XFILLER_1_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__119__A mprj_dat_i_core_bar\[5\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output580_A net1076 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1107_A net521 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_329_ net1842 net1467 vssd vssd vccd vccd net864 sky130_fd_sc_hd__and2_4
XFILLER_31_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output845_A net845 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1476_A net402 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] net1322 vssd vssd vccd vccd la_data_in_mprj_bar\[92\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_45_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1643_A net1644 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__301__B net454 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1908_A net1909 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__211__B net202 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_810 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2124_A net2125 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input207_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_114_ mprj_dat_i_core_bar\[0\] vssd vssd vccd vccd net881 sky130_fd_sc_hd__clkinv_2
XFILLER_10_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_045_ la_data_in_mprj_bar\[62\] vssd vssd vccd vccd net677 sky130_fd_sc_hd__clkinv_2
XFILLER_10_2375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2060 net2061 vssd vssd vccd vccd net2060 sky130_fd_sc_hd__buf_6
Xwire2071 net2072 vssd vssd vccd vccd net2071 sky130_fd_sc_hd__buf_6
XFILLER_1_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2082 net2083 vssd vssd vccd vccd net2082 sky130_fd_sc_hd__buf_6
XFILLER_38_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2093 mprj_logic1\[193\] vssd vssd vccd vccd net2093 sky130_fd_sc_hd__buf_6
XANTENNA_wire1057_A net473 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__401__A_N net1570 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1370 net434 vssd vssd vccd vccd net1370 sky130_fd_sc_hd__buf_6
XFILLER_21_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1381 net1382 vssd vssd vccd vccd net1381 sky130_fd_sc_hd__buf_6
XFILLER_53_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1392 net1393 vssd vssd vccd vccd net1392 sky130_fd_sc_hd__buf_6
XFILLER_1_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1224_A net1225 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output795_A net1005 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[20\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_50_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1760_A mprj_logic1\[446\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1858_A mprj_logic1\[338\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__312__A mprj_logic1\[17\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__B net197 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3746 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2074_A net2075 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input157_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput301 la_oenb_mprj[21] vssd vssd vccd vccd net301 sky130_fd_sc_hd__clkbuf_4
XANTENNA__424__A_N net338 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput312 la_oenb_mprj[31] vssd vssd vccd vccd net312 sky130_fd_sc_hd__buf_6
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput323 la_oenb_mprj[41] vssd vssd vccd vccd net323 sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput334 la_oenb_mprj[51] vssd vssd vccd vccd net334 sky130_fd_sc_hd__buf_6
XFILLER_2_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput345 la_oenb_mprj[61] vssd vssd vccd vccd net345 sky130_fd_sc_hd__clkbuf_4
Xinput356 la_oenb_mprj[71] vssd vssd vccd vccd net356 sky130_fd_sc_hd__buf_6
Xinput367 la_oenb_mprj[81] vssd vssd vccd vccd net367 sky130_fd_sc_hd__buf_6
XANTENNA_input324_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput378 la_oenb_mprj[91] vssd vssd vccd vccd net378 sky130_fd_sc_hd__buf_6
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput389 mprj_adr_o_core[10] vssd vssd vccd vccd net389 sky130_fd_sc_hd__buf_6
XFILLER_53_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input18_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_594_ net384 net1963 vssd vssd vccd vccd net843 sky130_fd_sc_hd__and2_4
XFILLER_16_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1774 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_5 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput808 net808 vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__buf_8
Xoutput819 net819 vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__buf_8
X_028_ la_data_in_mprj_bar\[45\] vssd vssd vccd vccd net658 sky130_fd_sc_hd__inv_2
XFILLER_28_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output543_A net1084 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__132__A mprj_dat_i_core_bar\[18\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1174_A net1175 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output808_A net808 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1439_A net1440 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] la_data_in_enable\[55\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[55\] sky130_fd_sc_hd__nand2_2
XFILLER_48_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__307__A net2199 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1975_A mprj_logic1\[292\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__447__A_N net1539 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__217__A mprj_logic1\[384\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input274_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2191_A mprj_logic1\[143\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input441_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput120 la_data_out_mprj[8] vssd vssd vccd vccd net120 sky130_fd_sc_hd__clkbuf_4
Xinput131 la_data_out_mprj[9] vssd vssd vccd vccd net131 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput142 la_iena_mprj[109] vssd vssd vccd vccd net142 sky130_fd_sc_hd__clkbuf_4
Xinput153 la_iena_mprj[119] vssd vssd vccd vccd net153 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput164 la_iena_mprj[13] vssd vssd vccd vccd net164 sky130_fd_sc_hd__clkbuf_4
XTAP_4641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 la_iena_mprj[23] vssd vssd vccd vccd net175 sky130_fd_sc_hd__buf_6
XTAP_4652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 la_iena_mprj[33] vssd vssd vccd vccd net186 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput197 la_iena_mprj[43] vssd vssd vccd vccd net197 sky130_fd_sc_hd__buf_4
XTAP_4674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_577_ net1537 net1994 vssd vssd vccd vccd net825 sky130_fd_sc_hd__and2_4
XFILLER_32_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output493_A net493 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__127__A mprj_dat_i_core_bar\[13\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output660_A net660 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output758_A net1052 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1291_A net1292 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput605 net605 vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_8
XFILLER_9_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1389_A net1390 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput616 net616 vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_8
XFILLER_29_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput627 net627 vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_8
XFILLER_42_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput638 net638 vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_8
XFILLER_29_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output925_A net1190 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput649 net649 vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_8
XFILLER_42_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1723_A net1724 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__037__A la_data_in_mprj_bar\[54\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_B la_data_in_enable\[34\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_47_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1903 net1904 vssd vssd vccd vccd net1903 sky130_fd_sc_hd__buf_6
XANTENNA__500__A net321 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1914 mprj_logic1\[317\] vssd vssd vccd vccd net1914 sky130_fd_sc_hd__buf_6
XFILLER_8_1678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1925 net1926 vssd vssd vccd vccd net1925 sky130_fd_sc_hd__buf_6
XFILLER_41_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1936 mprj_logic1\[310\] vssd vssd vccd vccd net1936 sky130_fd_sc_hd__buf_6
XFILLER_6_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1947 mprj_logic1\[305\] vssd vssd vccd vccd net1947 sky130_fd_sc_hd__buf_6
XTAP_3203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1958 mprj_logic1\[300\] vssd vssd vccd vccd net1958 sky130_fd_sc_hd__buf_6
XTAP_3214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1969 net1970 vssd vssd vccd vccd net1969 sky130_fd_sc_hd__buf_6
XTAP_3225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_500_ net321 net2058 vssd vssd vccd vccd net780 sky130_fd_sc_hd__and2_4
XFILLER_19_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 net1865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 net2115 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_225 mprj_logic1\[365\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2037_A net2038 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 net1528 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_431_ net1555 mprj_logic1\[136\] net90 vssd vssd vccd vccd net549 sky130_fd_sc_hd__and3b_2
XTAP_2557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 net2016 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 net1575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ net1704 net1366 vssd vssd vccd vccd net930 sky130_fd_sc_hd__and2_2
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_293_ net1726 net462 vssd vssd vccd vccd user_irq_enable\[2\] sky130_fd_sc_hd__and2_1
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input391_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input85_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output506_A net1121 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1137_A net579 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1304_A net1305 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output875_A net875 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] la_data_in_enable\[18\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[18\] sky130_fd_sc_hd__nand2_2
XFILLER_31_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1673_A mprj_logic1\[81\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[16\]_B la_data_in_enable\[16\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_44_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[100\]_B la_data_in_enable\[100\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__304__B net457 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1840_A mprj_logic1\[351\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput468 net1062 vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__buf_8
XANTENNA_wire1938_A mprj_logic1\[309\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput479 net479 vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__buf_8
XFILLER_9_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__320__A mprj_logic1\[25\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__214__B net206 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__230__A net1815 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1700 net1701 vssd vssd vccd vccd net1700 sky130_fd_sc_hd__buf_6
Xwire1711 mprj_logic1\[62\] vssd vssd vccd vccd net1711 sky130_fd_sc_hd__buf_6
Xwire1722 mprj_logic1\[462\] vssd vssd vccd vccd net1722 sky130_fd_sc_hd__buf_6
XANTENNA_wire2154_A mprj_logic1\[160\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input237_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1733 net1734 vssd vssd vccd vccd net1733 sky130_fd_sc_hd__buf_6
Xwire1744 net1745 vssd vssd vccd vccd net1744 sky130_fd_sc_hd__buf_6
XFILLER_46_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1755 net1756 vssd vssd vccd vccd net1755 sky130_fd_sc_hd__buf_6
Xwire1766 mprj_logic1\[443\] vssd vssd vccd vccd net1766 sky130_fd_sc_hd__buf_6
XTAP_3011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1777 mprj_logic1\[437\] vssd vssd vccd vccd net1777 sky130_fd_sc_hd__buf_6
XTAP_3033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1788 mprj_logic1\[431\] vssd vssd vccd vccd net1788 sky130_fd_sc_hd__buf_6
XFILLER_41_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1799 mprj_logic1\[424\] vssd vssd vccd vccd net1799 sky130_fd_sc_hd__buf_6
XTAP_3055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input404_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ net327 mprj_logic1\[119\] net71 vssd vssd vccd vccd net530 sky130_fd_sc_hd__and3b_4
XFILLER_19_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ mprj_logic1\[50\] net1346 vssd vssd vccd vccd net943 sky130_fd_sc_hd__and2_2
XFILLER_50_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_276_ net1765 net147 vssd vssd vccd vccd la_data_in_enable\[113\] sky130_fd_sc_hd__and2_4
XFILLER_13_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1087_A net1088 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__140__A mprj_dat_i_core_bar\[26\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1254_A net1255 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2530 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1421_A net414 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1519_A net390 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1888_A mprj_logic1\[325\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__315__A mprj_logic1\[20\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1182 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__050__A la_data_in_mprj_bar\[67\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1007 net1008 vssd vssd vccd vccd net1007 sky130_fd_sc_hd__buf_6
XFILLER_5_1604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1018 net782 vssd vssd vccd vccd net1018 sky130_fd_sc_hd__buf_6
Xwire1029 net762 vssd vssd vccd vccd net1029 sky130_fd_sc_hd__buf_6
XFILLER_0_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1915 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__209__B net200 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_130_ mprj_dat_i_core_bar\[16\] vssd vssd vccd vccd net888 sky130_fd_sc_hd__clkinv_2
XFILLER_7_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__225__A mprj_logic1\[392\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_061_ net978 vssd vssd vccd vccd net694 sky130_fd_sc_hd__clkinv_2
XFILLER_27_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input187_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input354_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input48_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1530 net373 vssd vssd vccd vccd net1530 sky130_fd_sc_hd__buf_6
XFILLER_21_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1541 net361 vssd vssd vccd vccd net1541 sky130_fd_sc_hd__buf_8
XFILLER_47_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1552 net349 vssd vssd vccd vccd net1552 sky130_fd_sc_hd__buf_6
XFILLER_46_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1563 net328 vssd vssd vccd vccd net1563 sky130_fd_sc_hd__buf_6
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1574 net309 vssd vssd vccd vccd net1574 sky130_fd_sc_hd__buf_6
XFILLER_38_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1585 net284 vssd vssd vccd vccd net1585 sky130_fd_sc_hd__buf_6
XFILLER_47_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1596 net272 vssd vssd vccd vccd net1596 sky130_fd_sc_hd__buf_4
XFILLER_46_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1002_A net1003 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_328_ mprj_logic1\[33\] net1472 vssd vssd vccd vccd net863 sky130_fd_sc_hd__and2_4
XFILLER_15_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output573_A net573 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__135__A mprj_dat_i_core_bar\[21\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_259_ net1797 net255 vssd vssd vccd vccd la_data_in_enable\[96\] sky130_fd_sc_hd__and2_4
XFILLER_31_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output740_A net740 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output838_A net838 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1371_A net433 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1469_A net1470 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1014 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__480__A_N net1595 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] net1329 vssd vssd vccd vccd la_data_in_mprj_bar\[85\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__045__A la_data_in_mprj_bar\[62\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_822 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_538 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input102_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2117_A net2118 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_113_ user_irq_bar\[2\] vssd vssd vccd vccd net959 sky130_fd_sc_hd__inv_2
XFILLER_7_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_044_ la_data_in_mprj_bar\[61\] vssd vssd vccd vccd net676 sky130_fd_sc_hd__clkinv_2
XFILLER_10_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2050 mprj_logic1\[211\] vssd vssd vccd vccd net2050 sky130_fd_sc_hd__buf_6
XFILLER_43_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2061 mprj_logic1\[204\] vssd vssd vccd vccd net2061 sky130_fd_sc_hd__buf_6
Xwire2072 mprj_logic1\[200\] vssd vssd vccd vccd net2072 sky130_fd_sc_hd__buf_6
Xwire2083 net2084 vssd vssd vccd vccd net2083 sky130_fd_sc_hd__buf_6
Xwire2094 net2095 vssd vssd vccd vccd net2094 sky130_fd_sc_hd__buf_6
XFILLER_47_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1360 net1361 vssd vssd vccd vccd net1360 sky130_fd_sc_hd__buf_6
Xwire1371 net433 vssd vssd vccd vccd net1371 sky130_fd_sc_hd__buf_6
Xwire1382 net426 vssd vssd vccd vccd net1382 sky130_fd_sc_hd__buf_6
Xwire1393 net421 vssd vssd vccd vccd net1393 sky130_fd_sc_hd__buf_6
XFILLER_19_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1217_A net1218 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output690_A net690 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output788_A net788 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output955_A net1307 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[13\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_28_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1753_A net1754 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__312__B net1405 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[1\]_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1920_A net1921 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] la_data_in_enable\[111\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[111\] sky130_fd_sc_hd__nand2_2
XFILLER_6_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__376__A_N net365 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput302 la_oenb_mprj[22] vssd vssd vccd vccd net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput313 la_oenb_mprj[32] vssd vssd vccd vccd net313 sky130_fd_sc_hd__buf_6
XFILLER_2_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput324 la_oenb_mprj[42] vssd vssd vccd vccd net324 sky130_fd_sc_hd__buf_4
XFILLER_40_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput335 la_oenb_mprj[52] vssd vssd vccd vccd net335 sky130_fd_sc_hd__buf_4
XANTENNA_wire2067_A net2068 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput346 la_oenb_mprj[62] vssd vssd vccd vccd net346 sky130_fd_sc_hd__buf_6
Xinput357 la_oenb_mprj[72] vssd vssd vccd vccd net357 sky130_fd_sc_hd__buf_6
XFILLER_2_3565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput368 la_oenb_mprj[82] vssd vssd vccd vccd net368 sky130_fd_sc_hd__buf_6
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput379 la_oenb_mprj[92] vssd vssd vccd vccd net379 sky130_fd_sc_hd__buf_6
XFILLER_29_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input317_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_593_ net383 net1965 vssd vssd vccd vccd net842 sky130_fd_sc_hd__and2_4
XFILLER_35_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_6 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput809 net809 vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__buf_8
X_027_ la_data_in_mprj_bar\[44\] vssd vssd vccd vccd net657 sky130_fd_sc_hd__inv_2
XFILLER_29_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output536_A net1093 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1167_A net1168 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__399__A_N net1572 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1190 net1191 vssd vssd vccd vccd net1190 sky130_fd_sc_hd__buf_8
XFILLER_39_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] la_data_in_enable\[48\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[48\] sky130_fd_sc_hd__nand2_2
XFILLER_34_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1501_A net1502 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__307__B net1437 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1870_A mprj_logic1\[331\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1968_A mprj_logic1\[297\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__323__A mprj_logic1\[28\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__A net1810 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2184_A net2185 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input267_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input434_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput110 la_data_out_mprj[80] vssd vssd vccd vccd net110 sky130_fd_sc_hd__buf_6
Xinput121 la_data_out_mprj[90] vssd vssd vccd vccd net121 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input30_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput132 la_iena_mprj[0] vssd vssd vccd vccd net132 sky130_fd_sc_hd__clkbuf_4
Xinput143 la_iena_mprj[10] vssd vssd vccd vccd net143 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput154 la_iena_mprj[11] vssd vssd vccd vccd net154 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput165 la_iena_mprj[14] vssd vssd vccd vccd net165 sky130_fd_sc_hd__clkbuf_4
XTAP_4642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 la_iena_mprj[24] vssd vssd vccd vccd net176 sky130_fd_sc_hd__buf_6
XTAP_4653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput187 la_iena_mprj[34] vssd vssd vccd vccd net187 sky130_fd_sc_hd__clkbuf_4
XTAP_4664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput198 la_iena_mprj[44] vssd vssd vccd vccd net198 sky130_fd_sc_hd__buf_4
XFILLER_36_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_576_ net1538 net1996 vssd vssd vccd vccd net823 sky130_fd_sc_hd__and2_4
XFILLER_16_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output486_A net486 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output653_A net653 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput606 net606 vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_8
XANTENNA__143__A mprj_dat_i_core_bar\[29\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput617 net617 vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_8
XANTENNA_wire1284_A net1285 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput628 net628 vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_8
Xoutput639 net639 vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_8
XFILLER_25_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output820_A net820 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output918_A net1211 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1451_A net408 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1716_A mprj_logic1\[58\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__A_N net327 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__053__A la_data_in_mprj_bar\[70\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1904 mprj_logic1\[320\] vssd vssd vccd vccd net1904 sky130_fd_sc_hd__buf_6
XFILLER_8_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__500__B net2058 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1915 net1916 vssd vssd vccd vccd net1915 sky130_fd_sc_hd__buf_6
Xwire1926 net1927 vssd vssd vccd vccd net1926 sky130_fd_sc_hd__buf_6
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1937 net1938 vssd vssd vccd vccd net1937 sky130_fd_sc_hd__buf_6
Xwire1948 net1949 vssd vssd vccd vccd net1948 sky130_fd_sc_hd__buf_6
XTAP_3204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1959 net1960 vssd vssd vccd vccd net1959 sky130_fd_sc_hd__buf_6
XTAP_3215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 net1865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 net2115 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 mprj_logic1\[386\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 net1588 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ net345 mprj_logic1\[135\] net89 vssd vssd vccd vccd net548 sky130_fd_sc_hd__and3b_4
XANTENNA_248 net2136 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 mprj_logic1\[78\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__228__A mprj_logic1\[395\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_361_ net1706 net1367 vssd vssd vccd vccd net929 sky130_fd_sc_hd__and2_2
XFILLER_13_3212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_292_ net1729 net461 vssd vssd vccd vccd user_irq_enable\[1\] sky130_fd_sc_hd__and2_1
XFILLER_42_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input384_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input78_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__B mprj_logic1\[115\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1032_A net759 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__437__A_N net1549 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__138__A mprj_dat_i_core_bar\[24\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_559_ net1555 net2022 vssd vssd vccd vccd net805 sky130_fd_sc_hd__and2_4
XFILLER_14_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output868_A net868 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1499_A net1500 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1666_A net1667 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput469 net1061 vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__buf_8
XANTENNA__601__A net1603 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1833_A net1834 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__320__B net1505 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__048__A la_data_in_mprj_bar\[65\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__511__A net293 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__230__B net1610 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1701 mprj_logic1\[69\] vssd vssd vccd vccd net1701 sky130_fd_sc_hd__buf_6
XFILLER_43_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1712 mprj_logic1\[61\] vssd vssd vccd vccd net1712 sky130_fd_sc_hd__buf_6
Xwire1723 net1724 vssd vssd vccd vccd net1723 sky130_fd_sc_hd__buf_6
XFILLER_24_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1734 mprj_logic1\[458\] vssd vssd vccd vccd net1734 sky130_fd_sc_hd__buf_6
Xwire1745 mprj_logic1\[453\] vssd vssd vccd vccd net1745 sky130_fd_sc_hd__buf_6
XTAP_3001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input132_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1756 mprj_logic1\[448\] vssd vssd vccd vccd net1756 sky130_fd_sc_hd__buf_6
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1767 net1768 vssd vssd vccd vccd net1767 sky130_fd_sc_hd__buf_6
XANTENNA_wire2147_A net2148 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1778 net1779 vssd vssd vccd vccd net1778 sky130_fd_sc_hd__buf_6
XTAP_3034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1789 net1790 vssd vssd vccd vccd net1789 sky130_fd_sc_hd__buf_6
XFILLER_19_4144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_413_ net326 mprj_logic1\[118\] net70 vssd vssd vccd vccd net529 sky130_fd_sc_hd__and3b_4
XTAP_2377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ mprj_logic1\[49\] net1348 vssd vssd vccd vccd net942 sky130_fd_sc_hd__and2_2
XFILLER_53_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_3930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_275_ net1767 net146 vssd vssd vccd vccd la_data_in_enable\[112\] sky130_fd_sc_hd__and2_4
XFILLER_32_2964 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__405__B mprj_logic1\[110\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output616_A net616 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1247_A net1248 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1414_A net1415 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] la_data_in_enable\[30\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[30\] sky130_fd_sc_hd__nand2_4
XFILLER_33_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__315__B net1520 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1950_A net1951 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__331__A net1823 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1008 net794 vssd vssd vccd vccd net1008 sky130_fd_sc_hd__buf_6
Xwire1019 net779 vssd vssd vccd vccd net1019 sky130_fd_sc_hd__buf_6
XFILLER_5_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__A net387 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__225__B net218 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_060_ la_data_in_mprj_bar\[77\] vssd vssd vccd vccd net693 sky130_fd_sc_hd__clkinv_2
XFILLER_23_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2097_A net2098 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__241__A mprj_logic1\[408\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input347_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1520 net1521 vssd vssd vccd vccd net1520 sky130_fd_sc_hd__buf_6
XFILLER_21_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1531 net372 vssd vssd vccd vccd net1531 sky130_fd_sc_hd__buf_6
XFILLER_19_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1542 net360 vssd vssd vccd vccd net1542 sky130_fd_sc_hd__buf_8
XFILLER_21_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1553 net348 vssd vssd vccd vccd net1553 sky130_fd_sc_hd__buf_6
XFILLER_24_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1564 net325 vssd vssd vccd vccd net1564 sky130_fd_sc_hd__buf_4
XFILLER_24_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1575 net307 vssd vssd vccd vccd net1575 sky130_fd_sc_hd__buf_6
Xwire1586 net283 vssd vssd vccd vccd net1586 sky130_fd_sc_hd__buf_6
Xwire1597 net270 vssd vssd vccd vccd net1597 sky130_fd_sc_hd__buf_6
XFILLER_47_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_327_ mprj_logic1\[32\] net1475 vssd vssd vccd vccd net862 sky130_fd_sc_hd__and2_4
XFILLER_15_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_258_ net1798 net254 vssd vssd vccd vccd la_data_in_enable\[95\] sky130_fd_sc_hd__and2_4
XFILLER_10_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output566_A net566 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_189_ net1831 net1612 vssd vssd vccd vccd la_data_in_enable\[26\] sky130_fd_sc_hd__and2_2
XFILLER_45_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output733_A net733 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1364_A net440 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] la_data_in_enable\[78\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[78\] sky130_fd_sc_hd__nand2_2
XFILLER_6_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1531_A net372 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1629_A net104 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1998_A net1999 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__A mprj_logic1\[31\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__061__A net978 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2012_A net2013 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__236__A mprj_logic1\[403\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input297_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_112_ user_irq_bar\[1\] vssd vssd vccd vccd net958 sky130_fd_sc_hd__clkinv_2
XFILLER_51_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_043_ la_data_in_mprj_bar\[60\] vssd vssd vccd vccd net675 sky130_fd_sc_hd__inv_2
XFILLER_10_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input60_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__402__C net58 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2040 net2041 vssd vssd vccd vccd net2040 sky130_fd_sc_hd__buf_6
Xwire2051 mprj_logic1\[210\] vssd vssd vccd vccd net2051 sky130_fd_sc_hd__buf_6
XFILLER_21_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2062 net2063 vssd vssd vccd vccd net2062 sky130_fd_sc_hd__buf_6
Xwire2073 net2074 vssd vssd vccd vccd net2073 sky130_fd_sc_hd__buf_6
XFILLER_19_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2084 mprj_logic1\[196\] vssd vssd vccd vccd net2084 sky130_fd_sc_hd__buf_6
XFILLER_19_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1350 net1351 vssd vssd vccd vccd net1350 sky130_fd_sc_hd__buf_6
Xwire2095 net2096 vssd vssd vccd vccd net2095 sky130_fd_sc_hd__buf_6
Xwire1361 net443 vssd vssd vccd vccd net1361 sky130_fd_sc_hd__buf_6
XFILLER_47_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1372 net1373 vssd vssd vccd vccd net1372 sky130_fd_sc_hd__buf_6
XFILLER_1_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1383 net1384 vssd vssd vccd vccd net1383 sky130_fd_sc_hd__buf_6
XFILLER_46_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1394 net1395 vssd vssd vccd vccd net1394 sky130_fd_sc_hd__buf_6
XFILLER_19_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_870 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output683_A net683 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output850_A net1268 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output948_A net1280 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1746_A net1747 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1913_A net1914 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] la_data_in_enable\[104\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[104\] sky130_fd_sc_hd__nand2_8
XFILLER_17_3700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__056__A la_data_in_mprj_bar\[73\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__503__B net2053 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput303 la_oenb_mprj[23] vssd vssd vccd vccd net303 sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput314 la_oenb_mprj[33] vssd vssd vccd vccd net314 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput325 la_oenb_mprj[43] vssd vssd vccd vccd net325 sky130_fd_sc_hd__buf_6
Xinput336 la_oenb_mprj[53] vssd vssd vccd vccd net336 sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput347 la_oenb_mprj[63] vssd vssd vccd vccd net347 sky130_fd_sc_hd__buf_6
XFILLER_22_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput358 la_oenb_mprj[73] vssd vssd vccd vccd net358 sky130_fd_sc_hd__buf_6
Xinput369 la_oenb_mprj[83] vssd vssd vccd vccd net369 sky130_fd_sc_hd__buf_6
XFILLER_2_3588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input212_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_592_ net382 net1967 vssd vssd vccd vccd net841 sky130_fd_sc_hd__and2_4
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__A_N net1606 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_7 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_026_ la_data_in_mprj_bar\[43\] vssd vssd vccd vccd net656 sky130_fd_sc_hd__inv_2
XANTENNA__413__B mprj_logic1\[118\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output529_A net1100 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1062_A net468 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1180 net1181 vssd vssd vccd vccd net1180 sky130_fd_sc_hd__buf_6
Xwire1191 net1192 vssd vssd vccd vccd net1191 sky130_fd_sc_hd__buf_6
XFILLER_1_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1327_A la_data_in_enable\[87\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1696_A net1697 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__A net1600 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1863_A net1864 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__323__B net1494 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__493__A_N net1582 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__514__A net296 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__B net227 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input162_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2177_A net2178 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput100 la_data_out_mprj[71] vssd vssd vccd vccd net100 sky130_fd_sc_hd__buf_6
XFILLER_2_4042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput111 la_data_out_mprj[81] vssd vssd vccd vccd net111 sky130_fd_sc_hd__buf_6
XFILLER_44_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput122 la_data_out_mprj[91] vssd vssd vccd vccd net122 sky130_fd_sc_hd__clkbuf_4
XTAP_4610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 la_iena_mprj[100] vssd vssd vccd vccd net133 sky130_fd_sc_hd__buf_4
XFILLER_23_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput144 la_iena_mprj[110] vssd vssd vccd vccd net144 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input427_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 la_iena_mprj[120] vssd vssd vccd vccd net155 sky130_fd_sc_hd__clkbuf_4
XTAP_4632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 la_iena_mprj[15] vssd vssd vccd vccd net166 sky130_fd_sc_hd__clkbuf_4
XTAP_4643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input23_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput177 la_iena_mprj[25] vssd vssd vccd vccd net177 sky130_fd_sc_hd__buf_6
XTAP_4654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 la_iena_mprj[35] vssd vssd vccd vccd net188 sky130_fd_sc_hd__clkbuf_4
XTAP_4665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput199 la_iena_mprj[45] vssd vssd vccd vccd net199 sky130_fd_sc_hd__buf_4
XFILLER_29_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_575_ net1539 net1998 vssd vssd vccd vccd net822 sky130_fd_sc_hd__and2_4
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__408__B mprj_logic1\[113\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output479_A net479 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_29_4157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput607 net607 vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_8
XFILLER_9_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput618 net618 vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_8
Xoutput629 net629 vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_8
XFILLER_29_2733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output646_A net646 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_009_ la_data_in_mprj_bar\[26\] vssd vssd vccd vccd net637 sky130_fd_sc_hd__inv_4
XFILLER_46_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1277_A net877 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output813_A net1047 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1444_A net1445 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] la_data_in_enable\[60\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[60\] sky130_fd_sc_hd__nand2_2
XFILLER_23_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1709_A mprj_logic1\[64\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__318__B net1512 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1980_A mprj_logic1\[289\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__334__A net1812 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_max_length1311_A wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1905 net1906 vssd vssd vccd vccd net1905 sky130_fd_sc_hd__buf_6
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1916 net1917 vssd vssd vccd vccd net1916 sky130_fd_sc_hd__buf_6
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1927 mprj_logic1\[313\] vssd vssd vccd vccd net1927 sky130_fd_sc_hd__buf_6
XFILLER_41_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1938 mprj_logic1\[309\] vssd vssd vccd vccd net1938 sky130_fd_sc_hd__buf_6
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1949 mprj_logic1\[304\] vssd vssd vccd vccd net1949 sky130_fd_sc_hd__buf_6
XFILLER_19_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_205 net1865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_216 net2115 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__509__A net291 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_227 mprj_logic1\[386\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 net1589 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 net26 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__228__B net221 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ net1708 net1368 vssd vssd vccd vccd net928 sky130_fd_sc_hd__and2_2
XFILLER_17_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_291_ net1732 net460 vssd vssd vccd vccd user_irq_enable\[0\] sky130_fd_sc_hd__and2_1
XFILLER_52_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__A net1808 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__389__A_N net300 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input377_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__410__C net67 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_558_ net345 mprj_logic1\[263\] vssd vssd vccd vccd net804 sky130_fd_sc_hd__and2_2
XANTENNA_wire1025_A net767 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output596_A net596 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_489_ net1586 net2088 net1598 vssd vssd vccd vccd net486 sky130_fd_sc_hd__and3b_4
XFILLER_20_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output763_A net1028 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1394_A net1395 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output930_A net1170 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1561_A net1562 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1659_A net1660 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__601__B net1943 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1826_A mprj_logic1\[360\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__329__A net1842 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__064__A net975 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput960 net960 vssd vssd vccd vccd user_reset sky130_fd_sc_hd__buf_8
XFILLER_9_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__511__B net2040 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1702 net1703 vssd vssd vccd vccd net1702 sky130_fd_sc_hd__buf_6
XFILLER_5_3789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1713 mprj_logic1\[60\] vssd vssd vccd vccd net1713 sky130_fd_sc_hd__buf_6
XFILLER_8_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1724 net1725 vssd vssd vccd vccd net1724 sky130_fd_sc_hd__buf_6
XFILLER_1_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1735 net1736 vssd vssd vccd vccd net1735 sky130_fd_sc_hd__buf_6
XFILLER_24_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1746 net1747 vssd vssd vccd vccd net1746 sky130_fd_sc_hd__buf_6
XTAP_3002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1757 net1758 vssd vssd vccd vccd net1757 sky130_fd_sc_hd__buf_6
Xwire1768 mprj_logic1\[442\] vssd vssd vccd vccd net1768 sky130_fd_sc_hd__buf_6
XTAP_3013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1779 mprj_logic1\[436\] vssd vssd vccd vccd net1779 sky130_fd_sc_hd__buf_6
XTAP_3035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2042_A net2043 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__239__A mprj_logic1\[406\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ net325 mprj_logic1\[117\] net69 vssd vssd vccd vccd net528 sky130_fd_sc_hd__and3b_4
XTAP_2367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ mprj_logic1\[48\] net1350 vssd vssd vccd vccd net941 sky130_fd_sc_hd__and2_2
XFILLER_52_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input90_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_274_ net1769 net145 vssd vssd vccd vccd la_data_in_enable\[111\] sky130_fd_sc_hd__and2_4
XFILLER_52_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__405__C net61 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[6\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_10_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__421__B mprj_logic1\[126\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__404__A_N net1569 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output511_A net1116 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output609_A net609 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1142_A net524 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1407_A net1408 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output880_A net1306 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] la_data_in_enable\[23\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[23\] sky130_fd_sc_hd__nand2_4
XFILLER_18_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1776_A mprj_logic1\[438\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__612__A net1591 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1943_A net1944 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__331__B net1457 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1009 net1010 vssd vssd vccd vccd net1009 sky130_fd_sc_hd__buf_6
XFILLER_20_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__059__A la_data_in_mprj_bar\[76\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__B net2049 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__522__A net305 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__427__A_N net1556 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__241__B net235 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2200 mprj_logic1\[11\] vssd vssd vccd vccd net2200 sky130_fd_sc_hd__buf_6
Xoutput790 net1011 vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__buf_8
XFILLER_1_4118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input242_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1510 net1511 vssd vssd vccd vccd net1510 sky130_fd_sc_hd__buf_6
XFILLER_1_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1521 net389 vssd vssd vccd vccd net1521 sky130_fd_sc_hd__buf_6
Xwire1532 net371 vssd vssd vccd vccd net1532 sky130_fd_sc_hd__buf_6
XFILLER_4_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1543 net359 vssd vssd vccd vccd net1543 sky130_fd_sc_hd__buf_6
XFILLER_48_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1554 net347 vssd vssd vccd vccd net1554 sky130_fd_sc_hd__buf_6
Xwire1565 net322 vssd vssd vccd vccd net1565 sky130_fd_sc_hd__buf_6
XFILLER_4_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1576 net1577 vssd vssd vccd vccd net1576 sky130_fd_sc_hd__buf_6
XFILLER_38_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1587 net281 vssd vssd vccd vccd net1587 sky130_fd_sc_hd__buf_6
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1598 net27 vssd vssd vccd vccd net1598 sky130_fd_sc_hd__buf_4
XFILLER_21_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_326_ mprj_logic1\[31\] net1477 vssd vssd vccd vccd net861 sky130_fd_sc_hd__and2_4
XFILLER_9_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__416__B mprj_logic1\[121\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_257_ net1799 net253 vssd vssd vccd vccd la_data_in_enable\[94\] sky130_fd_sc_hd__and2_4
XFILLER_32_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_188_ net1833 net1613 vssd vssd vccd vccd la_data_in_enable\[25\] sky130_fd_sc_hd__and2_2
XANTENNA_output559_A net559 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1092_A net537 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output726_A net726 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1357_A net446 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1524_A net1525 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__A net1596 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1893_A net1894 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__B net1477 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire977_A la_data_in_mprj_bar\[79\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[91\]_B net1323 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__342__A mprj_logic1\[47\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__517__A net300 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__236__B net230 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2005_A net2006 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_111_ user_irq_bar\[0\] vssd vssd vccd vccd net957 sky130_fd_sc_hd__clkinv_2
XFILLER_14_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input192_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_042_ la_data_in_mprj_bar\[59\] vssd vssd vccd vccd net673 sky130_fd_sc_hd__inv_2
XFILLER_50_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__252__A mprj_logic1\[419\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input457_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input53_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2030 mprj_logic1\[225\] vssd vssd vccd vccd net2030 sky130_fd_sc_hd__buf_6
Xwire2041 mprj_logic1\[216\] vssd vssd vccd vccd net2041 sky130_fd_sc_hd__buf_6
Xwire2052 mprj_logic1\[209\] vssd vssd vccd vccd net2052 sky130_fd_sc_hd__buf_6
XFILLER_38_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2063 mprj_logic1\[203\] vssd vssd vccd vccd net2063 sky130_fd_sc_hd__buf_6
Xwire2074 net2075 vssd vssd vccd vccd net2074 sky130_fd_sc_hd__buf_6
XFILLER_21_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1340 net85 vssd vssd vccd vccd net1340 sky130_fd_sc_hd__buf_6
Xwire2085 net2086 vssd vssd vccd vccd net2085 sky130_fd_sc_hd__buf_6
Xwire1351 net449 vssd vssd vccd vccd net1351 sky130_fd_sc_hd__buf_6
Xwire2096 mprj_logic1\[192\] vssd vssd vccd vccd net2096 sky130_fd_sc_hd__buf_6
Xwire1362 net442 vssd vssd vccd vccd net1362 sky130_fd_sc_hd__buf_6
XFILLER_43_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1373 net1374 vssd vssd vccd vccd net1373 sky130_fd_sc_hd__buf_6
XFILLER_47_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1384 net425 vssd vssd vccd vccd net1384 sky130_fd_sc_hd__buf_6
XFILLER_46_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1395 net1396 vssd vssd vccd vccd net1395 sky130_fd_sc_hd__buf_6
XFILLER_38_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_882 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1105_A net523 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_309_ net2179 net1417 vssd vssd vccd vccd net874 sky130_fd_sc_hd__and2_2
XFILLER_30_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[73\]_B la_data_in_enable\[73\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_47_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output843_A net843 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__162__A la_data_in_mprj_bar\[15\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1474_A net403 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] net1324 vssd vssd vccd vccd la_data_in_mprj_bar\[90\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1641_A net1642 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1739_A mprj_logic1\[456\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1906_A net1907 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__337__A mprj_logic1\[42\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__072__A net968 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput304 la_oenb_mprj[24] vssd vssd vccd vccd net304 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput315 la_oenb_mprj[34] vssd vssd vccd vccd net315 sky130_fd_sc_hd__buf_4
XFILLER_44_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput326 la_oenb_mprj[44] vssd vssd vccd vccd net326 sky130_fd_sc_hd__buf_6
Xinput337 la_oenb_mprj[54] vssd vssd vccd vccd net337 sky130_fd_sc_hd__buf_8
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput348 la_oenb_mprj[64] vssd vssd vccd vccd net348 sky130_fd_sc_hd__buf_6
XFILLER_40_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput359 la_oenb_mprj[74] vssd vssd vccd vccd net359 sky130_fd_sc_hd__buf_6
XFILLER_5_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_591_ net381 net1969 vssd vssd vccd vccd net840 sky130_fd_sc_hd__and2_4
XFILLER_35_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2122_A mprj_logic1\[181\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input205_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__247__A mprj_logic1\[414\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_025_ la_data_in_mprj_bar\[42\] vssd vssd vccd vccd net655 sky130_fd_sc_hd__inv_2
XANTENNA_8 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__413__C net70 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2766 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1170 net1171 vssd vssd vccd vccd net1170 sky130_fd_sc_hd__buf_8
XFILLER_19_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1181 net928 vssd vssd vccd vccd net1181 sky130_fd_sc_hd__buf_6
XFILLER_47_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1192 net1193 vssd vssd vccd vccd net1192 sky130_fd_sc_hd__buf_6
XFILLER_1_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__295__A_N net1576 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1222_A net915 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output793_A net793 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1689_A mprj_logic1\[74\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__B net1937 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1856_A mprj_logic1\[340\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__A net1583 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__067__A net973 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[37\]_B la_data_in_enable\[37\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_3174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[121\]_B la_data_in_enable\[121\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__514__B net2036 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A net314 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input155_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vssd vccd vccd net101 sky130_fd_sc_hd__buf_6
XFILLER_7_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput112 la_data_out_mprj[82] vssd vssd vccd vccd net112 sky130_fd_sc_hd__buf_6
Xinput123 la_data_out_mprj[92] vssd vssd vccd vccd net123 sky130_fd_sc_hd__clkbuf_4
XTAP_4600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput134 la_iena_mprj[101] vssd vssd vccd vccd net134 sky130_fd_sc_hd__clkbuf_4
XTAP_4611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 la_iena_mprj[111] vssd vssd vccd vccd net145 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput156 la_iena_mprj[121] vssd vssd vccd vccd net156 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input322_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput167 la_iena_mprj[16] vssd vssd vccd vccd net167 sky130_fd_sc_hd__clkbuf_4
XTAP_4644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 la_iena_mprj[26] vssd vssd vccd vccd net178 sky130_fd_sc_hd__buf_6
XTAP_4655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 la_iena_mprj[36] vssd vssd vccd vccd net189 sky130_fd_sc_hd__clkbuf_4
XTAP_4666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_574_ net1540 net2001 vssd vssd vccd vccd net821 sky130_fd_sc_hd__and2_4
XANTENNA_user_wb_dat_gates\[30\]_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__424__B mprj_logic1\[129\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B la_data_in_enable\[112\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_8_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput608 net608 vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_8
Xoutput619 net619 vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_8
X_008_ la_data_in_mprj_bar\[25\] vssd vssd vccd vccd net636 sky130_fd_sc_hd__inv_4
XFILLER_29_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output541_A net1087 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output639_A net639 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1172_A net1173 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output806_A net806 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1437_A net1438 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] la_data_in_enable\[53\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[53\] sky130_fd_sc_hd__nand2_4
XFILLER_48_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1604_A net264 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[21\]_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__615__A net1588 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1973_A net1974 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[19\]_B la_data_in_enable\[19\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_30_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__334__B net1442 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B net1316 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__350__A net1719 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__460__A_N net378 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input8_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1906 net1907 vssd vssd vccd vccd net1906 sky130_fd_sc_hd__buf_6
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1917 net1918 vssd vssd vccd vccd net1917 sky130_fd_sc_hd__buf_6
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1928 net1929 vssd vssd vccd vccd net1928 sky130_fd_sc_hd__buf_6
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1939 net1940 vssd vssd vccd vccd net1939 sky130_fd_sc_hd__buf_6
XFILLER_41_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 net1865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 net2116 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 mprj_logic1\[47\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__509__B net2044 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_239 net1592 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_290_ net1735 net162 vssd vssd vccd vccd la_data_in_enable\[127\] sky130_fd_sc_hd__and2_4
XFILLER_17_2682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__525__A net308 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__B net239 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input272_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__260__A net1795 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__419__B mprj_logic1\[124\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_557_ net344 mprj_logic1\[262\] vssd vssd vccd vccd net803 sky130_fd_sc_hd__and2_2
XFILLER_31_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1018_A net782 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_488_ net1587 net2091 net1608 vssd vssd vccd vccd net484 sky130_fd_sc_hd__and3b_4
XANTENNA_output491_A net491 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output589_A net1067 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output756_A net1034 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1387_A net1388 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__483__A_N net1592 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output923_A net1194 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__170__A net1859 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1721_A net1722 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__329__B net1467 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__345__A mprj_logic1\[50\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__080__A la_data_in_mprj_bar\[97\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput950 net1299 vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__buf_8
XFILLER_25_4375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1703 mprj_logic1\[68\] vssd vssd vccd vccd net1703 sky130_fd_sc_hd__buf_6
XFILLER_43_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1714 mprj_logic1\[5\] vssd vssd vccd vccd net1714 sky130_fd_sc_hd__buf_6
Xwire1725 net951 vssd vssd vccd vccd net1725 sky130_fd_sc_hd__buf_6
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1736 net1737 vssd vssd vccd vccd net1736 sky130_fd_sc_hd__buf_6
XFILLER_41_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1747 net1748 vssd vssd vccd vccd net1747 sky130_fd_sc_hd__buf_6
XTAP_3003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1758 mprj_logic1\[447\] vssd vssd vccd vccd net1758 sky130_fd_sc_hd__buf_6
XFILLER_2_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1769 net1770 vssd vssd vccd vccd net1769 sky130_fd_sc_hd__buf_6
XTAP_3014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__239__B net233 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2035_A mprj_logic1\[220\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ net324 mprj_logic1\[116\] net68 vssd vssd vccd vccd net527 sky130_fd_sc_hd__and3b_4
XFILLER_27_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_342_ mprj_logic1\[47\] net1352 vssd vssd vccd vccd net940 sky130_fd_sc_hd__and2_2
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__255__A net1801 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_273_ net1771 net144 vssd vssd vccd vccd la_data_in_enable\[110\] sky130_fd_sc_hd__and2_4
XFILLER_32_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input83_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__421__C net79 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output504_A net1123 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1135_A net474 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_609_ net1594 net1922 vssd vssd vccd vccd net733 sky130_fd_sc_hd__and2_4
XFILLER_53_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1302_A net950 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output873_A net873 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__165__A net1867 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] la_data_in_enable\[16\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[16\] sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[29\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_31_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1671_A mprj_logic1\[82\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1769_A net1770 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__612__B net1911 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1936_A mprj_logic1\[310\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] la_data_in_enable\[127\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[127\] sky130_fd_sc_hd__nand2_1
XFILLER_0_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__379__A_N net271 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__075__A net965 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_950 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__522__B mprj_logic1\[227\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput780 net1050 vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__buf_8
Xwire2201 net2202 vssd vssd vccd vccd net2201 sky130_fd_sc_hd__buf_6
Xoutput791 net1049 vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__buf_8
XFILLER_40_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1500 net396 vssd vssd vccd vccd net1500 sky130_fd_sc_hd__buf_6
XFILLER_8_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1511 net393 vssd vssd vccd vccd net1511 sky130_fd_sc_hd__buf_6
XFILLER_48_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input235_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1522 net1523 vssd vssd vccd vccd net1522 sky130_fd_sc_hd__buf_8
XFILLER_24_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2152_A net2153 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1533 net370 vssd vssd vccd vccd net1533 sky130_fd_sc_hd__buf_6
XFILLER_4_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1544 net358 vssd vssd vccd vccd net1544 sky130_fd_sc_hd__buf_6
XFILLER_38_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1555 net346 vssd vssd vccd vccd net1555 sky130_fd_sc_hd__buf_6
Xwire1566 net32 vssd vssd vccd vccd net1566 sky130_fd_sc_hd__buf_6
Xwire1577 net1578 vssd vssd vccd vccd net1577 sky130_fd_sc_hd__buf_6
XFILLER_24_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1588 net280 vssd vssd vccd vccd net1588 sky130_fd_sc_hd__buf_6
XFILLER_41_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1599 net269 vssd vssd vccd vccd net1599 sky130_fd_sc_hd__buf_4
XFILLER_41_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input402_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ mprj_logic1\[30\] net1482 vssd vssd vccd vccd net860 sky130_fd_sc_hd__and2_4
XFILLER_30_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__416__C net73 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_256_ net1800 net252 vssd vssd vccd vccd la_data_in_enable\[93\] sky130_fd_sc_hd__and2_4
XFILLER_7_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_187_ net1835 net1614 vssd vssd vccd vccd la_data_in_enable\[24\] sky130_fd_sc_hd__and2_2
XFILLER_48_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__432__B net2198 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1085_A net1086 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output719_A net1053 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1252_A net913 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1517_A net391 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__B net1928 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1886_A net1887 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__A net1580 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__342__B net1352 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[4\]_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__517__B net2033 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_110_ net979 vssd vssd vccd vccd net621 sky130_fd_sc_hd__clkinv_2
XFILLER_36_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__533__A net1568 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_041_ la_data_in_mprj_bar\[58\] vssd vssd vccd vccd net672 sky130_fd_sc_hd__inv_2
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__252__B net247 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input352_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input46_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2020 mprj_logic1\[266\] vssd vssd vccd vccd net2020 sky130_fd_sc_hd__buf_6
XFILLER_1_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2031 mprj_logic1\[224\] vssd vssd vccd vccd net2031 sky130_fd_sc_hd__buf_6
XFILLER_43_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2042 net2043 vssd vssd vccd vccd net2042 sky130_fd_sc_hd__buf_6
Xwire2053 net2054 vssd vssd vccd vccd net2053 sky130_fd_sc_hd__buf_6
XFILLER_1_3226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2064 net2065 vssd vssd vccd vccd net2064 sky130_fd_sc_hd__buf_6
Xwire1330 la_data_in_enable\[84\] vssd vssd vccd vccd net1330 sky130_fd_sc_hd__buf_8
Xwire2075 mprj_logic1\[199\] vssd vssd vccd vccd net2075 sky130_fd_sc_hd__buf_6
Xwire1341 net459 vssd vssd vccd vccd net1341 sky130_fd_sc_hd__buf_6
Xwire2086 net2087 vssd vssd vccd vccd net2086 sky130_fd_sc_hd__buf_6
XFILLER_21_3187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1352 net1353 vssd vssd vccd vccd net1352 sky130_fd_sc_hd__buf_6
XFILLER_5_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2097 net2098 vssd vssd vccd vccd net2097 sky130_fd_sc_hd__buf_6
XFILLER_21_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1363 net441 vssd vssd vccd vccd net1363 sky130_fd_sc_hd__buf_6
Xwire1374 net432 vssd vssd vccd vccd net1374 sky130_fd_sc_hd__buf_6
XFILLER_21_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1385 net1386 vssd vssd vccd vccd net1385 sky130_fd_sc_hd__buf_6
Xwire1396 net1397 vssd vssd vccd vccd net1396 sky130_fd_sc_hd__buf_6
XFILLER_46_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__427__B mprj_logic1\[132\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2814 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_308_ net2195 net1422 vssd vssd vccd vccd net873 sky130_fd_sc_hd__and2_4
XANTENNA_wire1000_A net1001 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output571_A net571 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_239_ mprj_logic1\[406\] net233 vssd vssd vccd vccd la_data_in_enable\[76\] sky130_fd_sc_hd__and2_4
XFILLER_10_3592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output836_A net994 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1467_A net1468 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] net1331 vssd vssd vccd vccd la_data_in_mprj_bar\[83\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_3098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1634_A mprj_logic1\[9\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__618__A net1585 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__337__B net1391 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__417__A_N net330 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__353__A net1716 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput305 la_oenb_mprj[25] vssd vssd vccd vccd net305 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput316 la_oenb_mprj[35] vssd vssd vccd vccd net316 sky130_fd_sc_hd__buf_6
XFILLER_2_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput327 la_oenb_mprj[45] vssd vssd vccd vccd net327 sky130_fd_sc_hd__buf_4
XFILLER_22_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput338 la_oenb_mprj[55] vssd vssd vccd vccd net338 sky130_fd_sc_hd__buf_4
XFILLER_5_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput349 la_oenb_mprj[65] vssd vssd vccd vccd net349 sky130_fd_sc_hd__buf_6
XFILLER_2_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_590_ net380 net1971 vssd vssd vccd vccd net839 sky130_fd_sc_hd__and2_4
XFILLER_2_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__A net1571 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input100_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2115_A net2116 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__263__A net1789 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_024_ la_data_in_mprj_bar\[41\] vssd vssd vccd vccd net654 sky130_fd_sc_hd__inv_2
XANTENNA_9 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1160 net1161 vssd vssd vccd vccd net1160 sky130_fd_sc_hd__buf_6
Xwire1171 net1172 vssd vssd vccd vccd net1171 sky130_fd_sc_hd__buf_6
Xwire1182 net1183 vssd vssd vccd vccd net1182 sky130_fd_sc_hd__buf_8
XFILLER_1_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1193 net925 vssd vssd vccd vccd net1193 sky130_fd_sc_hd__buf_6
XFILLER_47_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1048_A net802 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1215_A net1216 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output786_A net1013 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output953_A net2205 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__173__A net1856 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[11\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_51_2991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1751_A net1752 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1849_A mprj_logic1\[344\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__B net1886 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__348__A mprj_logic1\[53\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__083__A net993 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__530__B mprj_logic1\[235\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput102 la_data_out_mprj[73] vssd vssd vccd vccd net102 sky130_fd_sc_hd__buf_6
XFILLER_24_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput113 la_data_out_mprj[83] vssd vssd vccd vccd net113 sky130_fd_sc_hd__buf_6
XFILLER_7_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput124 la_data_out_mprj[93] vssd vssd vccd vccd net124 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2065_A mprj_logic1\[202\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input148_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput135 la_iena_mprj[102] vssd vssd vccd vccd net135 sky130_fd_sc_hd__clkbuf_4
XTAP_4612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput146 la_iena_mprj[112] vssd vssd vccd vccd net146 sky130_fd_sc_hd__buf_4
XFILLER_22_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 la_iena_mprj[122] vssd vssd vccd vccd net157 sky130_fd_sc_hd__buf_4
XTAP_4634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 la_iena_mprj[17] vssd vssd vccd vccd net168 sky130_fd_sc_hd__clkbuf_4
XTAP_4645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 la_iena_mprj[27] vssd vssd vccd vccd net179 sky130_fd_sc_hd__buf_4
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input315_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__258__A net1798 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_573_ net1541 net2003 vssd vssd vccd vccd net820 sky130_fd_sc_hd__and2_4
XTAP_3988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__424__C net82 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput609 net609 vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_8
XFILLER_29_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_007_ la_data_in_mprj_bar\[24\] vssd vssd vccd vccd net635 sky130_fd_sc_hd__clkinv_4
XFILLER_46_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__B net2188 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output534_A net1095 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1165_A net932 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1332_A la_data_in_enable\[80\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__168__A net1862 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] la_data_in_enable\[46\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[46\] sky130_fd_sc_hd__nand2_2
XFILLER_1_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__615__B net1902 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] la_data_in_enable\[8\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[8\] sky130_fd_sc_hd__nand2_2
XANTENNA__350__B net1383 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1907 mprj_logic1\[319\] vssd vssd vccd vccd net1907 sky130_fd_sc_hd__buf_6
XFILLER_41_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1918 mprj_logic1\[316\] vssd vssd vccd vccd net1918 sky130_fd_sc_hd__buf_6
Xwire1929 net1930 vssd vssd vccd vccd net1929 sky130_fd_sc_hd__buf_6
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__078__A net962 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_207 net1951 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 net2125 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_978 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_229 mprj_logic1\[78\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__525__B net2027 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__541__A net326 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2182_A net2183 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__260__B net256 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input432_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_625_ net1871 net132 vssd vssd vccd vccd la_data_in_enable\[0\] sky130_fd_sc_hd__and2_1
XTAP_3763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__419__C net77 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_556_ net342 mprj_logic1\[261\] vssd vssd vccd vccd net801 sky130_fd_sc_hd__and2_2
XFILLER_50_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_487_ net1588 net2094 net24 vssd vssd vccd vccd net483 sky130_fd_sc_hd__and3b_4
XFILLER_32_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__435__B net2194 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output484_A net484 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output651_A net651 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output749_A net749 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1282_A net1283 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output916_A net1217 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1714_A mprj_logic1\[5\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4258 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__345__B net1346 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__361__A net1706 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput940 net1238 vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__buf_8
XFILLER_5_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput951 net1723 vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_47_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1704 net1705 vssd vssd vccd vccd net1704 sky130_fd_sc_hd__buf_6
XFILLER_28_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1715 mprj_logic1\[59\] vssd vssd vccd vccd net1715 sky130_fd_sc_hd__buf_6
XFILLER_25_2985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1726 net1727 vssd vssd vccd vccd net1726 sky130_fd_sc_hd__buf_6
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1737 mprj_logic1\[457\] vssd vssd vccd vccd net1737 sky130_fd_sc_hd__buf_6
Xwire1748 mprj_logic1\[452\] vssd vssd vccd vccd net1748 sky130_fd_sc_hd__buf_6
XTAP_3004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1759 net1760 vssd vssd vccd vccd net1759 sky130_fd_sc_hd__buf_6
XFILLER_19_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ net323 mprj_logic1\[115\] net67 vssd vssd vccd vccd net526 sky130_fd_sc_hd__and3b_4
XTAP_2347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ mprj_logic1\[46\] net1354 vssd vssd vccd vccd net939 sky130_fd_sc_hd__and2_2
XFILLER_36_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__255__B net251 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_272_ net1773 net142 vssd vssd vccd vccd la_data_in_enable\[109\] sky130_fd_sc_hd__and2_4
XFILLER_10_3922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input382_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input76_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__271__A net1775 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_608_ net1595 net1925 vssd vssd vccd vccd net732 sky130_fd_sc_hd__and2_4
XTAP_3593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1030_A net761 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1128_A net498 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_539_ net324 net2024 vssd vssd vccd vccd net783 sky130_fd_sc_hd__and2_2
XFILLER_32_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__450__A_N net1536 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output866_A net866 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1497_A net397 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__181__A net1844 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1664_A net1665 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1831_A net1832 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1929_A net1930 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__356__A net1712 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__091__A net990 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput770 net770 vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__buf_8
Xoutput781 net781 vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__buf_8
XFILLER_47_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2202 mprj_logic1\[10\] vssd vssd vccd vccd net2202 sky130_fd_sc_hd__buf_6
Xoutput792 net1009 vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__buf_8
XFILLER_43_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1501 net1502 vssd vssd vccd vccd net1501 sky130_fd_sc_hd__buf_6
Xwire1512 net1513 vssd vssd vccd vccd net1512 sky130_fd_sc_hd__buf_6
XFILLER_38_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1523 net1524 vssd vssd vccd vccd net1523 sky130_fd_sc_hd__buf_6
XFILLER_21_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1534 net369 vssd vssd vccd vccd net1534 sky130_fd_sc_hd__buf_6
Xwire1545 net357 vssd vssd vccd vccd net1545 sky130_fd_sc_hd__buf_6
XFILLER_4_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input130_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1556 net341 vssd vssd vccd vccd net1556 sky130_fd_sc_hd__buf_6
XFILLER_38_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2145_A mprj_logic1\[163\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1567 net318 vssd vssd vccd vccd net1567 sky130_fd_sc_hd__buf_6
XFILLER_21_2668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1578 net3 vssd vssd vccd vccd net1578 sky130_fd_sc_hd__buf_6
XANTENNA_input228_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1589 net279 vssd vssd vccd vccd net1589 sky130_fd_sc_hd__buf_6
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__473__A_N net1603 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__266__A net1784 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ mprj_logic1\[29\] net1490 vssd vssd vccd vccd net858 sky130_fd_sc_hd__and2_4
XFILLER_32_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_255_ net1801 net251 vssd vssd vccd vccd la_data_in_enable\[92\] sky130_fd_sc_hd__and2_4
XFILLER_10_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_186_ net1837 net1615 vssd vssd vccd vccd la_data_in_enable\[23\] sky130_fd_sc_hd__and2_2
XFILLER_7_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__432__C net91 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1245_A net938 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1412_A net1413 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__176__A net1850 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1781_A mprj_logic1\[435\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1879_A net1880 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__B net1876 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[4\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__496__A_N net1579 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__086__A net992 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_040_ la_data_in_mprj_bar\[57\] vssd vssd vccd vccd net671 sky130_fd_sc_hd__inv_2
XFILLER_49_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2095_A net2096 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input178_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input345_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2010 net2011 vssd vssd vccd vccd net2010 sky130_fd_sc_hd__buf_6
Xwire2021 mprj_logic1\[265\] vssd vssd vccd vccd net2021 sky130_fd_sc_hd__buf_6
Xwire2032 mprj_logic1\[223\] vssd vssd vccd vccd net2032 sky130_fd_sc_hd__buf_6
XFILLER_21_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input39_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2043 mprj_logic1\[215\] vssd vssd vccd vccd net2043 sky130_fd_sc_hd__buf_6
Xwire2054 mprj_logic1\[208\] vssd vssd vccd vccd net2054 sky130_fd_sc_hd__buf_6
XFILLER_43_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1320 la_data_in_enable\[94\] vssd vssd vccd vccd net1320 sky130_fd_sc_hd__buf_6
Xwire2065 mprj_logic1\[202\] vssd vssd vccd vccd net2065 sky130_fd_sc_hd__buf_6
Xwire2076 net2077 vssd vssd vccd vccd net2076 sky130_fd_sc_hd__buf_6
Xwire1331 la_data_in_enable\[83\] vssd vssd vccd vccd net1331 sky130_fd_sc_hd__buf_6
XFILLER_1_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1342 net1343 vssd vssd vccd vccd net1342 sky130_fd_sc_hd__buf_6
Xwire2087 mprj_logic1\[195\] vssd vssd vccd vccd net2087 sky130_fd_sc_hd__buf_6
XFILLER_1_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1353 net448 vssd vssd vccd vccd net1353 sky130_fd_sc_hd__buf_6
Xwire2098 mprj_logic1\[191\] vssd vssd vccd vccd net2098 sky130_fd_sc_hd__buf_6
XFILLER_5_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1364 net440 vssd vssd vccd vccd net1364 sky130_fd_sc_hd__buf_6
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1375 net431 vssd vssd vccd vccd net1375 sky130_fd_sc_hd__buf_6
Xwire1386 net424 vssd vssd vccd vccd net1386 sky130_fd_sc_hd__buf_6
Xwire1397 net420 vssd vssd vccd vccd net1397 sky130_fd_sc_hd__buf_6
XFILLER_1_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__427__C net1340 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_307_ net2199 net1437 vssd vssd vccd vccd net870 sky130_fd_sc_hd__and2_2
XFILLER_50_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_238_ mprj_logic1\[405\] net232 vssd vssd vccd vccd la_data_in_enable\[75\] sky130_fd_sc_hd__and2_4
XANTENNA__443__B net2182 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output564_A net564 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__369__A_N net260 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_169_ net1861 net226 vssd vssd vccd vccd la_data_in_enable\[6\] sky130_fd_sc_hd__and2_2
XFILLER_7_796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1195_A net1196 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output731_A net731 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output829_A net829 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] la_data_in_enable\[76\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[76\] sky130_fd_sc_hd__nand2_8
XFILLER_23_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1627_A net106 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__618__B net1892 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1996_A net1997 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__353__B net1378 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput306 la_oenb_mprj[26] vssd vssd vccd vccd net306 sky130_fd_sc_hd__buf_4
Xinput317 la_oenb_mprj[36] vssd vssd vccd vccd net317 sky130_fd_sc_hd__buf_6
Xinput328 la_oenb_mprj[46] vssd vssd vccd vccd net328 sky130_fd_sc_hd__buf_6
Xinput339 la_oenb_mprj[56] vssd vssd vccd vccd net339 sky130_fd_sc_hd__buf_4
XFILLER_22_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__B mprj_logic1\[233\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2010_A net2011 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2108_A net2109 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__544__A net1561 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input295_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__263__B net133 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_023_ la_data_in_mprj_bar\[40\] vssd vssd vccd vccd net653 sky130_fd_sc_hd__inv_2
XANTENNA_input462_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1150 net1151 vssd vssd vccd vccd net1150 sky130_fd_sc_hd__buf_8
XFILLER_48_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1161 net933 vssd vssd vccd vccd net1161 sky130_fd_sc_hd__buf_6
XFILLER_40_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1172 net1173 vssd vssd vccd vccd net1172 sky130_fd_sc_hd__buf_6
XFILLER_1_2334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1183 net1184 vssd vssd vccd vccd net1183 sky130_fd_sc_hd__buf_6
Xwire1194 net1195 vssd vssd vccd vccd net1194 sky130_fd_sc_hd__buf_8
XFILLER_34_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__438__B net2191 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1110_A net518 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1208_A net1209 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output779_A net1019 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output946_A net1289 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1577_A net1578 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1744_A net1745 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1911_A net1912 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] la_data_in_enable\[102\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[102\] sky130_fd_sc_hd__nand2_4
XANTENNA__348__B net1387 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__364__A net1700 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput103 la_data_out_mprj[74] vssd vssd vccd vccd net103 sky130_fd_sc_hd__buf_6
Xinput114 la_data_out_mprj[84] vssd vssd vccd vccd net114 sky130_fd_sc_hd__buf_6
XFILLER_24_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput125 la_data_out_mprj[94] vssd vssd vccd vccd net125 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 la_iena_mprj[103] vssd vssd vccd vccd net136 sky130_fd_sc_hd__clkbuf_4
XTAP_4613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput147 la_iena_mprj[113] vssd vssd vccd vccd net147 sky130_fd_sc_hd__buf_4
XTAP_4624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 la_iena_mprj[123] vssd vssd vccd vccd net158 sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput169 la_iena_mprj[18] vssd vssd vccd vccd net169 sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire2058_A net2059 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__539__A net324 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input210_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_572_ net1542 net2005 vssd vssd vccd vccd net819 sky130_fd_sc_hd__and2_4
XFILLER_29_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input308_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__274__A net1769 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_006_ la_data_in_mprj_bar\[23\] vssd vssd vccd vccd net634 sky130_fd_sc_hd__clkinv_4
XFILLER_29_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__C net1633 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__407__A_N net319 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output527_A net1102 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1060_A net470 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1158_A net1159 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1325_A la_data_in_enable\[89\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output896_A net896 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] la_data_in_enable\[39\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[39\] sky130_fd_sc_hd__nand2_2
XFILLER_23_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__184__A net1840 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1694_A net1695 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1861_A mprj_logic1\[336\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1959_A net1960 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1908 net1909 vssd vssd vccd vccd net1908 sky130_fd_sc_hd__buf_6
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1919 net1920 vssd vssd vccd vccd net1919 sky130_fd_sc_hd__buf_6
XFILLER_41_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__359__A net1709 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 net1954 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 net2132 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__094__A net988 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input160_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input258_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2175_A net2176 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input425_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__269__A net1778 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_624_ net1579 net1872 vssd vssd vccd vccd net749 sky130_fd_sc_hd__and2_4
XTAP_4498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_555_ net1556 mprj_logic1\[260\] vssd vssd vccd vccd net800 sky130_fd_sc_hd__and2_4
XFILLER_35_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_486_ net1589 net2097 net23 vssd vssd vccd vccd net482 sky130_fd_sc_hd__and3b_4
XFILLER_18_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__435__C net1338 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output477_A net1054 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__451__B net2165 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output644_A net644 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1275_A net879 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output811_A net811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1442_A net1443 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__179__A net1846 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_702 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__361__B net1367 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput930 net1170 vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__buf_8
Xoutput941 net1235 vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__buf_8
Xoutput952 net952 vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_5_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1705 mprj_logic1\[67\] vssd vssd vccd vccd net1705 sky130_fd_sc_hd__buf_6
Xwire1716 mprj_logic1\[58\] vssd vssd vccd vccd net1716 sky130_fd_sc_hd__buf_6
XFILLER_28_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1727 net1728 vssd vssd vccd vccd net1727 sky130_fd_sc_hd__buf_6
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__089__A la_data_in_mprj_bar\[106\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1738 net1739 vssd vssd vccd vccd net1738 sky130_fd_sc_hd__buf_6
Xwire1749 net1750 vssd vssd vccd vccd net1749 sky130_fd_sc_hd__buf_6
XTAP_3005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ mprj_logic1\[45\] net1356 vssd vssd vccd vccd net938 sky130_fd_sc_hd__and2_4
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__536__B mprj_logic1\[241\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_971 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_271_ net1775 net141 vssd vssd vccd vccd la_data_in_enable\[108\] sky130_fd_sc_hd__and2_4
XFILLER_13_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__552__A net338 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input375_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__271__B net141 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input69_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_607_ net1596 net1928 vssd vssd vccd vccd net731 sky130_fd_sc_hd__and2_4
XFILLER_45_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__B net2175 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_538_ net323 mprj_logic1\[243\] vssd vssd vccd vccd net782 sky130_fd_sc_hd__and2_4
XTAP_2893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output594_A net594 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_469_ net1607 net2133 net5 vssd vssd vccd vccd net464 sky130_fd_sc_hd__and3b_2
XFILLER_32_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output761_A net1030 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output859_A net859 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1392_A net1393 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__181__B net169 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1657_A net1658 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__356__B net1375 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B net1320 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3738 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput760 net1031 vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__buf_8
XFILLER_5_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput771 net771 vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__buf_8
XFILLER_40_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput782 net1018 vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__buf_8
XFILLER_8_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2203 net2204 vssd vssd vccd vccd net2203 sky130_fd_sc_hd__buf_6
Xoutput793 net793 vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__buf_8
XFILLER_47_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1502 net1503 vssd vssd vccd vccd net1502 sky130_fd_sc_hd__buf_6
Xwire1513 net1514 vssd vssd vccd vccd net1513 sky130_fd_sc_hd__buf_6
XFILLER_24_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1524 net1525 vssd vssd vccd vccd net1524 sky130_fd_sc_hd__buf_6
Xwire1535 net368 vssd vssd vccd vccd net1535 sky130_fd_sc_hd__buf_6
Xwire1546 net356 vssd vssd vccd vccd net1546 sky130_fd_sc_hd__buf_6
XFILLER_41_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1557 net34 vssd vssd vccd vccd net1557 sky130_fd_sc_hd__buf_4
Xwire1568 net317 vssd vssd vccd vccd net1568 sky130_fd_sc_hd__buf_6
XFILLER_38_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1579 net290 vssd vssd vccd vccd net1579 sky130_fd_sc_hd__buf_6
XANTENNA_input123_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2040_A net2041 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2138_A mprj_logic1\[171\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__A net333 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__266__B net136 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_323_ mprj_logic1\[28\] net1494 vssd vssd vccd vccd net857 sky130_fd_sc_hd__and2_4
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_B net1329 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_254_ net1802 net250 vssd vssd vccd vccd la_data_in_enable\[91\] sky130_fd_sc_hd__and2_4
XFILLER_32_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__282__A net1753 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_185_ net1839 net174 vssd vssd vccd vccd la_data_in_enable\[22\] sky130_fd_sc_hd__and2_4
XFILLER_45_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[4\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1140_A net546 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1238_A net1239 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1405_A net1406 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] la_data_in_enable\[21\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[21\] sky130_fd_sc_hd__nand2_1
XFILLER_50_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_B la_data_in_enable\[76\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__192__A net1828 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1774_A mprj_logic1\[439\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1941_A net1942 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__367__A net1692 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2088_A net2089 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2000 mprj_logic1\[280\] vssd vssd vccd vccd net2000 sky130_fd_sc_hd__buf_6
Xoutput590 net1136 vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__buf_8
XFILLER_44_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2011 mprj_logic1\[274\] vssd vssd vccd vccd net2011 sky130_fd_sc_hd__buf_6
XFILLER_21_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2022 mprj_logic1\[264\] vssd vssd vccd vccd net2022 sky130_fd_sc_hd__buf_6
XANTENNA_input240_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2033 mprj_logic1\[222\] vssd vssd vccd vccd net2033 sky130_fd_sc_hd__buf_6
XANTENNA_input338_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2044 mprj_logic1\[214\] vssd vssd vccd vccd net2044 sky130_fd_sc_hd__buf_6
XFILLER_21_2400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2055 net2056 vssd vssd vccd vccd net2055 sky130_fd_sc_hd__buf_6
XFILLER_40_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__440__A_N net1546 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1321 la_data_in_enable\[93\] vssd vssd vccd vccd net1321 sky130_fd_sc_hd__buf_6
Xwire2066 net2067 vssd vssd vccd vccd net2066 sky130_fd_sc_hd__buf_6
Xwire2077 net2078 vssd vssd vccd vccd net2077 sky130_fd_sc_hd__buf_6
XFILLER_8_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1332 la_data_in_enable\[80\] vssd vssd vccd vccd net1332 sky130_fd_sc_hd__buf_6
XFILLER_38_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1343 net458 vssd vssd vccd vccd net1343 sky130_fd_sc_hd__buf_6
Xwire2088 net2089 vssd vssd vccd vccd net2088 sky130_fd_sc_hd__buf_6
Xwire2099 net2100 vssd vssd vccd vccd net2099 sky130_fd_sc_hd__buf_6
Xwire1354 net1355 vssd vssd vccd vccd net1354 sky130_fd_sc_hd__buf_6
Xwire1365 net439 vssd vssd vccd vccd net1365 sky130_fd_sc_hd__buf_6
XFILLER_19_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1376 net430 vssd vssd vccd vccd net1376 sky130_fd_sc_hd__buf_6
XFILLER_38_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1387 net1388 vssd vssd vccd vccd net1387 sky130_fd_sc_hd__buf_6
Xwire1398 net1399 vssd vssd vccd vccd net1398 sky130_fd_sc_hd__buf_6
XANTENNA__277__A net1763 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_370 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_306_ net2200 net1485 vssd vssd vccd vccd net859 sky130_fd_sc_hd__and2_4
XFILLER_10_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_237_ mprj_logic1\[404\] net231 vssd vssd vccd vccd la_data_in_enable\[74\] sky130_fd_sc_hd__and2_4
XANTENNA__443__C net1630 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_168_ net1862 net215 vssd vssd vccd vccd la_data_in_enable\[5\] sky130_fd_sc_hd__and2_2
XFILLER_13_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output557_A net1139 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_099_ la_data_in_mprj_bar\[116\] vssd vssd vccd vccd net609 sky130_fd_sc_hd__inv_2
XANTENNA_wire1090_A net539 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1188_A net1189 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output724_A net724 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1355_A net447 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] la_data_in_enable\[69\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[69\] sky130_fd_sc_hd__nand2_4
XFILLER_39_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1522_A net1523 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__187__A net1835 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1891_A mprj_logic1\[324\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1989_A mprj_logic1\[285\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__463__A_N net381 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput307 la_oenb_mprj[27] vssd vssd vccd vccd net307 sky130_fd_sc_hd__buf_6
Xinput318 la_oenb_mprj[37] vssd vssd vccd vccd net318 sky130_fd_sc_hd__buf_6
Xinput329 la_oenb_mprj[47] vssd vssd vccd vccd net329 sky130_fd_sc_hd__buf_6
XFILLER_6_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__097__A net985 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_B net1312 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__544__B mprj_logic1\[249\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2003_A net2004 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input190_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input288_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_022_ la_data_in_mprj_bar\[39\] vssd vssd vccd vccd net651 sky130_fd_sc_hd__inv_2
XFILLER_6_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__A net1554 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input455_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input51_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1140 net546 vssd vssd vccd vccd net1140 sky130_fd_sc_hd__buf_6
XFILLER_1_3058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1151 net1152 vssd vssd vccd vccd net1151 sky130_fd_sc_hd__buf_6
Xwire1162 net1163 vssd vssd vccd vccd net1162 sky130_fd_sc_hd__buf_8
XFILLER_48_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1173 net930 vssd vssd vccd vccd net1173 sky130_fd_sc_hd__buf_6
Xwire1184 net1185 vssd vssd vccd vccd net1184 sky130_fd_sc_hd__buf_6
XFILLER_38_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1195 net1196 vssd vssd vccd vccd net1195 sky130_fd_sc_hd__buf_6
XANTENNA__438__C net1335 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__454__B net2156 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_B la_data_in_enable\[115\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_wire1103_A net526 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__486__A_N net1589 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output841_A net841 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output939_A net1241 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1472_A net1473 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1904_A mprj_logic1\[320\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[24\]_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[106\]_B la_data_in_enable\[106\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__364__B net1364 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput104 la_data_out_mprj[75] vssd vssd vccd vccd net104 sky130_fd_sc_hd__buf_6
XFILLER_40_2105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput115 la_data_out_mprj[85] vssd vssd vccd vccd net115 sky130_fd_sc_hd__buf_6
Xinput126 la_data_out_mprj[95] vssd vssd vccd vccd net126 sky130_fd_sc_hd__clkbuf_4
XTAP_4603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 la_iena_mprj[104] vssd vssd vccd vccd net137 sky130_fd_sc_hd__clkbuf_4
XTAP_4614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 la_iena_mprj[114] vssd vssd vccd vccd net148 sky130_fd_sc_hd__clkbuf_4
XTAP_4625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput159 la_iena_mprj[124] vssd vssd vccd vccd net159 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__539__B net2024 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[15\]_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_571_ net1543 net2007 vssd vssd vccd vccd net818 sky130_fd_sc_hd__and2_4
XTAP_3968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2120_A mprj_logic1\[182\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input203_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__555__A net1556 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__274__B net145 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input99_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__A net1735 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_005_ la_data_in_mprj_bar\[22\] vssd vssd vccd vccd net633 sky130_fd_sc_hd__clkinv_2
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__B net2169 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1053_A net719 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_958 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1220_A net1221 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output791_A net1049 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1318_A la_data_in_enable\[96\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1687_A mprj_logic1\[75\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1854_A net1855 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1909 net1910 vssd vssd vccd vccd net1909 sky130_fd_sc_hd__buf_6
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__359__B net1369 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 net1956 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2070_A net2071 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input153_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2168_A mprj_logic1\[155\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__269__B net139 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input320_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input418_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_623_ net1580 net1876 vssd vssd vccd vccd net748 sky130_fd_sc_hd__and2_4
XFILLER_22_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_554_ net340 mprj_logic1\[259\] vssd vssd vccd vccd net799 sky130_fd_sc_hd__and2_4
XTAP_3798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__285__A net1746 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_485_ net1590 net2099 net1611 vssd vssd vccd vccd net481 sky130_fd_sc_hd__and3b_4
XFILLER_31_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__451__C net1622 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output637_A net637 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1170_A net1171 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1268_A net1269 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output804_A net996 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1435_A net1436 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] la_data_in_enable\[51\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[51\] sky130_fd_sc_hd__nand2_4
XFILLER_40_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_714 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__195__A net1824 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1214 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1971_A mprj_logic1\[295\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput920 net1205 vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput931 net1166 vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__buf_8
Xoutput942 net1232 vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__buf_8
XFILLER_8_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput953 net2205 vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_9_3885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input6_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1706 net1707 vssd vssd vccd vccd net1706 sky130_fd_sc_hd__buf_6
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1717 mprj_logic1\[57\] vssd vssd vccd vccd net1717 sky130_fd_sc_hd__buf_6
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1728 mprj_logic1\[460\] vssd vssd vccd vccd net1728 sky130_fd_sc_hd__buf_6
XFILLER_3_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1739 mprj_logic1\[456\] vssd vssd vccd vccd net1739 sky130_fd_sc_hd__buf_6
XFILLER_25_2998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_270_ net1777 net140 vssd vssd vccd vccd la_data_in_enable\[107\] sky130_fd_sc_hd__and2_1
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__552__B mprj_logic1\[257\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input270_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input368_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_606_ net1597 net1931 vssd vssd vccd vccd net729 sky130_fd_sc_hd__and2_4
XTAP_3573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_91 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_537_ net1565 mprj_logic1\[242\] vssd vssd vccd vccd net781 sky130_fd_sc_hd__and2_4
XTAP_2872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__446__C net1627 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_468_ net1527 net2135 net130 vssd vssd vccd vccd net589 sky130_fd_sc_hd__and3b_4
XANTENNA_wire1016_A net1017 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output587_A net1069 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_399_ net1572 mprj_logic1\[104\] net55 vssd vssd vccd vccd net514 sky130_fd_sc_hd__and3b_2
XFILLER_31_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__B mprj_logic1\[167\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output754_A net1036 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1385_A net1386 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output921_A net1202 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] net1317 vssd vssd vccd vccd la_data_in_mprj_bar\[99\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_29_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1817_A mprj_logic1\[37\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__372__B net1682 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2980 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[7\]_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput750 net1040 vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__buf_8
Xoutput761 net1030 vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__buf_8
Xoutput772 net772 vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__buf_8
XFILLER_5_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput783 net1016 vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__buf_8
XFILLER_40_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2204 mprj_logic1\[0\] vssd vssd vccd vccd net2204 sky130_fd_sc_hd__buf_6
Xoutput794 net1007 vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__buf_8
XFILLER_5_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1503 net1504 vssd vssd vccd vccd net1503 sky130_fd_sc_hd__buf_6
XFILLER_24_1015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1514 net392 vssd vssd vccd vccd net1514 sky130_fd_sc_hd__buf_6
XFILLER_43_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1525 net1526 vssd vssd vccd vccd net1525 sky130_fd_sc_hd__buf_6
XFILLER_24_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1536 net367 vssd vssd vccd vccd net1536 sky130_fd_sc_hd__buf_6
XFILLER_1_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1547 net355 vssd vssd vccd vccd net1547 sky130_fd_sc_hd__buf_6
XFILLER_24_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1558 net334 vssd vssd vccd vccd net1558 sky130_fd_sc_hd__buf_6
XFILLER_3_3292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1569 net316 vssd vssd vccd vccd net1569 sky130_fd_sc_hd__buf_6
XFILLER_38_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__B mprj_logic1\[252\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input116_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2033_A mprj_logic1\[222\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ mprj_logic1\[27\] net1498 vssd vssd vccd vccd net856 sky130_fd_sc_hd__and2_4
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2200_A mprj_logic1\[11\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__563__A net1551 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_253_ mprj_logic1\[420\] net249 vssd vssd vccd vccd la_data_in_enable\[90\] sky130_fd_sc_hd__and2_4
XFILLER_14_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input81_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_184_ net1840 net173 vssd vssd vccd vccd la_data_in_enable\[21\] sky130_fd_sc_hd__and2_1
XFILLER_52_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output502_A net1144 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__457__B net2146 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1133_A net1134 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1300_A net1301 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output871_A net871 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] la_data_in_enable\[14\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[14\] sky130_fd_sc_hd__nand2_4
XFILLER_31_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[27\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_33_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__192__B net181 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1767_A net1768 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1934_A net1935 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] la_data_in_enable\[125\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[125\] sky130_fd_sc_hd__nand2_4
XFILLER_9_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__367__B net1359 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__A_N net303 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput580 net1076 vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__buf_8
XFILLER_40_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2001 net2002 vssd vssd vccd vccd net2001 sky130_fd_sc_hd__buf_6
XFILLER_25_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput591 net591 vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_8
Xwire2012 net2013 vssd vssd vccd vccd net2012 sky130_fd_sc_hd__buf_6
XFILLER_27_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2023 mprj_logic1\[251\] vssd vssd vccd vccd net2023 sky130_fd_sc_hd__buf_4
XFILLER_8_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2034 mprj_logic1\[221\] vssd vssd vccd vccd net2034 sky130_fd_sc_hd__buf_6
Xwire1300 net1301 vssd vssd vccd vccd net1300 sky130_fd_sc_hd__buf_6
Xwire2045 net2046 vssd vssd vccd vccd net2045 sky130_fd_sc_hd__buf_6
Xwire2056 mprj_logic1\[207\] vssd vssd vccd vccd net2056 sky130_fd_sc_hd__buf_6
XFILLER_21_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1322 la_data_in_enable\[92\] vssd vssd vccd vccd net1322 sky130_fd_sc_hd__buf_6
XFILLER_5_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2067 net2068 vssd vssd vccd vccd net2067 sky130_fd_sc_hd__buf_6
XANTENNA_wire2150_A net2151 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input233_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2078 mprj_logic1\[198\] vssd vssd vccd vccd net2078 sky130_fd_sc_hd__buf_6
Xwire1333 la_data_in_enable\[79\] vssd vssd vccd vccd net1333 sky130_fd_sc_hd__buf_6
XFILLER_5_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1344 net1345 vssd vssd vccd vccd net1344 sky130_fd_sc_hd__buf_6
Xwire2089 net2090 vssd vssd vccd vccd net2089 sky130_fd_sc_hd__buf_6
XFILLER_38_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__558__A net345 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1355 net447 vssd vssd vccd vccd net1355 sky130_fd_sc_hd__buf_6
Xwire1366 net438 vssd vssd vccd vccd net1366 sky130_fd_sc_hd__buf_6
XFILLER_21_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1377 net429 vssd vssd vccd vccd net1377 sky130_fd_sc_hd__buf_6
XFILLER_35_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1388 net423 vssd vssd vccd vccd net1388 sky130_fd_sc_hd__buf_6
XFILLER_38_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1399 net1400 vssd vssd vccd vccd net1399 sky130_fd_sc_hd__buf_6
XANTENNA_input400_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__277__B net148 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__293__A net1726 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ net2201 net1522 vssd vssd vccd vccd net848 sky130_fd_sc_hd__and2_2
XFILLER_15_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_236_ mprj_logic1\[403\] net230 vssd vssd vccd vccd la_data_in_enable\[73\] sky130_fd_sc_hd__and2_4
XFILLER_10_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_167_ net1863 net204 vssd vssd vccd vccd la_data_in_enable\[4\] sky130_fd_sc_hd__and2_1
XFILLER_6_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_098_ net984 vssd vssd vccd vccd net608 sky130_fd_sc_hd__inv_2
XFILLER_26_3024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1083_A net544 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output717_A net717 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1250_A net924 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1348_A net1349 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__187__B net1614 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1515_A net1516 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1884_A net1885 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire968_A la_data_in_mprj_bar\[89\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput308 la_oenb_mprj[28] vssd vssd vccd vccd net308 sky130_fd_sc_hd__buf_4
XFILLER_9_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput319 la_oenb_mprj[38] vssd vssd vccd vccd net319 sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2859 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_021_ la_data_in_mprj_bar\[38\] vssd vssd vccd vccd net650 sky130_fd_sc_hd__inv_2
XFILLER_10_2124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input183_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__B net2021 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input350_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input448_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input44_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1130 net496 vssd vssd vccd vccd net1130 sky130_fd_sc_hd__buf_6
XFILLER_40_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__288__A net1740 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1141 net535 vssd vssd vccd vccd net1141 sky130_fd_sc_hd__buf_6
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1152 net1153 vssd vssd vccd vccd net1152 sky130_fd_sc_hd__buf_6
Xwire1163 net1164 vssd vssd vccd vccd net1163 sky130_fd_sc_hd__buf_6
XFILLER_38_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1174 net1175 vssd vssd vccd vccd net1174 sky130_fd_sc_hd__buf_8
Xwire1185 net927 vssd vssd vccd vccd net1185 sky130_fd_sc_hd__buf_6
XFILLER_34_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1196 net1197 vssd vssd vccd vccd net1196 sky130_fd_sc_hd__buf_6
XFILLER_35_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__454__C net1619 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_219_ mprj_logic1\[386\] net211 vssd vssd vccd vccd la_data_in_enable\[56\] sky130_fd_sc_hd__and2_2
XFILLER_32_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1298_A net945 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__470__B net2132 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output834_A net995 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1465_A net1466 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] la_data_in_enable\[81\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[81\] sky130_fd_sc_hd__nand2_1
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__198__A mprj_logic1\[365\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_606 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_672 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__430__A_N net345 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__380__B net1663 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput105 la_data_out_mprj[76] vssd vssd vccd vccd net105 sky130_fd_sc_hd__buf_6
Xinput116 la_data_out_mprj[86] vssd vssd vccd vccd net116 sky130_fd_sc_hd__buf_6
XFILLER_44_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput127 la_data_out_mprj[96] vssd vssd vccd vccd net127 sky130_fd_sc_hd__clkbuf_4
XTAP_4604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 la_iena_mprj[105] vssd vssd vccd vccd net138 sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput149 la_iena_mprj[115] vssd vssd vccd vccd net149 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[15\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_570_ net1544 net2009 vssd vssd vccd vccd net817 sky130_fd_sc_hd__and2_4
XTAP_3958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__555__B mprj_logic1\[260\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2113_A net2114 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input398_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__571__A net1543 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_004_ la_data_in_mprj_bar\[21\] vssd vssd vccd vccd net632 sky130_fd_sc_hd__inv_2
XFILLER_46_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__B net162 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__449__C net1624 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1046_A net824 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__465__B net2139 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1213_A net918 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__453__A_N net1533 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output784_A net784 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output951_A net1723 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1847_A net1848 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__375__B net1674 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2063_A mprj_logic1\[203\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input146_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_622_ net1581 net1879 vssd vssd vccd vccd net747 sky130_fd_sc_hd__and2_4
XFILLER_22_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input313_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__476__A_N net1600 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__566__A net1548 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_553_ net339 mprj_logic1\[258\] vssd vssd vccd vccd net798 sky130_fd_sc_hd__and2_2
XTAP_3788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__285__B net157 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_484_ net1591 net2102 net21 vssd vssd vccd vccd net480 sky130_fd_sc_hd__and3b_4
XFILLER_35_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output532_A net1097 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1163_A net1164 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1330_A la_data_in_enable\[84\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1428_A net1429 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] la_data_in_enable\[44\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[44\] sky130_fd_sc_hd__nand2_2
XFILLER_18_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1797_A mprj_logic1\[426\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1964_A mprj_logic1\[299\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput910 net910 vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_8
Xoutput921 net1202 vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__buf_8
Xoutput932 net1162 vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__buf_8
Xoutput943 net1229 vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_4379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] la_data_in_enable\[6\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[6\] sky130_fd_sc_hd__nand2_2
XFILLER_25_2900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput954 net954 vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_3_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1707 mprj_logic1\[66\] vssd vssd vccd vccd net1707 sky130_fd_sc_hd__buf_6
XFILLER_3_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1718 mprj_logic1\[56\] vssd vssd vccd vccd net1718 sky130_fd_sc_hd__buf_6
XFILLER_41_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1729 net1730 vssd vssd vccd vccd net1729 sky130_fd_sc_hd__buf_6
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input263_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2180_A net2181 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input430_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__296__A mprj_logic1\[1\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_605_ net1599 net1934 vssd vssd vccd vccd net728 sky130_fd_sc_hd__and2_2
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_536_ net320 mprj_logic1\[241\] vssd vssd vccd vccd net779 sky130_fd_sc_hd__and2_4
XFILLER_15_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_467_ net1528 net2136 net129 vssd vssd vccd vccd net588 sky130_fd_sc_hd__and3b_4
XFILLER_14_962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_398_ net1574 mprj_logic1\[103\] net53 vssd vssd vccd vccd net512 sky130_fd_sc_hd__and3b_4
XANTENNA_output482_A net482 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1009_A net1010 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__462__C net124 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output747_A net747 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1280_A net1281 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1378_A net428 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output914_A net1223 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3818 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1712_A mprj_logic1\[61\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[7\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput740 net740 vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__buf_8
XFILLER_5_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput751 net1039 vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput762 net1029 vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__buf_8
XFILLER_5_3514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput773 net1024 vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__buf_8
Xoutput784 net784 vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__buf_8
XFILLER_40_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2205 net2206 vssd vssd vccd vccd net2205 sky130_fd_sc_hd__buf_6
Xoutput795 net1005 vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__buf_8
XFILLER_5_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1504 net395 vssd vssd vccd vccd net1504 sky130_fd_sc_hd__buf_6
XFILLER_41_2042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1515 net1516 vssd vssd vccd vccd net1515 sky130_fd_sc_hd__buf_6
Xwire1526 net388 vssd vssd vccd vccd net1526 sky130_fd_sc_hd__buf_6
XFILLER_5_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1537 net366 vssd vssd vccd vccd net1537 sky130_fd_sc_hd__buf_6
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[7\]_B la_data_in_enable\[7\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1548 net353 vssd vssd vccd vccd net1548 sky130_fd_sc_hd__buf_6
Xwire1559 net330 vssd vssd vccd vccd net1559 sky130_fd_sc_hd__buf_6
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2026_A mprj_logic1\[236\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input109_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ mprj_logic1\[26\] net1501 vssd vssd vccd vccd net855 sky130_fd_sc_hd__and2_2
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_252_ mprj_logic1\[419\] net247 vssd vssd vccd vccd la_data_in_enable\[89\] sky130_fd_sc_hd__and2_4
XANTENNA__563__B net2018 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_183_ net1841 net172 vssd vssd vccd vccd la_data_in_enable\[20\] sky130_fd_sc_hd__and2_1
XANTENNA_input380_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input74_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__457__C net1616 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1126_A net500 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_519_ net302 net2031 vssd vssd vccd vccd net761 sky130_fd_sc_hd__and2_4
XFILLER_35_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__473__B net2126 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output864_A net864 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1495_A net1496 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1662_A mprj_logic1\[86\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1927_A mprj_logic1\[313\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] la_data_in_enable\[118\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[118\] sky130_fd_sc_hd__nand2_2
XFILLER_3_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__383__B net1657 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput570 net570 vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__buf_8
XFILLER_44_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput581 net1075 vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__buf_8
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2002 mprj_logic1\[279\] vssd vssd vccd vccd net2002 sky130_fd_sc_hd__buf_6
XFILLER_40_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput592 net592 vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_8
XFILLER_5_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2013 mprj_logic1\[273\] vssd vssd vccd vccd net2013 sky130_fd_sc_hd__buf_6
Xwire2024 mprj_logic1\[244\] vssd vssd vccd vccd net2024 sky130_fd_sc_hd__buf_4
XFILLER_43_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2035 mprj_logic1\[220\] vssd vssd vccd vccd net2035 sky130_fd_sc_hd__buf_6
Xwire1301 net1302 vssd vssd vccd vccd net1301 sky130_fd_sc_hd__buf_6
XFILLER_8_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2046 mprj_logic1\[213\] vssd vssd vccd vccd net2046 sky130_fd_sc_hd__buf_6
XFILLER_21_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1312 la_data_in_enable\[124\] vssd vssd vccd vccd net1312 sky130_fd_sc_hd__buf_8
Xwire2057 mprj_logic1\[206\] vssd vssd vccd vccd net2057 sky130_fd_sc_hd__buf_6
Xwire2068 mprj_logic1\[201\] vssd vssd vccd vccd net2068 sky130_fd_sc_hd__buf_6
Xwire1323 la_data_in_enable\[91\] vssd vssd vccd vccd net1323 sky130_fd_sc_hd__buf_6
XFILLER_43_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1334 net99 vssd vssd vccd vccd net1334 sky130_fd_sc_hd__buf_6
Xwire2079 net2080 vssd vssd vccd vccd net2079 sky130_fd_sc_hd__buf_6
XFILLER_19_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1345 net452 vssd vssd vccd vccd net1345 sky130_fd_sc_hd__buf_6
XANTENNA__558__B mprj_logic1\[263\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1356 net1357 vssd vssd vccd vccd net1356 sky130_fd_sc_hd__buf_6
XFILLER_5_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2143_A mprj_logic1\[165\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input226_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1367 net437 vssd vssd vccd vccd net1367 sky130_fd_sc_hd__buf_6
Xwire1378 net428 vssd vssd vccd vccd net1378 sky130_fd_sc_hd__buf_6
Xwire1389 net1390 vssd vssd vccd vccd net1389 sky130_fd_sc_hd__buf_6
XFILLER_34_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__574__A net1540 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__293__B net462 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_304_ net1634 net457 vssd vssd vccd vccd net948 sky130_fd_sc_hd__and2_4
XFILLER_10_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_235_ mprj_logic1\[402\] net229 vssd vssd vccd vccd la_data_in_enable\[72\] sky130_fd_sc_hd__and2_4
XFILLER_32_2553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_166_ net1865 net193 vssd vssd vccd vccd la_data_in_enable\[3\] sky130_fd_sc_hd__and2_1
XFILLER_49_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_097_ net985 vssd vssd vccd vccd net607 sky130_fd_sc_hd__clkinv_2
XFILLER_45_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1076_A net580 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__468__B net2135 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1890 net1891 vssd vssd vccd vccd net1890 sky130_fd_sc_hd__buf_6
XFILLER_37_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1410_A net1411 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1508_A net394 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_190 net1818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1638 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1877_A net1878 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput309 la_oenb_mprj[29] vssd vssd vccd vccd net309 sky130_fd_sc_hd__buf_6
XFILLER_29_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__B net1668 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_16_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_020_ la_data_in_mprj_bar\[37\] vssd vssd vccd vccd net649 sky130_fd_sc_hd__clkinv_2
XFILLER_14_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2093_A mprj_logic1\[193\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input176_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input343_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__569__A net1545 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input37_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1120 net507 vssd vssd vccd vccd net1120 sky130_fd_sc_hd__buf_6
XFILLER_19_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1131 net495 vssd vssd vccd vccd net1131 sky130_fd_sc_hd__buf_6
XFILLER_25_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__288__B net160 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1142 net524 vssd vssd vccd vccd net1142 sky130_fd_sc_hd__buf_6
XFILLER_40_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1153 net936 vssd vssd vccd vccd net1153 sky130_fd_sc_hd__buf_6
Xwire1164 net1165 vssd vssd vccd vccd net1164 sky130_fd_sc_hd__buf_6
XFILLER_5_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1175 net1176 vssd vssd vccd vccd net1175 sky130_fd_sc_hd__buf_6
XFILLER_5_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1186 net1187 vssd vssd vccd vccd net1186 sky130_fd_sc_hd__buf_8
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1197 net923 vssd vssd vccd vccd net1197 sky130_fd_sc_hd__buf_6
XFILLER_34_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_218_ mprj_logic1\[385\] net210 vssd vssd vccd vccd la_data_in_enable\[55\] sky130_fd_sc_hd__and2_2
XFILLER_45_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output562_A net562 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_149_ la_data_in_mprj_bar\[2\] vssd vssd vccd vccd net641 sky130_fd_sc_hd__inv_2
XFILLER_7_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__C net6 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output827_A net827 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__382__A_N net292 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1360_A net1361 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1458_A net1459 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] la_data_in_enable\[74\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[74\] sky130_fd_sc_hd__nand2_4
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1625_A net108 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1994_A net1995 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_684 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__380__C net26 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput106 la_data_out_mprj[77] vssd vssd vccd vccd net106 sky130_fd_sc_hd__buf_6
XFILLER_41_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput117 la_data_out_mprj[87] vssd vssd vccd vccd net117 sky130_fd_sc_hd__buf_6
XFILLER_2_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput128 la_data_out_mprj[97] vssd vssd vccd vccd net128 sky130_fd_sc_hd__clkbuf_4
XTAP_4605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput139 la_iena_mprj[106] vssd vssd vccd vccd net139 sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2106_A net2107 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1546 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input293_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__571__B net2007 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_90 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_003_ la_data_in_mprj_bar\[20\] vssd vssd vccd vccd net631 sky130_fd_sc_hd__inv_2
XFILLER_29_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input460_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__299__A mprj_logic1\[4\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1039_A net751 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1206_A net1207 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output777_A net777 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__481__B net2110 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output944_A net1226 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1742_A net1743 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__002__A la_data_in_mprj_bar\[19\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] la_data_in_enable\[100\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[100\] sky130_fd_sc_hd__nand2_1
XFILLER_39_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__391__B net1641 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input139_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2056_A mprj_logic1\[207\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_621_ net1582 net1883 vssd vssd vccd vccd net746 sky130_fd_sc_hd__and2_4
XTAP_4468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_552_ net338 mprj_logic1\[257\] vssd vssd vccd vccd net797 sky130_fd_sc_hd__and2_4
XANTENNA__566__B net2015 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input306_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_483_ net1592 net2105 net20 vssd vssd vccd vccd net479 sky130_fd_sc_hd__and3b_4
XFILLER_44_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__582__A net1532 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output525_A net1104 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1156_A net1157 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__420__A_N net334 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__476__B net2121 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1323_A la_data_in_enable\[91\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output894_A net894 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] la_data_in_enable\[37\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[37\] sky130_fd_sc_hd__nand2_4
XFILLER_23_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1692_A net1693 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1957_A net1958 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput900 net900 vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_8
XFILLER_9_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput911 net911 vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_8
XFILLER_25_4347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput922 net1198 vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__buf_8
Xoutput933 net1158 vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__buf_8
Xoutput944 net1226 vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__buf_8
XFILLER_28_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput955 net1307 vssd vssd vccd vccd user_clock sky130_fd_sc_hd__buf_8
XFILLER_45_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[30\]_B la_data_in_enable\[30\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1708 mprj_logic1\[65\] vssd vssd vccd vccd net1708 sky130_fd_sc_hd__buf_6
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1719 mprj_logic1\[55\] vssd vssd vccd vccd net1719 sky130_fd_sc_hd__buf_4
XFILLER_45_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__386__B net1650 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B la_data_in_enable\[97\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2173_A net2174 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input256_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__443__A_N net1543 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input423_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__577__A net1537 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_604_ net1600 net1937 vssd vssd vccd vccd net727 sky130_fd_sc_hd__and2_4
XTAP_4298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_716 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_535_ net319 net2025 vssd vssd vccd vccd net778 sky130_fd_sc_hd__and2_1
XFILLER_35_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_B net1326 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_466_ net384 net2137 net128 vssd vssd vccd vccd net587 sky130_fd_sc_hd__and3b_4
XFILLER_53_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_397_ net308 mprj_logic1\[102\] net52 vssd vssd vccd vccd net511 sky130_fd_sc_hd__and3b_4
XFILLER_35_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output475_A net1056 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output642_A net642 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1273_A net849 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1440_A net1441 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1538_A net364 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B net1333 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__466__A_N net384 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput730 net1042 vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__buf_8
XFILLER_9_3651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput741 net1041 vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__buf_8
XFILLER_25_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput752 net1038 vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__buf_8
XFILLER_47_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput763 net1028 vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__buf_8
Xoutput774 net1022 vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__buf_8
XFILLER_5_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput785 net1015 vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__buf_8
Xwire2206 net2207 vssd vssd vccd vccd net2206 sky130_fd_sc_hd__buf_6
XFILLER_25_3476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput796 net796 vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__buf_8
XFILLER_48_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1505 net1506 vssd vssd vccd vccd net1505 sky130_fd_sc_hd__buf_6
Xwire1516 net1517 vssd vssd vccd vccd net1516 sky130_fd_sc_hd__buf_6
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2054 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1527 net386 vssd vssd vccd vccd net1527 sky130_fd_sc_hd__buf_6
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1538 net364 vssd vssd vccd vccd net1538 sky130_fd_sc_hd__buf_6
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1549 net352 vssd vssd vccd vccd net1549 sky130_fd_sc_hd__buf_6
XFILLER_38_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ mprj_logic1\[25\] net1505 vssd vssd vccd vccd net854 sky130_fd_sc_hd__and2_4
XFILLER_42_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2019_A mprj_logic1\[267\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_251_ net1804 net246 vssd vssd vccd vccd la_data_in_enable\[88\] sky130_fd_sc_hd__and2_4
XFILLER_32_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_182_ net1843 net170 vssd vssd vccd vccd la_data_in_enable\[19\] sky130_fd_sc_hd__and2_2
XFILLER_49_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input373_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input67_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__100__A net983 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_518_ net301 net2032 vssd vssd vccd vccd net760 sky130_fd_sc_hd__and2_4
XTAP_2682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output592_A net592 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1119_A net508 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_449_ net1537 net2169 net1624 vssd vssd vccd vccd net569 sky130_fd_sc_hd__and3b_4
XFILLER_15_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__489__A_N net1586 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output857_A net857 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1488_A net1489 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1655_A net1656 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__383__C net37 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2590 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput560 net560 vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__buf_8
XFILLER_40_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput571 net571 vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__buf_8
XFILLER_43_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput582 net1074 vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__buf_8
XFILLER_44_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2003 net2004 vssd vssd vccd vccd net2003 sky130_fd_sc_hd__buf_6
Xoutput593 net593 vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_8
XFILLER_8_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2014 mprj_logic1\[272\] vssd vssd vccd vccd net2014 sky130_fd_sc_hd__buf_6
XFILLER_47_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2025 mprj_logic1\[240\] vssd vssd vccd vccd net2025 sky130_fd_sc_hd__buf_6
XFILLER_47_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2036 mprj_logic1\[219\] vssd vssd vccd vccd net2036 sky130_fd_sc_hd__buf_6
XFILLER_43_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2047 net2048 vssd vssd vccd vccd net2047 sky130_fd_sc_hd__buf_6
XFILLER_25_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1302 net950 vssd vssd vccd vccd net1302 sky130_fd_sc_hd__buf_6
XFILLER_8_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2058 net2059 vssd vssd vccd vccd net2058 sky130_fd_sc_hd__buf_6
Xwire1313 la_data_in_enable\[123\] vssd vssd vccd vccd net1313 sky130_fd_sc_hd__buf_6
Xwire2069 net2070 vssd vssd vccd vccd net2069 sky130_fd_sc_hd__buf_6
XFILLER_21_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1324 la_data_in_enable\[90\] vssd vssd vccd vccd net1324 sky130_fd_sc_hd__buf_8
XFILLER_25_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1335 net97 vssd vssd vccd vccd net1335 sky130_fd_sc_hd__buf_6
XFILLER_21_2436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1346 net1347 vssd vssd vccd vccd net1346 sky130_fd_sc_hd__buf_6
XFILLER_21_2447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1357 net446 vssd vssd vccd vccd net1357 sky130_fd_sc_hd__buf_6
Xwire1368 net436 vssd vssd vccd vccd net1368 sky130_fd_sc_hd__buf_6
Xwire1379 net1380 vssd vssd vccd vccd net1379 sky130_fd_sc_hd__buf_6
XFILLER_28_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input121_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input219_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2136_A mprj_logic1\[172\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__574__B net2001 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_B la_data_in_enable\[127\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_303_ net1654 net456 vssd vssd vccd vccd net947 sky130_fd_sc_hd__and2_1
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_234_ mprj_logic1\[401\] net228 vssd vssd vccd vccd la_data_in_enable\[71\] sky130_fd_sc_hd__and2_4
XFILLER_7_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__590__A net380 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_165_ net1867 net182 vssd vssd vccd vccd la_data_in_enable\[2\] sky130_fd_sc_hd__and2_1
XFILLER_6_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[2\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_32_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_096_ net986 vssd vssd vccd vccd net606 sky130_fd_sc_hd__inv_2
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_powergood_check_mprj_vdd_logic1 net952 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__468__C net130 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output605_A net605 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1880 net1881 vssd vssd vccd vccd net1880 sky130_fd_sc_hd__buf_6
XANTENNA_wire1236_A net1237 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1891 mprj_logic1\[324\] vssd vssd vccd vccd net1891 sky130_fd_sc_hd__buf_6
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__484__B net2102 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_B la_data_in_enable\[118\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1403_A net1404 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_180 net1811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_191 net1818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1772_A mprj_logic1\[440\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4322 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__005__A la_data_in_mprj_bar\[22\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[27\]_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__C net131 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__B net1635 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[109\]_B la_data_in_enable\[109\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_24_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2086_A net2087 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input169_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__569__B net2010 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input336_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[18\]_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1110 net518 vssd vssd vccd vccd net1110 sky130_fd_sc_hd__buf_6
XFILLER_25_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1121 net506 vssd vssd vccd vccd net1121 sky130_fd_sc_hd__buf_6
Xwire1132 net494 vssd vssd vccd vccd net1132 sky130_fd_sc_hd__buf_6
XFILLER_5_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1143 net513 vssd vssd vccd vccd net1143 sky130_fd_sc_hd__buf_6
Xwire1154 net1155 vssd vssd vccd vccd net1154 sky130_fd_sc_hd__buf_8
XFILLER_1_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1165 net932 vssd vssd vccd vccd net1165 sky130_fd_sc_hd__buf_6
Xwire1176 net1177 vssd vssd vccd vccd net1176 sky130_fd_sc_hd__buf_6
XFILLER_38_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1187 net1188 vssd vssd vccd vccd net1187 sky130_fd_sc_hd__buf_6
XFILLER_5_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1198 net1199 vssd vssd vccd vccd net1198 sky130_fd_sc_hd__buf_8
XFILLER_53_3907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__585__A net1529 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_217_ mprj_logic1\[384\] net209 vssd vssd vccd vccd la_data_in_enable\[54\] sky130_fd_sc_hd__and2_1
XFILLER_10_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_148_ la_data_in_mprj_bar\[1\] vssd vssd vccd vccd net630 sky130_fd_sc_hd__inv_2
XFILLER_13_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output555_A net555 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_079_ la_data_in_mprj_bar\[96\] vssd vssd vccd vccd net714 sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1186_A net1187 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output722_A net722 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__479__B net2115 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1353_A net448 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] la_data_in_enable\[67\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[67\] sky130_fd_sc_hd__nand2_4
XFILLER_1_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1520_A net1521 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1618_A net116 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1987_A mprj_logic1\[286\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire973_A la_data_in_mprj_bar\[84\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput107 la_data_out_mprj[78] vssd vssd vccd vccd net107 sky130_fd_sc_hd__buf_6
XFILLER_22_3232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput118 la_data_out_mprj[88] vssd vssd vccd vccd net118 sky130_fd_sc_hd__buf_6
XANTENNA__389__B net1645 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput129 la_data_out_mprj[98] vssd vssd vccd vccd net129 sky130_fd_sc_hd__clkbuf_4
XTAP_4606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2001_A net2002 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input286_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_80 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_002_ la_data_in_mprj_bar\[19\] vssd vssd vccd vccd net629 sky130_fd_sc_hd__inv_2
XFILLER_11_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_91 mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input453_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__299__B net1342 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1101_A net528 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__481__C net18 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output937_A net1146 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1470_A net1471 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1568_A net317 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1735_A net1736 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1902_A net1903 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_620_ net1583 net1886 vssd vssd vccd vccd net745 sky130_fd_sc_hd__and2_4
XFILLER_22_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2049_A net2050 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_551_ net337 mprj_logic1\[256\] vssd vssd vccd vccd net796 sky130_fd_sc_hd__and2_4
XTAP_3768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input201_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_482_ net1593 net2108 net19 vssd vssd vccd vccd net478 sky130_fd_sc_hd__and3b_4
XFILLER_32_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__372__A_N net321 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__582__B net1984 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input97_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__103__A la_data_in_mprj_bar\[120\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3758 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output518_A net1110 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput460 user_irq_ena[0] vssd vssd vccd vccd net460 sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1051_A net769 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3632 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__492__B net2079 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1685_A mprj_logic1\[76\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput901 net901 vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_8
Xoutput912 net912 vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_8
XANTENNA_wire1852_A net1853 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput923 net1194 vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_28_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput934 net1154 vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput945 net1294 vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__buf_8
Xoutput956 net956 vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__buf_8
XFILLER_45_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1709 mprj_logic1\[64\] vssd vssd vccd vccd net1709 sky130_fd_sc_hd__buf_6
XFILLER_25_2968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__386__C net40 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__395__A_N net306 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input151_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2166_A mprj_logic1\[156\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input249_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__577__B net1994 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input416_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_603_ net1601 net1939 vssd vssd vccd vccd net726 sky130_fd_sc_hd__and2_4
XTAP_4288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_534_ net1567 mprj_logic1\[239\] vssd vssd vccd vccd net777 sky130_fd_sc_hd__and2_4
XFILLER_15_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__A net383 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ net383 net2139 net127 vssd vssd vccd vccd net586 sky130_fd_sc_hd__and3b_4
XTAP_2897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_396_ net1575 mprj_logic1\[101\] net51 vssd vssd vccd vccd net510 sky130_fd_sc_hd__and3b_4
XFILLER_13_3551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output468_A net1062 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1099_A net530 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output635_A net635 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1266_A net1267 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output802_A net1048 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__487__B net2094 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1433_A net1434 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput290 la_oenb_mprj[127] vssd vssd vccd vccd net290 sky130_fd_sc_hd__buf_6
XFILLER_3_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__008__A la_data_in_mprj_bar\[25\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput720 net720 vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__buf_8
XFILLER_47_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput731 net731 vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__buf_8
Xoutput742 net742 vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__buf_8
XFILLER_9_3663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput753 net1037 vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__buf_8
XFILLER_43_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput764 net1027 vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__buf_8
XFILLER_47_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput775 net775 vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__buf_8
XFILLER_9_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput786 net1013 vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__buf_8
Xwire2207 net2208 vssd vssd vccd vccd net2207 sky130_fd_sc_hd__buf_6
Xoutput797 net1004 vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__buf_8
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1506 net1507 vssd vssd vccd vccd net1506 sky130_fd_sc_hd__buf_6
XFILLER_24_1018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1517 net391 vssd vssd vccd vccd net1517 sky130_fd_sc_hd__buf_6
XFILLER_24_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1528 net385 vssd vssd vccd vccd net1528 sky130_fd_sc_hd__buf_6
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1539 net363 vssd vssd vccd vccd net1539 sky130_fd_sc_hd__buf_8
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__397__B mprj_logic1\[102\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_250_ net1805 net245 vssd vssd vccd vccd la_data_in_enable\[87\] sky130_fd_sc_hd__and2_4
XFILLER_36_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_181_ net1844 net169 vssd vssd vccd vccd la_data_in_enable\[18\] sky130_fd_sc_hd__and2_1
XFILLER_52_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input199_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__A_N net323 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input366_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_gates\[1\] user_irq_core[1] user_irq_enable\[1\] vssd vssd vccd vccd user_irq_bar\[1\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_8_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__588__A net378 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_517_ net300 net2033 vssd vssd vccd vccd net759 sky130_fd_sc_hd__and2_4
XTAP_2672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ net1538 net2171 net1625 vssd vssd vccd vccd net567 sky130_fd_sc_hd__and3b_4
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output585_A net1071 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3370 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_379_ net271 net1666 net15 vssd vssd vccd vccd net474 sky130_fd_sc_hd__and3b_4
XFILLER_35_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output752_A net1038 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1383_A net1384 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] la_data_in_enable\[97\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[97\] sky130_fd_sc_hd__nand2_8
XFILLER_6_3825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1648_A net1649 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__498__A net299 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__A_N net1553 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput550 net550 vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__buf_8
Xoutput561 net561 vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__buf_8
XFILLER_27_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput572 net572 vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__buf_8
XFILLER_47_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput583 net1073 vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__buf_8
Xwire2004 mprj_logic1\[278\] vssd vssd vccd vccd net2004 sky130_fd_sc_hd__buf_6
Xoutput594 net594 vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_8
XFILLER_5_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2015 mprj_logic1\[271\] vssd vssd vccd vccd net2015 sky130_fd_sc_hd__buf_6
XFILLER_8_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2026 mprj_logic1\[236\] vssd vssd vccd vccd net2026 sky130_fd_sc_hd__buf_6
Xwire2037 net2038 vssd vssd vccd vccd net2037 sky130_fd_sc_hd__buf_6
XFILLER_25_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1303 net1304 vssd vssd vccd vccd net1303 sky130_fd_sc_hd__buf_6
Xwire2048 mprj_logic1\[212\] vssd vssd vccd vccd net2048 sky130_fd_sc_hd__buf_6
XFILLER_43_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__201__A mprj_logic1\[368\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2059 mprj_logic1\[205\] vssd vssd vccd vccd net2059 sky130_fd_sc_hd__buf_6
XFILLER_21_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1314 la_data_in_enable\[114\] vssd vssd vccd vccd net1314 sky130_fd_sc_hd__buf_6
Xwire1325 la_data_in_enable\[89\] vssd vssd vccd vccd net1325 sky130_fd_sc_hd__buf_8
XFILLER_25_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1336 net96 vssd vssd vccd vccd net1336 sky130_fd_sc_hd__buf_6
Xwire1347 net451 vssd vssd vccd vccd net1347 sky130_fd_sc_hd__buf_6
XFILLER_3_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1358 net445 vssd vssd vccd vccd net1358 sky130_fd_sc_hd__buf_6
Xwire1369 net435 vssd vssd vccd vccd net1369 sky130_fd_sc_hd__buf_6
XFILLER_38_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2031_A mprj_logic1\[224\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input114_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2129_A mprj_logic1\[177\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ net1676 net455 vssd vssd vccd vccd net946 sky130_fd_sc_hd__and2_2
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_233_ net1810 net227 vssd vssd vccd vccd la_data_in_enable\[70\] sky130_fd_sc_hd__and2_2
XFILLER_50_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__590__B net1971 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_164_ net1869 net171 vssd vssd vccd vccd la_data_in_enable\[1\] sky130_fd_sc_hd__and2_1
XFILLER_10_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_095_ net987 vssd vssd vccd vccd net605 sky130_fd_sc_hd__clkinv_2
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1870 mprj_logic1\[331\] vssd vssd vccd vccd net1870 sky130_fd_sc_hd__buf_6
XANTENNA_output500_A net1126 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1881 net1882 vssd vssd vccd vccd net1881 sky130_fd_sc_hd__buf_6
XFILLER_37_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1892 net1893 vssd vssd vccd vccd net1892 sky130_fd_sc_hd__buf_6
XFILLER_20_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1131_A net495 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1229_A net1230 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__456__A_N net1530 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__484__C net21 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_170 net1585 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_181 net1811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_192 net1820 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] la_data_in_enable\[12\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[12\] sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[25\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_50_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1765_A net1766 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1932_A net1933 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__021__A la_data_in_mprj_bar\[38\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[27\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] net1313 vssd vssd vccd vccd la_data_in_mprj_bar\[123\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_2_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2079_A net2080 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1100 net529 vssd vssd vccd vccd net1100 sky130_fd_sc_hd__buf_6
XANTENNA_user_wb_dat_gates\[18\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1111 net517 vssd vssd vccd vccd net1111 sky130_fd_sc_hd__buf_6
Xwire1122 net505 vssd vssd vccd vccd net1122 sky130_fd_sc_hd__buf_6
XFILLER_43_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input231_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1133 net1134 vssd vssd vccd vccd net1133 sky130_fd_sc_hd__buf_6
XANTENNA_input329_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__479__A_N net272 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1144 net502 vssd vssd vccd vccd net1144 sky130_fd_sc_hd__buf_6
Xwire1155 net1156 vssd vssd vccd vccd net1155 sky130_fd_sc_hd__buf_6
Xwire1166 net1167 vssd vssd vccd vccd net1166 sky130_fd_sc_hd__buf_8
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1177 net929 vssd vssd vccd vccd net1177 sky130_fd_sc_hd__buf_6
Xwire1188 net1189 vssd vssd vccd vccd net1188 sky130_fd_sc_hd__buf_6
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1199 net1200 vssd vssd vccd vccd net1199 sky130_fd_sc_hd__buf_6
XFILLER_38_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__585__B net1977 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_216_ mprj_logic1\[383\] net208 vssd vssd vccd vccd la_data_in_enable\[53\] sky130_fd_sc_hd__and2_2
XFILLER_11_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__106__A net981 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_147_ la_data_in_mprj_bar\[0\] vssd vssd vccd vccd net591 sky130_fd_sc_hd__inv_2
XFILLER_13_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_078_ net962 vssd vssd vccd vccd net713 sky130_fd_sc_hd__clkinv_4
XFILLER_45_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output548_A net1079 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1081_A net545 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1179_A net1180 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__479__C net16 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output715_A net715 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1346_A net1347 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__495__B net2069 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1513_A net1514 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1882_A mprj_logic1\[327\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire966_A la_data_in_mprj_bar\[91\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__016__A la_data_in_mprj_bar\[33\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput108 la_data_out_mprj[79] vssd vssd vccd vccd net108 sky130_fd_sc_hd__buf_6
XANTENNA__389__C net44 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput119 la_data_out_mprj[89] vssd vssd vccd vccd net119 sky130_fd_sc_hd__clkbuf_4
XTAP_4607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_70 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_001_ la_data_in_mprj_bar\[18\] vssd vssd vccd vccd net628 sky130_fd_sc_hd__inv_2
XFILLER_29_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_81 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_92 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input181_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2196_A mprj_logic1\[139\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input446_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input42_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__596__A net1527 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output498_A net1128 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1296_A net1297 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output832_A net832 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1463_A net1464 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1630_A net103 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1728_A mprj_logic1\[460\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput90 la_data_out_mprj[62] vssd vssd vccd vccd net90 sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_550_ net336 mprj_logic1\[255\] vssd vssd vccd vccd net795 sky130_fd_sc_hd__and2_2
XFILLER_17_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_481_ net1594 net2110 net18 vssd vssd vccd vccd net477 sky130_fd_sc_hd__and3b_1
XFILLER_16_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2111_A mprj_logic1\[186\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2209_A net953 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input396_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput450 mprj_dat_o_core[7] vssd vssd vccd vccd net450 sky130_fd_sc_hd__buf_6
XFILLER_23_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput461 user_irq_ena[1] vssd vssd vccd vccd net461 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1044_A net846 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3644 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1211_A net1212 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output782_A net1018 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1309_A net955 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__492__C net30 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3254 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1678_A net1679 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput902 net902 vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_8
XFILLER_29_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput913 net1251 vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput924 net1249 vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_9_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput935 net1246 vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_25_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput946 net1289 vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__buf_8
Xoutput957 net957 vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_8
XFILLER_3_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1845_A mprj_logic1\[347\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_442 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__204__A net1822 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3090 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input144_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2061_A mprj_logic1\[204\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2159_A net2160 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_602_ net1602 net1941 vssd vssd vccd vccd net725 sky130_fd_sc_hd__and2_4
XTAP_4278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input311_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input409_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_533_ net1568 mprj_logic1\[238\] vssd vssd vccd vccd net776 sky130_fd_sc_hd__and2_4
XFILLER_2_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__B net1965 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ net382 net2140 net126 vssd vssd vccd vccd net585 sky130_fd_sc_hd__and3b_4
XTAP_2898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_395_ net306 mprj_logic1\[100\] net50 vssd vssd vccd vccd net509 sky130_fd_sc_hd__and3b_4
XFILLER_35_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output530_A net1099 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1161_A net933 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1259_A net856 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__487__C net24 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput280 la_oenb_mprj[118] vssd vssd vccd vccd net280 sky130_fd_sc_hd__buf_6
Xinput291 la_oenb_mprj[12] vssd vssd vccd vccd net291 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] la_data_in_enable\[42\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[42\] sky130_fd_sc_hd__nand2_2
XFILLER_18_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1795_A net1796 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1962_A mprj_logic1\[2\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput710 net710 vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_8
Xoutput721 net721 vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__buf_8
XANTENNA__024__A la_data_in_mprj_bar\[41\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput732 net732 vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__buf_8
XFILLER_47_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput743 net743 vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__buf_8
Xoutput754 net1036 vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__buf_8
XFILLER_9_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput765 net1026 vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] la_data_in_enable\[4\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[4\] sky130_fd_sc_hd__nand2_1
Xoutput776 net776 vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__buf_8
XFILLER_25_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput787 net787 vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__buf_8
Xwire2208 net2209 vssd vssd vccd vccd net2208 sky130_fd_sc_hd__buf_6
Xoutput798 net1002 vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__buf_8
XFILLER_42_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1507 net1508 vssd vssd vccd vccd net1507 sky130_fd_sc_hd__buf_6
XFILLER_5_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1518 net1519 vssd vssd vccd vccd net1518 sky130_fd_sc_hd__buf_6
XFILLER_21_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1529 net374 vssd vssd vccd vccd net1529 sky130_fd_sc_hd__buf_6
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__397__C net52 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_180_ net1845 net168 vssd vssd vccd vccd la_data_in_enable\[17\] sky130_fd_sc_hd__and2_4
XFILLER_10_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input261_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_622 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input359_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__588__B net1973 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_516_ net298 net2034 vssd vssd vccd vccd net757 sky130_fd_sc_hd__and2_4
XTAP_2673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__109__A net980 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_447_ net1539 net2173 net1626 vssd vssd vccd vccd net566 sky130_fd_sc_hd__and3b_4
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1007_A net1008 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_378_ net387 net1668 net131 vssd vssd vccd vccd net590 sky130_fd_sc_hd__and3b_4
XANTENNA_output480_A net480 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output578_A net1077 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output745_A net745 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__385__A_N net295 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1376_A net430 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output912_A net912 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__498__B net2062 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1543_A net359 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1710_A mprj_logic1\[63\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1808_A mprj_logic1\[411\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire996_A net804 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__019__A la_data_in_mprj_bar\[36\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput540 net1089 vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__buf_8
XFILLER_25_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput551 net551 vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__buf_8
XFILLER_9_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput562 net562 vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__buf_8
Xoutput573 net573 vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__buf_8
XFILLER_43_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput584 net1072 vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__buf_8
Xwire2005 net2006 vssd vssd vccd vccd net2005 sky130_fd_sc_hd__buf_6
Xoutput595 net595 vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_8
XFILLER_21_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2016 mprj_logic1\[270\] vssd vssd vccd vccd net2016 sky130_fd_sc_hd__buf_6
Xwire2027 mprj_logic1\[230\] vssd vssd vccd vccd net2027 sky130_fd_sc_hd__buf_6
Xwire2038 mprj_logic1\[218\] vssd vssd vccd vccd net2038 sky130_fd_sc_hd__buf_6
XFILLER_25_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1304 net1305 vssd vssd vccd vccd net1304 sky130_fd_sc_hd__buf_6
Xwire2049 net2050 vssd vssd vccd vccd net2049 sky130_fd_sc_hd__buf_6
Xwire1315 la_data_in_enable\[107\] vssd vssd vccd vccd net1315 sky130_fd_sc_hd__buf_6
XFILLER_8_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1326 la_data_in_enable\[88\] vssd vssd vccd vccd net1326 sky130_fd_sc_hd__buf_8
Xwire1337 net95 vssd vssd vccd vccd net1337 sky130_fd_sc_hd__buf_6
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1348 net1349 vssd vssd vccd vccd net1348 sky130_fd_sc_hd__buf_6
XFILLER_28_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1359 net444 vssd vssd vccd vccd net1359 sky130_fd_sc_hd__buf_6
XFILLER_3_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_301_ net1698 net454 vssd vssd vccd vccd net945 sky130_fd_sc_hd__and2_4
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_232_ net1813 net225 vssd vssd vccd vccd la_data_in_enable\[69\] sky130_fd_sc_hd__and2_2
XFILLER_24_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_163_ la_data_in_mprj_bar\[16\] vssd vssd vccd vccd net626 sky130_fd_sc_hd__clkinv_2
XFILLER_32_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_094_ net988 vssd vssd vccd vccd net604 sky130_fd_sc_hd__clkinv_2
XANTENNA_input72_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__599__A net1605 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1860 mprj_logic1\[337\] vssd vssd vccd vccd net1860 sky130_fd_sc_hd__buf_6
Xwire1871 mprj_logic1\[330\] vssd vssd vccd vccd net1871 sky130_fd_sc_hd__buf_6
Xwire1882 mprj_logic1\[327\] vssd vssd vccd vccd net1882 sky130_fd_sc_hd__buf_6
XFILLER_24_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1893 net1894 vssd vssd vccd vccd net1893 sky130_fd_sc_hd__buf_6
XFILLER_18_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1124_A net503 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_160 net1370 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_171 net1742 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_182 net1811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 net1820 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output862_A net1254 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[18\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1660_A mprj_logic1\[87\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1758_A mprj_logic1\[447\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__302__A net1676 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1925_A net1926 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] la_data_in_enable\[116\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[116\] sky130_fd_sc_hd__nand2_4
XFILLER_28_128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__400__A_N net312 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__212__A mprj_logic1\[379\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1101 net528 vssd vssd vccd vccd net1101 sky130_fd_sc_hd__buf_6
XFILLER_0_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1112 net516 vssd vssd vccd vccd net1112 sky130_fd_sc_hd__buf_6
Xwire1123 net504 vssd vssd vccd vccd net1123 sky130_fd_sc_hd__buf_6
XFILLER_5_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1134 net485 vssd vssd vccd vccd net1134 sky130_fd_sc_hd__buf_6
XFILLER_43_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1145 net463 vssd vssd vccd vccd net1145 sky130_fd_sc_hd__buf_6
Xwire1156 net1157 vssd vssd vccd vccd net1156 sky130_fd_sc_hd__buf_6
Xwire1167 net1168 vssd vssd vccd vccd net1167 sky130_fd_sc_hd__buf_6
XANTENNA_wire2141_A mprj_logic1\[168\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input224_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1178 net1179 vssd vssd vccd vccd net1178 sky130_fd_sc_hd__buf_8
XFILLER_1_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1189 net926 vssd vssd vccd vccd net1189 sky130_fd_sc_hd__buf_6
XFILLER_28_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_215_ mprj_logic1\[382\] net207 vssd vssd vccd vccd la_data_in_enable\[52\] sky130_fd_sc_hd__and2_2
XFILLER_11_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_146_ mprj_ack_i_core_bar vssd vssd vccd vccd net847 sky130_fd_sc_hd__inv_2
XFILLER_32_1685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_077_ net963 vssd vssd vccd vccd net712 sky130_fd_sc_hd__inv_2
XFILLER_10_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__122__A mprj_dat_i_core_bar\[8\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1074_A net582 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__423__A_N net337 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output610_A net610 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1241_A net1242 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__495__C net1560 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1690 net1691 vssd vssd vccd vccd net1690 sky130_fd_sc_hd__buf_6
XFILLER_4_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1506_A net1507 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput109 la_data_out_mprj[7] vssd vssd vccd vccd net109 sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2206 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__207__A net1819 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_60 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_000_ la_data_in_mprj_bar\[17\] vssd vssd vccd vccd net627 sky130_fd_sc_hd__clkinv_2
XANTENNA_71 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_82 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_93 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2091_A net2092 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input174_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2189_A net2190 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__A_N net1540 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input341_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input439_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input35_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__596__B net1955 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output560_A net560 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output658_A net658 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_129_ mprj_dat_i_core_bar\[15\] vssd vssd vccd vccd net887 sky130_fd_sc_hd__inv_2
XANTENNA_wire1191_A net1192 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1289_A net1290 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output825_A net825 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1456_A net407 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] la_data_in_enable\[72\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[72\] sky130_fd_sc_hd__nand2_4
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1623_A net111 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1992_A net1993 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__A_N net1607 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput80 la_data_out_mprj[53] vssd vssd vccd vccd net80 sky130_fd_sc_hd__clkbuf_4
Xinput91 la_data_out_mprj[63] vssd vssd vccd vccd net91 sky130_fd_sc_hd__buf_4
XFILLER_43_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[33\]_B la_data_in_enable\[33\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_480_ net1595 net2112 net17 vssd vssd vccd vccd net476 sky130_fd_sc_hd__and3b_2
XFILLER_26_952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3756 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input291_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input389_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2506 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput440 mprj_dat_o_core[27] vssd vssd vccd vccd net440 sky130_fd_sc_hd__buf_6
Xinput451 mprj_dat_o_core[8] vssd vssd vccd vccd net451 sky130_fd_sc_hd__buf_6
Xinput462 user_irq_ena[2] vssd vssd vccd vccd net462 sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1037_A net753 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1204_A net921 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output775_A net775 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output942_A net1232 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput903 net903 vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_8
Xoutput914 net1223 vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_B la_data_in_enable\[15\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xoutput925 net1190 vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__buf_8
XFILLER_47_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput936 net1150 vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_9_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput947 net1284 vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__buf_8
Xoutput958 net958 vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_8
XFILLER_42_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1740_A net1741 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1838_A mprj_logic1\[353\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__A net2155 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__204__B net195 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input137_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_601_ net1603 net1943 vssd vssd vccd vccd net724 sky130_fd_sc_hd__and2_4
XTAP_4268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_532_ net1569 mprj_logic1\[237\] vssd vssd vccd vccd net775 sky130_fd_sc_hd__and2_4
XTAP_2822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input304_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_463_ net381 net2141 net125 vssd vssd vccd vccd net584 sky130_fd_sc_hd__and3b_4
XTAP_2877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_394_ net305 net1635 net49 vssd vssd vccd vccd net508 sky130_fd_sc_hd__and3b_4
XFILLER_31_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output523_A net1105 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__130__A mprj_dat_i_core_bar\[16\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1154_A net1155 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput270 la_oenb_mprj[109] vssd vssd vccd vccd net270 sky130_fd_sc_hd__buf_6
XFILLER_20_3579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput281 la_oenb_mprj[119] vssd vssd vccd vccd net281 sky130_fd_sc_hd__buf_6
XFILLER_7_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput292 la_oenb_mprj[13] vssd vssd vccd vccd net292 sky130_fd_sc_hd__buf_4
XFILLER_36_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1321_A la_data_in_enable\[93\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1419_A net1420 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] la_data_in_enable\[35\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[35\] sky130_fd_sc_hd__nand2_1
XFILLER_51_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1690_A net1691 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1788_A mprj_logic1\[431\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__305__A net2201 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1955_A net1956 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput700 net700 vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_8
XFILLER_9_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput711 net711 vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_8
Xoutput722 net722 vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__buf_8
Xoutput733 net733 vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__buf_8
Xoutput744 net744 vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__buf_8
Xoutput755 net1035 vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__buf_8
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput766 net766 vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__buf_8
XFILLER_9_3687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput777 net777 vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__buf_8
XFILLER_5_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput788 net788 vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__buf_8
XFILLER_25_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput799 net799 vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__buf_8
Xwire2209 net953 vssd vssd vccd vccd net2209 sky130_fd_sc_hd__buf_6
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1508 net394 vssd vssd vccd vccd net1508 sky130_fd_sc_hd__buf_6
XFILLER_28_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1519 net390 vssd vssd vccd vccd net1519 sky130_fd_sc_hd__buf_6
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__215__A mprj_logic1\[382\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1750 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2171_A net2172 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input254_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input421_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_515_ net297 net2035 vssd vssd vccd vccd net756 sky130_fd_sc_hd__and2_2
XTAP_2652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_446_ net1540 net2175 net1627 vssd vssd vccd vccd net565 sky130_fd_sc_hd__and3b_4
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_377_ net376 net1670 net120 vssd vssd vccd vccd net579 sky130_fd_sc_hd__and3b_4
XFILLER_48_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output473_A net1057 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output640_A net640 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output738_A net738 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3755 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1271_A net1272 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1369_A net435 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1536_A net367 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__035__A la_data_in_mprj_bar\[52\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput530 net1099 vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__buf_8
Xoutput541 net1087 vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__buf_8
Xoutput552 net552 vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__buf_8
XFILLER_25_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput563 net563 vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__buf_8
XFILLER_47_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput574 net574 vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__buf_8
Xoutput585 net1071 vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__buf_8
Xwire2006 mprj_logic1\[277\] vssd vssd vccd vccd net2006 sky130_fd_sc_hd__buf_6
Xoutput596 net596 vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_8
Xwire2017 mprj_logic1\[269\] vssd vssd vccd vccd net2017 sky130_fd_sc_hd__buf_6
XFILLER_5_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2028 mprj_logic1\[228\] vssd vssd vccd vccd net2028 sky130_fd_sc_hd__buf_6
XFILLER_25_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2039 mprj_logic1\[217\] vssd vssd vccd vccd net2039 sky130_fd_sc_hd__buf_6
Xwire1305 net949 vssd vssd vccd vccd net1305 sky130_fd_sc_hd__buf_6
Xwire1316 la_data_in_enable\[103\] vssd vssd vccd vccd net1316 sky130_fd_sc_hd__buf_6
Xwire1327 la_data_in_enable\[87\] vssd vssd vccd vccd net1327 sky130_fd_sc_hd__buf_8
Xwire1338 net94 vssd vssd vccd vccd net1338 sky130_fd_sc_hd__buf_6
Xwire1349 net450 vssd vssd vccd vccd net1349 sky130_fd_sc_hd__buf_6
XFILLER_41_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3924 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_858 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_300_ net1714 net1341 vssd vssd vccd vccd net950 sky130_fd_sc_hd__and2_4
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2017_A mprj_logic1\[269\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_231_ net1814 net1609 vssd vssd vccd vccd la_data_in_enable\[68\] sky130_fd_sc_hd__and2_2
XFILLER_32_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_162_ la_data_in_mprj_bar\[15\] vssd vssd vccd vccd net625 sky130_fd_sc_hd__clkinv_2
XFILLER_10_3534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_093_ net989 vssd vssd vccd vccd net603 sky130_fd_sc_hd__inv_2
XANTENNA_input371_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_910 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input65_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__599__B net1948 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1850 net1851 vssd vssd vccd vccd net1850 sky130_fd_sc_hd__buf_6
XFILLER_21_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1861 mprj_logic1\[336\] vssd vssd vccd vccd net1861 sky130_fd_sc_hd__buf_6
XFILLER_24_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1872 net1873 vssd vssd vccd vccd net1872 sky130_fd_sc_hd__buf_6
Xwire1883 net1884 vssd vssd vccd vccd net1883 sky130_fd_sc_hd__buf_6
Xwire1894 mprj_logic1\[323\] vssd vssd vccd vccd net1894 sky130_fd_sc_hd__buf_6
XTAP_3150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 net141 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 net1370 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 net1742 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_183 net1813 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output590_A net1136 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 net1820 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1117_A net510 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output688_A net688 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ net344 mprj_logic1\[134\] net88 vssd vssd vccd vccd net547 sky130_fd_sc_hd__and3b_4
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output855_A net1260 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1486_A net1487 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1653_A mprj_logic1\[90\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__302__B net455 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput1 caravel_clk vssd vssd vccd vccd net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] la_data_in_enable\[109\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[109\] sky130_fd_sc_hd__nand2_8
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__212__B net203 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1102 net527 vssd vssd vccd vccd net1102 sky130_fd_sc_hd__buf_6
XFILLER_5_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1113 net515 vssd vssd vccd vccd net1113 sky130_fd_sc_hd__buf_6
XFILLER_22_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1124 net503 vssd vssd vccd vccd net1124 sky130_fd_sc_hd__buf_6
Xwire1135 net474 vssd vssd vccd vccd net1135 sky130_fd_sc_hd__buf_6
XFILLER_19_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1146 net1147 vssd vssd vccd vccd net1146 sky130_fd_sc_hd__buf_8
XFILLER_5_2477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1157 net934 vssd vssd vccd vccd net1157 sky130_fd_sc_hd__buf_6
XFILLER_47_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1168 net1169 vssd vssd vccd vccd net1168 sky130_fd_sc_hd__buf_6
Xwire1179 net1180 vssd vssd vccd vccd net1179 sky130_fd_sc_hd__buf_6
XFILLER_19_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2134_A mprj_logic1\[174\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input217_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3754 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_214_ mprj_logic1\[381\] net206 vssd vssd vccd vccd la_data_in_enable\[51\] sky130_fd_sc_hd__and2_2
XFILLER_7_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_145_ mprj_dat_i_core_bar\[31\] vssd vssd vccd vccd net905 sky130_fd_sc_hd__clkinv_2
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[0\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_076_ net964 vssd vssd vccd vccd net711 sky130_fd_sc_hd__inv_2
XFILLER_23_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1067_A net589 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output603_A net603 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1680 net1681 vssd vssd vccd vccd net1680 sky130_fd_sc_hd__buf_6
XFILLER_39_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1691 mprj_logic1\[73\] vssd vssd vccd vccd net1691 sky130_fd_sc_hd__buf_6
XFILLER_34_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1401_A net1402 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[30\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1770_A mprj_logic1\[441\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1868_A mprj_logic1\[332\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__313__A mprj_logic1\[18\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__398__A_N net1574 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__207__B net198 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_50 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_61 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_72 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_83 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_94 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2084_A mprj_logic1\[196\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input167_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input334_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input28_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_128_ mprj_dat_i_core_bar\[14\] vssd vssd vccd vccd net886 sky130_fd_sc_hd__inv_2
XFILLER_29_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output553_A net553 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__133__A mprj_dat_i_core_bar\[19\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_059_ la_data_in_mprj_bar\[76\] vssd vssd vccd vccd net692 sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1184_A net1185 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output720_A net720 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output818_A net818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1351_A net449 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1449_A net1450 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] la_data_in_enable\[65\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[65\] sky130_fd_sc_hd__nand2_4
XFILLER_40_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1616_A net118 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__308__A net2195 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1985_A mprj_logic1\[287\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire971_A la_data_in_mprj_bar\[86\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput70 la_data_out_mprj[44] vssd vssd vccd vccd net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_4239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput81 la_data_out_mprj[54] vssd vssd vccd vccd net81 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput92 la_data_out_mprj[64] vssd vssd vccd vccd net92 sky130_fd_sc_hd__buf_4
XFILLER_45_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__218__A mprj_logic1\[385\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__413__A_N net326 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input284_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input451_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3936 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vssd vccd vccd net430 sky130_fd_sc_hd__buf_6
XFILLER_23_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput441 mprj_dat_o_core[28] vssd vssd vccd vccd net441 sky130_fd_sc_hd__buf_6
XFILLER_48_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput452 mprj_dat_o_core[9] vssd vssd vccd vccd net452 sky130_fd_sc_hd__buf_6
XFILLER_2_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output768_A net768 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1399_A net1400 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output935_A net1246 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput904 net904 vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_8
Xoutput915 net1220 vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput926 net1186 vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__buf_8
Xoutput937 net1146 vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_47_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput948 net1280 vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__buf_8
XFILLER_25_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput959 net959 vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_8
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1733_A net1734 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__B net1412 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1900_A net1901 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__436__A_N net1550 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__038__A la_data_in_mprj_bar\[55\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__501__A net332 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_600_ net1604 net1945 vssd vssd vccd vccd net723 sky130_fd_sc_hd__and2_4
XTAP_4258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2047_A net2048 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_531_ net315 net2026 vssd vssd vccd vccd net774 sky130_fd_sc_hd__and2_1
XTAP_2812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_462_ net380 mprj_logic1\[167\] net124 vssd vssd vccd vccd net583 sky130_fd_sc_hd__and3b_4
XFILLER_13_4200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_393_ net304 net1637 net48 vssd vssd vccd vccd net507 sky130_fd_sc_hd__and3b_4
XFILLER_25_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input95_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output516_A net1112 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput260 la_oenb_mprj[0] vssd vssd vccd vccd net260 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput271 la_oenb_mprj[10] vssd vssd vccd vccd net271 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput282 la_oenb_mprj[11] vssd vssd vccd vccd net282 sky130_fd_sc_hd__buf_4
Xinput293 la_oenb_mprj[14] vssd vssd vccd vccd net293 sky130_fd_sc_hd__buf_4
XANTENNA_wire1147_A net1148 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__459__A_N net377 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1314_A la_data_in_enable\[114\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] la_data_in_enable\[28\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[28\] sky130_fd_sc_hd__nand2_4
XFILLER_53_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1683_A mprj_logic1\[77\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__305__B net1522 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput701 net701 vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_8
Xoutput712 net712 vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_8
XANTENNA_wire1850_A net1851 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput723 net723 vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__buf_8
XANTENNA_wire1948_A net1949 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput734 net734 vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__buf_8
XFILLER_29_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput745 net745 vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__buf_8
Xoutput756 net1034 vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__buf_8
XFILLER_42_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput767 net1025 vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__buf_8
Xoutput778 net1020 vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__buf_8
Xoutput789 net789 vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__buf_8
XFILLER_42_4484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__321__A mprj_logic1\[26\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_powergood_check_mprj2_vdd_logic1 net954 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1509 net1510 vssd vssd vccd vccd net1509 sky130_fd_sc_hd__buf_6
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__215__B net207 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__231__A net1814 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input247_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3834 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input414_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_514_ net296 net2036 vssd vssd vccd vccd net755 sky130_fd_sc_hd__and2_4
XTAP_2653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_445_ net1541 net2177 net1628 vssd vssd vccd vccd net564 sky130_fd_sc_hd__and3b_4
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ net365 net1672 net109 vssd vssd vccd vccd net568 sky130_fd_sc_hd__and3b_4
XFILLER_31_2216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output466_A net1064 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1097_A net532 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output633_A net633 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__141__A mprj_dat_i_core_bar\[27\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1264_A net1265 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output800_A net1000 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1529_A net374 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1898_A net1899 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__316__A mprj_logic1\[21\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput520 net1108 vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__buf_8
Xoutput531 net1098 vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__buf_8
XFILLER_44_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput542 net1085 vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__buf_8
XFILLER_9_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput553 net553 vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__buf_8
XFILLER_43_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput564 net564 vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__buf_8
Xoutput575 net575 vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__buf_8
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__051__A la_data_in_mprj_bar\[68\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput586 net1070 vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__buf_8
Xwire2007 net2008 vssd vssd vccd vccd net2007 sky130_fd_sc_hd__buf_6
Xoutput597 net597 vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_8
Xwire2018 mprj_logic1\[268\] vssd vssd vccd vccd net2018 sky130_fd_sc_hd__buf_6
Xwire2029 mprj_logic1\[226\] vssd vssd vccd vccd net2029 sky130_fd_sc_hd__buf_6
XFILLER_5_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1306 net880 vssd vssd vccd vccd net1306 sky130_fd_sc_hd__buf_6
XFILLER_5_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1317 la_data_in_enable\[99\] vssd vssd vccd vccd net1317 sky130_fd_sc_hd__buf_6
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1328 la_data_in_enable\[86\] vssd vssd vccd vccd net1328 sky130_fd_sc_hd__buf_8
XFILLER_41_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1339 net93 vssd vssd vccd vccd net1339 sky130_fd_sc_hd__buf_6
XFILLER_38_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_230_ net1815 net1610 vssd vssd vccd vccd la_data_in_enable\[67\] sky130_fd_sc_hd__and2_2
XFILLER_23_583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__226__A mprj_logic1\[393\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_161_ la_data_in_mprj_bar\[14\] vssd vssd vccd vccd net624 sky130_fd_sc_hd__clkinv_2
XFILLER_32_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input197_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_092_ la_data_in_mprj_bar\[109\] vssd vssd vccd vccd net601 sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input364_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input58_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1840 mprj_logic1\[351\] vssd vssd vccd vccd net1840 sky130_fd_sc_hd__buf_6
XFILLER_24_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1851 mprj_logic1\[343\] vssd vssd vccd vccd net1851 sky130_fd_sc_hd__buf_6
XFILLER_20_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1862 mprj_logic1\[335\] vssd vssd vccd vccd net1862 sky130_fd_sc_hd__buf_6
XFILLER_1_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1873 net1874 vssd vssd vccd vccd net1873 sky130_fd_sc_hd__buf_6
Xwire1884 net1885 vssd vssd vccd vccd net1884 sky130_fd_sc_hd__buf_6
XTAP_3140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1895 net1896 vssd vssd vccd vccd net1895 sky130_fd_sc_hd__buf_6
XTAP_3151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_151 net312 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 net1379 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_173 net1742 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 net1813 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 net1829 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ net342 mprj_logic1\[133\] net86 vssd vssd vccd vccd net545 sky130_fd_sc_hd__and3b_4
XFILLER_18_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output583_A net1073 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__136__A mprj_dat_i_core_bar\[22\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_359_ net1709 net1369 vssd vssd vccd vccd net927 sky130_fd_sc_hd__and2_1
XFILLER_35_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output750_A net1040 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1381_A net1382 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1479_A net1480 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] net1319 vssd vssd vccd vccd la_data_in_mprj_bar\[95\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_44_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1646_A net1647 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput2 caravel_clk2 vssd vssd vccd vccd net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__046__A la_data_in_mprj_bar\[63\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1103 net526 vssd vssd vccd vccd net1103 sky130_fd_sc_hd__buf_6
XFILLER_5_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1114 net514 vssd vssd vccd vccd net1114 sky130_fd_sc_hd__buf_6
XFILLER_48_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1125 net501 vssd vssd vccd vccd net1125 sky130_fd_sc_hd__buf_6
XFILLER_9_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1136 net590 vssd vssd vccd vccd net1136 sky130_fd_sc_hd__buf_6
Xwire1147 net1148 vssd vssd vccd vccd net1147 sky130_fd_sc_hd__buf_6
Xwire1158 net1159 vssd vssd vccd vccd net1158 sky130_fd_sc_hd__buf_8
XFILLER_0_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1169 net931 vssd vssd vccd vccd net1169 sky130_fd_sc_hd__buf_6
XFILLER_38_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input112_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_213_ mprj_logic1\[380\] net205 vssd vssd vccd vccd la_data_in_enable\[50\] sky130_fd_sc_hd__and2_2
XFILLER_10_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_144_ mprj_dat_i_core_bar\[30\] vssd vssd vccd vccd net904 sky130_fd_sc_hd__clkinv_2
XFILLER_32_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_075_ net965 vssd vssd vccd vccd net710 sky130_fd_sc_hd__inv_2
XFILLER_27_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__403__B mprj_logic1\[108\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1670 net1671 vssd vssd vccd vccd net1670 sky130_fd_sc_hd__buf_6
XFILLER_20_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1681 mprj_logic1\[78\] vssd vssd vccd vccd net1681 sky130_fd_sc_hd__buf_6
XFILLER_18_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1692 net1693 vssd vssd vccd vccd net1692 sky130_fd_sc_hd__buf_6
XFILLER_0_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1227_A net1228 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output798_A net1002 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] la_data_in_enable\[10\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[10\] sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[23\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_50_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1596_A net272 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1763_A net1764 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__313__B net1401 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1930_A mprj_logic1\[312\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] la_data_in_enable\[121\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[121\] sky130_fd_sc_hd__nand2_4
XFILLER_39_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_40 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_51 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_62 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_73 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_84 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_95 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__504__A net365 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2077_A net2078 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input327_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_954 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__492__A_N net1583 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_49_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_127_ mprj_dat_i_core_bar\[13\] vssd vssd vccd vccd net885 sky130_fd_sc_hd__inv_2
XFILLER_29_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_058_ la_data_in_mprj_bar\[75\] vssd vssd vccd vccd net691 sky130_fd_sc_hd__inv_2
XFILLER_45_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output546_A net1140 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output713_A net713 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1344_A net1345 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2190 mprj_logic1\[144\] vssd vssd vccd vccd net2190 sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] la_data_in_enable\[58\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[58\] sky130_fd_sc_hd__nand2_2
XFILLER_19_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1511_A net393 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__308__B net1422 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1880_A net1881 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1978_A mprj_logic1\[290\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire964_A la_data_in_mprj_bar\[93\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__324__A mprj_logic1\[29\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput60 la_data_out_mprj[35] vssd vssd vccd vccd net60 sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput71 la_data_out_mprj[45] vssd vssd vccd vccd net71 sky130_fd_sc_hd__clkbuf_4
Xinput82 la_data_out_mprj[55] vssd vssd vccd vccd net82 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput93 la_data_out_mprj[65] vssd vssd vccd vccd net93 sky130_fd_sc_hd__buf_6
XFILLER_41_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__234__A mprj_logic1\[401\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2194_A mprj_logic1\[140\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input277_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input444_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input40_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput420 mprj_cyc_o_core vssd vssd vccd vccd net420 sky130_fd_sc_hd__buf_6
Xinput431 mprj_dat_o_core[19] vssd vssd vccd vccd net431 sky130_fd_sc_hd__buf_6
XFILLER_40_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput442 mprj_dat_o_core[29] vssd vssd vccd vccd net442 sky130_fd_sc_hd__buf_6
XANTENNA__400__C net56 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput453 mprj_iena_wb vssd vssd vccd vccd net453 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output496_A net1130 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__144__A mprj_dat_i_core_bar\[30\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A_N net298 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1294_A net1295 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput905 net905 vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_8
XFILLER_49_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput916 net1217 vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output830_A net830 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput927 net1182 vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_28_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput938 net1244 vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__buf_8
XANTENNA_output928_A net1178 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput949 net1303 vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__buf_8
XFILLER_45_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1461_A net406 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1559_A net330 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1726_A net1727 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__054__A la_data_in_mprj_bar\[71\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__501__B net2057 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_530_ net314 mprj_logic1\[235\] vssd vssd vccd vccd net773 sky130_fd_sc_hd__and2_4
XTAP_3558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__229__A mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_461_ net379 net2142 net123 vssd vssd vccd vccd net582 sky130_fd_sc_hd__and3b_4
XFILLER_35_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_392_ net303 net1639 net47 vssd vssd vccd vccd net506 sky130_fd_sc_hd__and3b_4
XFILLER_17_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2207_A net2208 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input394_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input88_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__411__B mprj_logic1\[116\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput250 la_iena_mprj[91] vssd vssd vccd vccd net250 sky130_fd_sc_hd__clkbuf_4
Xinput261 la_oenb_mprj[100] vssd vssd vccd vccd net261 sky130_fd_sc_hd__buf_6
Xinput272 la_oenb_mprj[110] vssd vssd vccd vccd net272 sky130_fd_sc_hd__buf_6
Xinput283 la_oenb_mprj[120] vssd vssd vccd vccd net283 sky130_fd_sc_hd__buf_6
XFILLER_23_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output509_A net1118 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput294 la_oenb_mprj[15] vssd vssd vccd vccd net294 sky130_fd_sc_hd__clkbuf_4
XFILLER_53_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1042_A net1043 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__139__A mprj_dat_i_core_bar\[25\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output780_A net1050 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1307_A net1308 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output878_A net1276 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1676_A net1677 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput702 net702 vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_8
XFILLER_9_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput713 net713 vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_8
Xoutput724 net724 vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__buf_8
XFILLER_9_3645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput735 net735 vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__buf_8
XANTENNA__602__A net1602 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput746 net746 vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__buf_8
XFILLER_29_2861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput757 net1033 vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__buf_8
XFILLER_47_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1843_A mprj_logic1\[349\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput768 net768 vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__buf_8
Xoutput779 net1019 vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__buf_8
XANTENNA__321__B net1501 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__403__A_N net315 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__049__A la_data_in_mprj_bar\[66\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__512__A net294 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__231__B net1609 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input142_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2157_A net2158 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input407_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_513_ net295 net2037 vssd vssd vccd vccd net754 sky130_fd_sc_hd__and2_4
XTAP_2632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_444_ net1542 net2180 net1629 vssd vssd vccd vccd net563 sky130_fd_sc_hd__and3b_4
XTAP_2687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_375_ net354 net1674 net98 vssd vssd vccd vccd net557 sky130_fd_sc_hd__and3b_4
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__406__B mprj_logic1\[111\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__426__A_N net340 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1257_A net858 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1424_A net1425 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] la_data_in_enable\[40\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[40\] sky130_fd_sc_hd__nand2_2
XFILLER_24_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1793_A net1794 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__316__B net1518 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1960_A net1961 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[90\]_B net1324 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput510 net1117 vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__buf_8
XANTENNA__332__A net1817 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput521 net1107 vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__buf_8
XFILLER_9_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput532 net1097 vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__buf_8
XFILLER_44_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput543 net1084 vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__buf_8
Xoutput554 net554 vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] la_data_in_enable\[2\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[2\] sky130_fd_sc_hd__nand2_1
Xoutput565 net565 vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__buf_8
XFILLER_5_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput576 net576 vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__buf_8
Xoutput587 net1069 vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__buf_8
Xwire2008 mprj_logic1\[276\] vssd vssd vccd vccd net2008 sky130_fd_sc_hd__buf_6
Xoutput598 net598 vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_8
Xwire2019 mprj_logic1\[267\] vssd vssd vccd vccd net2019 sky130_fd_sc_hd__buf_6
XFILLER_25_3278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1307 net1308 vssd vssd vccd vccd net1307 sky130_fd_sc_hd__buf_6
XFILLER_3_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1318 la_data_in_enable\[96\] vssd vssd vccd vccd net1318 sky130_fd_sc_hd__buf_8
Xwire1329 la_data_in_enable\[85\] vssd vssd vccd vccd net1329 sky130_fd_sc_hd__buf_8
XFILLER_20_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__507__A net271 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_160_ la_data_in_mprj_bar\[13\] vssd vssd vccd vccd net623 sky130_fd_sc_hd__clkinv_2
XANTENNA__226__B net219 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_091_ net990 vssd vssd vccd vccd net600 sky130_fd_sc_hd__inv_2
XFILLER_32_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_B la_data_in_enable\[81\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__449__A_N net1537 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__242__A mprj_logic1\[409\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input357_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1830 mprj_logic1\[357\] vssd vssd vccd vccd net1830 sky130_fd_sc_hd__buf_6
XFILLER_19_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1841 mprj_logic1\[350\] vssd vssd vccd vccd net1841 sky130_fd_sc_hd__buf_6
XFILLER_24_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1852 net1853 vssd vssd vccd vccd net1852 sky130_fd_sc_hd__buf_6
Xwire1863 net1864 vssd vssd vccd vccd net1863 sky130_fd_sc_hd__buf_6
Xwire1874 net1875 vssd vssd vccd vccd net1874 sky130_fd_sc_hd__buf_6
XFILLER_37_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1885 mprj_logic1\[326\] vssd vssd vccd vccd net1885 sky130_fd_sc_hd__buf_6
XTAP_3141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1896 net1897 vssd vssd vccd vccd net1896 sky130_fd_sc_hd__buf_6
XTAP_3152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 mprj_logic1\[390\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_152 net336 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 net1381 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 net1787 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 net1813 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_196 net1829 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_427_ net1556 mprj_logic1\[132\] net1340 vssd vssd vccd vccd net544 sky130_fd_sc_hd__and3b_4
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_358_ net1710 net1370 vssd vssd vccd vccd net926 sky130_fd_sc_hd__and2_1
XFILLER_50_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1005_A net1006 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output576_A net576 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_289_ net1738 net161 vssd vssd vccd vccd la_data_in_enable\[126\] sky130_fd_sc_hd__and2_4
XFILLER_31_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[72\]_B la_data_in_enable\[72\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_output743_A net743 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1374_A net432 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] net1326 vssd vssd vccd vccd la_data_in_mprj_bar\[88\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1541_A net361 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1639_A net1640 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput3 caravel_rstn vssd vssd vccd vccd net3 sky130_fd_sc_hd__buf_6
XFILLER_4_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire994_A net836 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__327__A mprj_logic1\[32\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__062__A net977 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1104 net525 vssd vssd vccd vccd net1104 sky130_fd_sc_hd__buf_6
XFILLER_44_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1115 net512 vssd vssd vccd vccd net1115 sky130_fd_sc_hd__buf_6
Xwire1126 net500 vssd vssd vccd vccd net1126 sky130_fd_sc_hd__buf_6
XFILLER_5_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1137 net579 vssd vssd vccd vccd net1137 sky130_fd_sc_hd__buf_6
XFILLER_47_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1148 net1149 vssd vssd vccd vccd net1148 sky130_fd_sc_hd__buf_6
XFILLER_21_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1159 net1160 vssd vssd vccd vccd net1159 sky130_fd_sc_hd__buf_6
XFILLER_0_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2022_A mprj_logic1\[264\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__237__A mprj_logic1\[404\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_690 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_212_ mprj_logic1\[379\] net203 vssd vssd vccd vccd la_data_in_enable\[49\] sky130_fd_sc_hd__and2_1
XFILLER_10_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_143_ mprj_dat_i_core_bar\[29\] vssd vssd vccd vccd net902 sky130_fd_sc_hd__clkinv_2
XFILLER_52_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input70_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_074_ net966 vssd vssd vccd vccd net709 sky130_fd_sc_hd__inv_2
XFILLER_45_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__403__C net59 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1660 mprj_logic1\[87\] vssd vssd vccd vccd net1660 sky130_fd_sc_hd__buf_6
Xwire1671 mprj_logic1\[82\] vssd vssd vccd vccd net1671 sky130_fd_sc_hd__buf_6
XFILLER_1_2844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1682 net1683 vssd vssd vccd vccd net1682 sky130_fd_sc_hd__buf_6
Xwire1693 mprj_logic1\[72\] vssd vssd vccd vccd net1693 sky130_fd_sc_hd__buf_6
XFILLER_18_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1122_A net505 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output860_A net1256 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[16\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1491_A net1492 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire990 la_data_in_mprj_bar\[108\] vssd vssd vccd vccd net990 sky130_fd_sc_hd__buf_6
XFILLER_41_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1756_A mprj_logic1\[448\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__610__A net1593 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1923_A net1924 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] net1314 vssd vssd vccd vccd la_data_in_mprj_bar\[114\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_602 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__057__A la_data_in_mprj_bar\[74\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_30 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_41 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_52 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_63 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_74 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[36\]_B la_data_in_enable\[36\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_85 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_96 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__504__B net2052 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_B la_data_in_enable\[120\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_46_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__520__A net303 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input222_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_126_ mprj_dat_i_core_bar\[12\] vssd vssd vccd vccd net884 sky130_fd_sc_hd__inv_2
XANTENNA__414__B mprj_logic1\[119\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B la_data_in_enable\[111\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_057_ la_data_in_mprj_bar\[74\] vssd vssd vccd vccd net690 sky130_fd_sc_hd__inv_2
XFILLER_7_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output539_A net1090 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1072_A net584 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_4190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2180 net2181 vssd vssd vccd vccd net2180 sky130_fd_sc_hd__buf_6
XFILLER_43_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2191 mprj_logic1\[143\] vssd vssd vccd vccd net2191 sky130_fd_sc_hd__buf_6
XANTENNA_wire1337_A net95 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1490 net1491 vssd vssd vccd vccd net1490 sky130_fd_sc_hd__buf_6
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1504_A net395 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[20\]_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__605__A net1599 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1873_A net1874 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__324__B net1490 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[102\]_B la_data_in_enable\[102\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_3402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput50 la_data_out_mprj[26] vssd vssd vccd vccd net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput61 la_data_out_mprj[36] vssd vssd vccd vccd net61 sky130_fd_sc_hd__clkbuf_4
Xinput72 la_data_out_mprj[46] vssd vssd vccd vccd net72 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput83 la_data_out_mprj[56] vssd vssd vccd vccd net83 sky130_fd_sc_hd__buf_4
XFILLER_28_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput94 la_data_out_mprj[66] vssd vssd vccd vccd net94 sky130_fd_sc_hd__buf_6
XFILLER_28_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[11\]_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__515__A net297 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__234__B net228 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input172_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__250__A net1805 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input437_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput410 mprj_adr_o_core[2] vssd vssd vccd vccd net410 sky130_fd_sc_hd__buf_6
Xinput421 mprj_dat_o_core[0] vssd vssd vccd vccd net421 sky130_fd_sc_hd__buf_6
XFILLER_24_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input33_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput432 mprj_dat_o_core[1] vssd vssd vccd vccd net432 sky130_fd_sc_hd__buf_6
XFILLER_0_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput443 mprj_dat_o_core[2] vssd vssd vccd vccd net443 sky130_fd_sc_hd__buf_6
XFILLER_40_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput454 mprj_sel_o_core[0] vssd vssd vccd vccd net454 sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__409__B mprj_logic1\[114\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output489_A net489 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output656_A net656 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_109_ net980 vssd vssd vccd vccd net620 sky130_fd_sc_hd__clkinv_2
Xoutput906 net906 vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_8
Xoutput917 net1214 vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_45_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput928 net1178 vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__buf_8
XFILLER_7_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1287_A net1288 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput939 net1241 vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_45_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output823_A net823 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1454_A net1455 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] la_data_in_enable\[70\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[70\] sky130_fd_sc_hd__nand2_4
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1621_A net113 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__319__B net1509 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1990_A net1991 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__335__A net1809 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__A_N net1593 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__070__A net970 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ net378 net2143 net122 vssd vssd vccd vccd net581 sky130_fd_sc_hd__and3b_4
XTAP_2847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__229__B net222 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_391_ net302 net1641 net46 vssd vssd vccd vccd net505 sky130_fd_sc_hd__and3b_4
XFILLER_53_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2102_A net2103 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__245__A net1807 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input387_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput240 la_iena_mprj[82] vssd vssd vccd vccd net240 sky130_fd_sc_hd__buf_4
XFILLER_20_3549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput251 la_iena_mprj[92] vssd vssd vccd vccd net251 sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput262 la_oenb_mprj[101] vssd vssd vccd vccd net262 sky130_fd_sc_hd__buf_6
Xinput273 la_oenb_mprj[111] vssd vssd vccd vccd net273 sky130_fd_sc_hd__buf_6
XFILLER_48_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput284 la_oenb_mprj[121] vssd vssd vccd vccd net284 sky130_fd_sc_hd__buf_6
Xinput295 la_oenb_mprj[16] vssd vssd vccd vccd net295 sky130_fd_sc_hd__buf_4
XFILLER_18_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1035_A net755 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_589_ net379 net1972 vssd vssd vccd vccd net838 sky130_fd_sc_hd__and2_4
XFILLER_18_3489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1202_A net1203 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output773_A net1024 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__155__A la_data_in_mprj_bar\[8\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output940_A net1238 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput703 net703 vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_8
XANTENNA_wire1571_A net312 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput714 net714 vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_8
XANTENNA_wire1669_A mprj_logic1\[83\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput725 net725 vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__buf_8
XFILLER_47_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput736 net736 vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__buf_8
XANTENNA__602__B net1941 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput747 net747 vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__buf_8
Xoutput758 net1052 vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__buf_8
XFILLER_42_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput769 net1051 vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__buf_8
XFILLER_47_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1836_A mprj_logic1\[354\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__065__A la_data_in_mprj_bar\[82\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__512__B net2039 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2052_A mprj_logic1\[209\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__378__A_N net387 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ net294 net2039 vssd vssd vccd vccd net753 sky130_fd_sc_hd__and2_4
XFILLER_19_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input302_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ net1543 net2182 net1630 vssd vssd vccd vccd net562 sky130_fd_sc_hd__and3b_4
XTAP_2677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ net343 net1678 net87 vssd vssd vccd vccd net546 sky130_fd_sc_hd__and3b_4
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output521_A net1107 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1152_A net1153 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1417_A net1418 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] la_data_in_enable\[33\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[33\] sky130_fd_sc_hd__nand2_4
XFILLER_51_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__613__A net1590 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1953_A net1954 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput500 net1126 vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__buf_8
Xoutput511 net1116 vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__buf_8
Xoutput522 net1106 vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__buf_8
XANTENNA__332__B net1452 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput533 net1096 vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__buf_8
XFILLER_47_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput544 net1082 vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__buf_8
Xoutput555 net555 vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__buf_8
XFILLER_47_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput566 net566 vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput577 net577 vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__buf_8
XFILLER_5_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput588 net1068 vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__buf_8
Xwire2009 mprj_logic1\[275\] vssd vssd vccd vccd net2009 sky130_fd_sc_hd__buf_6
Xoutput599 net599 vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_8
XFILLER_42_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1308 net1309 vssd vssd vccd vccd net1308 sky130_fd_sc_hd__buf_6
XFILLER_25_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1319 la_data_in_enable\[95\] vssd vssd vccd vccd net1319 sky130_fd_sc_hd__buf_6
XFILLER_25_2589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__507__B net2047 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_090_ net991 vssd vssd vccd vccd net599 sky130_fd_sc_hd__clkinv_2
XFILLER_13_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__523__A net306 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input252_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1820 mprj_logic1\[373\] vssd vssd vccd vccd net1820 sky130_fd_sc_hd__buf_6
Xwire1831 net1832 vssd vssd vccd vccd net1831 sky130_fd_sc_hd__buf_6
XFILLER_24_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1842 mprj_logic1\[34\] vssd vssd vccd vccd net1842 sky130_fd_sc_hd__buf_6
XFILLER_21_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1853 mprj_logic1\[342\] vssd vssd vccd vccd net1853 sky130_fd_sc_hd__buf_6
Xwire1864 mprj_logic1\[334\] vssd vssd vccd vccd net1864 sky130_fd_sc_hd__buf_6
XFILLER_19_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1875 mprj_logic1\[329\] vssd vssd vccd vccd net1875 sky130_fd_sc_hd__buf_6
XFILLER_18_324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1886 net1887 vssd vssd vccd vccd net1886 sky130_fd_sc_hd__buf_6
XFILLER_37_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1897 mprj_logic1\[322\] vssd vssd vccd vccd net1897 sky130_fd_sc_hd__buf_6
XTAP_3153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 mprj_logic1\[390\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_153 net1352 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_164 net1401 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 net1787 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 net1818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_426_ net340 mprj_logic1\[131\] net84 vssd vssd vccd vccd net543 sky130_fd_sc_hd__and3b_4
XANTENNA_197 net1829 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__417__B mprj_logic1\[122\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ net1711 net1371 vssd vssd vccd vccd net925 sky130_fd_sc_hd__and2_1
XFILLER_32_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_288_ net1740 net160 vssd vssd vccd vccd la_data_in_enable\[125\] sky130_fd_sc_hd__and2_4
XANTENNA_output471_A net1059 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output569_A net569 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_740 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output736_A net736 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1367_A net437 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1534_A net369 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput4 la_data_out_mprj[0] vssd vssd vccd vccd net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1701_A mprj_logic1\[69\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__608__A net1595 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__327__B net1475 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire987_A la_data_in_mprj_bar\[112\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__343__A mprj_logic1\[48\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1105 net523 vssd vssd vccd vccd net1105 sky130_fd_sc_hd__buf_6
XFILLER_40_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1116 net511 vssd vssd vccd vccd net1116 sky130_fd_sc_hd__buf_6
Xwire1127 net499 vssd vssd vccd vccd net1127 sky130_fd_sc_hd__buf_6
XFILLER_9_1893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1138 net568 vssd vssd vccd vccd net1138 sky130_fd_sc_hd__buf_6
Xwire1149 net937 vssd vssd vccd vccd net1149 sky130_fd_sc_hd__buf_6
XFILLER_27_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__A net301 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__237__B net231 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2015_A mprj_logic1\[271\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__416__A_N net329 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_211_ mprj_logic1\[378\] net202 vssd vssd vccd vccd la_data_in_enable\[48\] sky130_fd_sc_hd__and2_1
XFILLER_49_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_142_ mprj_dat_i_core_bar\[28\] vssd vssd vccd vccd net901 sky130_fd_sc_hd__clkinv_2
XFILLER_32_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__253__A mprj_logic1\[420\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_073_ net967 vssd vssd vccd vccd net708 sky130_fd_sc_hd__clkinv_2
XFILLER_10_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input63_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1650 net1651 vssd vssd vccd vccd net1650 sky130_fd_sc_hd__buf_6
XFILLER_21_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1661 net1662 vssd vssd vccd vccd net1661 sky130_fd_sc_hd__buf_6
XFILLER_47_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1672 net1673 vssd vssd vccd vccd net1672 sky130_fd_sc_hd__buf_6
Xwire1683 mprj_logic1\[77\] vssd vssd vccd vccd net1683 sky130_fd_sc_hd__buf_6
XFILLER_19_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1694 net1695 vssd vssd vccd vccd net1694 sky130_fd_sc_hd__buf_6
XFILLER_19_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1115_A net512 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output686_A net686 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_409_ net322 mprj_logic1\[114\] net66 vssd vssd vccd vccd net525 sky130_fd_sc_hd__and3b_4
XFILLER_50_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output853_A net1262 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__163__A la_data_in_mprj_bar\[16\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1484_A net400 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire980 la_data_in_mprj_bar\[126\] vssd vssd vccd vccd net980 sky130_fd_sc_hd__buf_6
XFILLER_31_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire991 la_data_in_mprj_bar\[107\] vssd vssd vccd vccd net991 sky130_fd_sc_hd__buf_6
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1749_A net1750 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__610__B net1919 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1916_A net1917 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] net1315 vssd vssd vccd vccd la_data_in_mprj_bar\[107\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__439__A_N net1547 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__338__A mprj_logic1\[43\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_20 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_31 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_42 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_53 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_64 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_75 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__073__A net967 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_86 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_97 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__520__B net2030 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3750 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input215_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2132_A mprj_logic1\[175\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__248__A mprj_logic1\[415\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_125_ mprj_dat_i_core_bar\[11\] vssd vssd vccd vccd net883 sky130_fd_sc_hd__inv_2
XFILLER_32_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__C net71 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_056_ la_data_in_mprj_bar\[73\] vssd vssd vccd vccd net689 sky130_fd_sc_hd__inv_2
XFILLER_10_2485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__430__B mprj_logic1\[135\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1065_A net465 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2170 mprj_logic1\[154\] vssd vssd vccd vccd net2170 sky130_fd_sc_hd__buf_6
XFILLER_21_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2181 mprj_logic1\[149\] vssd vssd vccd vccd net2181 sky130_fd_sc_hd__buf_6
Xwire2192 mprj_logic1\[142\] vssd vssd vccd vccd net2192 sky130_fd_sc_hd__buf_6
XFILLER_43_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1480 net1481 vssd vssd vccd vccd net1480 sky130_fd_sc_hd__buf_6
Xwire1491 net1492 vssd vssd vccd vccd net1491 sky130_fd_sc_hd__buf_6
XANTENNA_wire1232_A net1233 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1699_A mprj_logic1\[6\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__605__B net1934 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput40 la_data_out_mprj[17] vssd vssd vccd vccd net40 sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1866_A mprj_logic1\[333\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput51 la_data_out_mprj[27] vssd vssd vccd vccd net51 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput62 la_data_out_mprj[37] vssd vssd vccd vccd net62 sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput73 la_data_out_mprj[47] vssd vssd vccd vccd net73 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput84 la_data_out_mprj[57] vssd vssd vccd vccd net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput95 la_data_out_mprj[67] vssd vssd vccd vccd net95 sky130_fd_sc_hd__buf_6
XFILLER_45_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__621__A net1582 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__340__B net1356 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__068__A net972 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[11\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__515__B net2035 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__531__A net315 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input165_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2082_A net2083 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2278 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput400 mprj_adr_o_core[20] vssd vssd vccd vccd net400 sky130_fd_sc_hd__buf_6
XFILLER_2_4353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput411 mprj_adr_o_core[30] vssd vssd vccd vccd net411 sky130_fd_sc_hd__buf_6
XFILLER_40_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput422 mprj_dat_o_core[10] vssd vssd vccd vccd net422 sky130_fd_sc_hd__buf_6
XFILLER_7_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input332_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput433 mprj_dat_o_core[20] vssd vssd vccd vccd net433 sky130_fd_sc_hd__buf_6
XFILLER_48_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput444 mprj_dat_o_core[30] vssd vssd vccd vccd net444 sky130_fd_sc_hd__buf_6
XFILLER_0_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput455 mprj_sel_o_core[1] vssd vssd vccd vccd net455 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input26_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__409__C net66 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__425__B mprj_logic1\[130\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_108_ la_data_in_mprj_bar\[125\] vssd vssd vccd vccd net619 sky130_fd_sc_hd__inv_2
XFILLER_9_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput907 net907 vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_8
XFILLER_49_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output551_A net551 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput918 net1211 vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__buf_8
Xoutput929 net1174 vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__buf_8
XANTENNA_output649_A net649 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_039_ la_data_in_mprj_bar\[56\] vssd vssd vccd vccd net670 sky130_fd_sc_hd__inv_2
XANTENNA_wire1182_A net1183 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output816_A net816 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1447_A net1448 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] la_data_in_enable\[63\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[63\] sky130_fd_sc_hd__nand2_4
XFILLER_36_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__616__A net1587 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1983_A mprj_logic1\[288\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__335__B net1432 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__351__A net1718 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_390_ net301 net1643 net45 vssd vssd vccd vccd net504 sky130_fd_sc_hd__and3b_4
XFILLER_52_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__526__A net1574 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__245__B net240 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input282_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__A net1793 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput230 la_iena_mprj[73] vssd vssd vccd vccd net230 sky130_fd_sc_hd__clkbuf_4
Xinput241 la_iena_mprj[83] vssd vssd vccd vccd net241 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput252 la_iena_mprj[93] vssd vssd vccd vccd net252 sky130_fd_sc_hd__clkbuf_4
Xinput263 la_oenb_mprj[102] vssd vssd vccd vccd net263 sky130_fd_sc_hd__buf_6
Xinput274 la_oenb_mprj[112] vssd vssd vccd vccd net274 sky130_fd_sc_hd__buf_6
XFILLER_49_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput285 la_oenb_mprj[122] vssd vssd vccd vccd net285 sky130_fd_sc_hd__buf_6
XFILLER_18_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput296 la_oenb_mprj[17] vssd vssd vccd vccd net296 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_588_ net378 net1973 vssd vssd vccd vccd net837 sky130_fd_sc_hd__and2_4
XFILLER_34_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_970 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output766_A net766 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1397_A net420 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1080 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output933_A net1158 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput704 net704 vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_8
XFILLER_29_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput715 net715 vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_8
XANTENNA__171__A net1858 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput726 net726 vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__buf_8
XFILLER_42_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput737 net737 vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__buf_8
XFILLER_47_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1564_A net325 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput748 net748 vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__buf_8
XFILLER_7_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput759 net1032 vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__buf_8
XFILLER_42_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1731_A mprj_logic1\[459\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1829_A mprj_logic1\[358\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__346__A mprj_logic1\[51\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__081__A la_data_in_mprj_bar\[98\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input128_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2045_A net2046 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ net293 net2040 vssd vssd vccd vccd net752 sky130_fd_sc_hd__and2_4
XTAP_3368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ net1544 net2184 net1631 vssd vssd vccd vccd net561 sky130_fd_sc_hd__and3b_4
XFILLER_19_3788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__256__A net1800 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_373_ net332 net1680 net76 vssd vssd vccd vccd net535 sky130_fd_sc_hd__and3b_4
XFILLER_39_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input93_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[9\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_29_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__422__C net80 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output514_A net1114 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1145_A net463 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1312_A la_data_in_enable\[124\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__A_N net264 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__166__A net1865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] la_data_in_enable\[26\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[26\] sky130_fd_sc_hd__nand2_4
XFILLER_14_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1681_A mprj_logic1\[78\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1779_A mprj_logic1\[436\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__613__B net1908 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput501 net1125 vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__buf_8
Xoutput512 net1115 vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__buf_8
XFILLER_5_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput523 net1105 vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__buf_8
XFILLER_25_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput534 net1095 vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__buf_8
XFILLER_44_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1946_A net1947 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput545 net1081 vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__buf_8
XFILLER_25_3236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput556 net556 vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput567 net567 vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__buf_8
XFILLER_5_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput578 net1077 vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__buf_8
Xoutput589 net1067 vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__buf_8
XFILLER_47_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1309 net955 vssd vssd vccd vccd net1309 sky130_fd_sc_hd__buf_6
XFILLER_38_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_358 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__076__A net964 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__523__B net2028 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2162_A net2163 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input245_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1810 mprj_logic1\[400\] vssd vssd vccd vccd net1810 sky130_fd_sc_hd__buf_6
XFILLER_41_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1821 mprj_logic1\[372\] vssd vssd vccd vccd net1821 sky130_fd_sc_hd__buf_6
Xwire1832 mprj_logic1\[356\] vssd vssd vccd vccd net1832 sky130_fd_sc_hd__buf_6
XFILLER_46_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1843 mprj_logic1\[349\] vssd vssd vccd vccd net1843 sky130_fd_sc_hd__buf_6
XFILLER_21_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1854 net1855 vssd vssd vccd vccd net1854 sky130_fd_sc_hd__buf_6
XTAP_3110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1865 net1866 vssd vssd vccd vccd net1865 sky130_fd_sc_hd__buf_6
XTAP_3121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input412_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1876 net1877 vssd vssd vccd vccd net1876 sky130_fd_sc_hd__buf_6
XFILLER_46_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1887 net1888 vssd vssd vccd vccd net1887 sky130_fd_sc_hd__buf_6
XANTENNA__495__A_N net1580 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1898 net1899 vssd vssd vccd vccd net1898 sky130_fd_sc_hd__buf_6
XFILLER_19_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 mprj_logic1\[252\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_121 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 mprj_logic1\[395\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 net1352 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 net1401 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 net1787 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_425_ net339 mprj_logic1\[130\] net83 vssd vssd vccd vccd net542 sky130_fd_sc_hd__and3b_2
XANTENNA_187 net1818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_198 net1837 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__417__C net74 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_356_ net1712 net1375 vssd vssd vccd vccd net923 sky130_fd_sc_hd__and2_1
XFILLER_31_2027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_287_ net1742 net159 vssd vssd vccd vccd la_data_in_enable\[124\] sky130_fd_sc_hd__and2_2
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__B net2197 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output464_A net1066 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1095_A net534 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output729_A net729 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1262_A net1263 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput5 la_data_out_mprj[100] vssd vssd vccd vccd net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__608__B net1925 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1896_A net1897 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__624__A net1579 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__343__B net1350 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1106 net522 vssd vssd vccd vccd net1106 sky130_fd_sc_hd__buf_6
XFILLER_9_1872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1117 net510 vssd vssd vccd vccd net1117 sky130_fd_sc_hd__buf_6
Xwire1128 net498 vssd vssd vccd vccd net1128 sky130_fd_sc_hd__buf_6
XFILLER_38_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1139 net557 vssd vssd vccd vccd net1139 sky130_fd_sc_hd__buf_6
XFILLER_19_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4426 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__B net2032 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_210_ mprj_logic1\[377\] net201 vssd vssd vccd vccd la_data_in_enable\[47\] sky130_fd_sc_hd__and2_1
XFILLER_51_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__534__A net1567 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_141_ mprj_dat_i_core_bar\[27\] vssd vssd vccd vccd net900 sky130_fd_sc_hd__clkinv_2
XFILLER_49_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input195_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__253__B net249 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_072_ net968 vssd vssd vccd vccd net706 sky130_fd_sc_hd__clkinv_2
XFILLER_10_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input362_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input56_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1640 mprj_logic1\[97\] vssd vssd vccd vccd net1640 sky130_fd_sc_hd__buf_6
XFILLER_1_2824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1651 mprj_logic1\[91\] vssd vssd vccd vccd net1651 sky130_fd_sc_hd__buf_6
XFILLER_5_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1662 mprj_logic1\[86\] vssd vssd vccd vccd net1662 sky130_fd_sc_hd__buf_6
XFILLER_19_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1673 mprj_logic1\[81\] vssd vssd vccd vccd net1673 sky130_fd_sc_hd__buf_6
XFILLER_47_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1684 net1685 vssd vssd vccd vccd net1684 sky130_fd_sc_hd__buf_6
XFILLER_24_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1695 mprj_logic1\[71\] vssd vssd vccd vccd net1695 sky130_fd_sc_hd__buf_6
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__428__B mprj_logic1\[133\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ net320 mprj_logic1\[113\] net64 vssd vssd vccd vccd net523 sky130_fd_sc_hd__and3b_4
XFILLER_32_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output581_A net1075 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1108_A net520 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_339_ mprj_logic1\[44\] net1360 vssd vssd vccd vccd net935 sky130_fd_sc_hd__and2_1
XFILLER_35_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire970 la_data_in_mprj_bar\[87\] vssd vssd vccd vccd net970 sky130_fd_sc_hd__buf_6
XANTENNA_output846_A net1044 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire981 la_data_in_mprj_bar\[123\] vssd vssd vccd vccd net981 sky130_fd_sc_hd__buf_6
Xwire992 la_data_in_mprj_bar\[103\] vssd vssd vccd vccd net992 sky130_fd_sc_hd__buf_6
XFILLER_45_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1477_A net1478 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] net1321 vssd vssd vccd vccd la_data_in_mprj_bar\[93\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_41_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1644_A mprj_logic1\[95\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1811_A mprj_logic1\[3\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1909_A net1910 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__619__A net1584 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__338__B net1372 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_10 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_21 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_32 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__354__A net1715 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_43 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_54 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_65 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_76 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_87 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_98 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__529__A net1570 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__248__B net243 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2125_A mprj_logic1\[179\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input208_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__264__A net1787 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_124_ mprj_dat_i_core_bar\[10\] vssd vssd vccd vccd net882 sky130_fd_sc_hd__inv_2
XFILLER_32_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_055_ la_data_in_mprj_bar\[72\] vssd vssd vccd vccd net688 sky130_fd_sc_hd__inv_2
XFILLER_49_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__430__C net89 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2160 net2161 vssd vssd vccd vccd net2160 sky130_fd_sc_hd__buf_6
Xwire2171 net2172 vssd vssd vccd vccd net2171 sky130_fd_sc_hd__buf_6
XFILLER_1_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2182 net2183 vssd vssd vccd vccd net2182 sky130_fd_sc_hd__buf_6
Xwire2193 mprj_logic1\[141\] vssd vssd vccd vccd net2193 sky130_fd_sc_hd__buf_6
XANTENNA_wire1058_A net472 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1470 net1471 vssd vssd vccd vccd net1470 sky130_fd_sc_hd__buf_6
XFILLER_53_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1481 net401 vssd vssd vccd vccd net1481 sky130_fd_sc_hd__buf_6
Xwire1492 net1493 vssd vssd vccd vccd net1492 sky130_fd_sc_hd__buf_6
XFILLER_34_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1225_A net914 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output796_A net796 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__174__A net1854 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[21\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_30_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput30 la_data_out_mprj[123] vssd vssd vccd vccd net30 sky130_fd_sc_hd__buf_4
XFILLER_50_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput41 la_data_out_mprj[18] vssd vssd vccd vccd net41 sky130_fd_sc_hd__clkbuf_4
Xinput52 la_data_out_mprj[28] vssd vssd vccd vccd net52 sky130_fd_sc_hd__clkbuf_4
Xinput63 la_data_out_mprj[38] vssd vssd vccd vccd net63 sky130_fd_sc_hd__clkbuf_4
Xinput74 la_data_out_mprj[48] vssd vssd vccd vccd net74 sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1761_A net1762 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput85 la_data_out_mprj[58] vssd vssd vccd vccd net85 sky130_fd_sc_hd__buf_6
XFILLER_41_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput96 la_data_out_mprj[68] vssd vssd vccd vccd net96 sky130_fd_sc_hd__buf_6
XANTENNA_wire1859_A net1860 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__621__B net1883 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__406__A_N net318 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__349__A mprj_logic1\[54\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__531__B net2026 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2075_A mprj_logic1\[199\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input158_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput401 mprj_adr_o_core[21] vssd vssd vccd vccd net401 sky130_fd_sc_hd__buf_6
Xinput412 mprj_adr_o_core[31] vssd vssd vccd vccd net412 sky130_fd_sc_hd__buf_6
XFILLER_22_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput423 mprj_dat_o_core[11] vssd vssd vccd vccd net423 sky130_fd_sc_hd__buf_6
XFILLER_40_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput434 mprj_dat_o_core[21] vssd vssd vccd vccd net434 sky130_fd_sc_hd__buf_6
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput445 mprj_dat_o_core[31] vssd vssd vccd vccd net445 sky130_fd_sc_hd__buf_6
XFILLER_2_4387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput456 mprj_sel_o_core[2] vssd vssd vccd vccd net456 sky130_fd_sc_hd__buf_4
XANTENNA_input325_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__259__A net1797 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input19_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__425__C net83 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_107_ la_data_in_mprj_bar\[124\] vssd vssd vccd vccd net618 sky130_fd_sc_hd__clkinv_2
XFILLER_32_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput908 net908 vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_8
Xoutput919 net1208 vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__buf_8
XFILLER_45_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__429__A_N net344 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_038_ la_data_in_mprj_bar\[55\] vssd vssd vccd vccd net669 sky130_fd_sc_hd__inv_2
XANTENNA__441__B net2186 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output544_A net1082 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1175_A net1176 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output809_A net809 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1342_A net1343 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__169__A net1861 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] la_data_in_enable\[56\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[56\] sky130_fd_sc_hd__nand2_2
XFILLER_19_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__616__B net1898 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1976_A mprj_logic1\[291\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__351__B net1381 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__079__A la_data_in_mprj_bar\[96\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__526__B mprj_logic1\[231\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__542__A net327 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2192_A mprj_logic1\[142\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__B net257 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input442_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_iena_mprj[64] vssd vssd vccd vccd net220 sky130_fd_sc_hd__buf_4
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput231 la_iena_mprj[74] vssd vssd vccd vccd net231 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput242 la_iena_mprj[84] vssd vssd vccd vccd net242 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput253 la_iena_mprj[94] vssd vssd vccd vccd net253 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput264 la_oenb_mprj[103] vssd vssd vccd vccd net264 sky130_fd_sc_hd__buf_6
Xinput275 la_oenb_mprj[113] vssd vssd vccd vccd net275 sky130_fd_sc_hd__buf_6
XFILLER_2_3483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput286 la_oenb_mprj[123] vssd vssd vccd vccd net286 sky130_fd_sc_hd__buf_6
Xinput297 la_oenb_mprj[18] vssd vssd vccd vccd net297 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_587_ net377 net1975 vssd vssd vccd vccd net836 sky130_fd_sc_hd__and2_2
XFILLER_32_724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__436__B net2193 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output494_A net1132 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_982 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output661_A net661 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output759_A net1032 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1292_A net1293 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput705 net705 vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_8
Xoutput716 net716 vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_8
XFILLER_29_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput727 net727 vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__buf_8
Xoutput738 net738 vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__buf_8
XFILLER_42_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput749 net749 vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__buf_8
XANTENNA_output926_A net1186 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_2897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1724_A net1725 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_890 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__346__B net1344 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[93\]_B net1321 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__362__A net1704 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_510_ net292 net2042 vssd vssd vccd vccd net751 sky130_fd_sc_hd__and2_4
XFILLER_22_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__537__A net1565 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ net1545 net2186 net1632 vssd vssd vccd vccd net560 sky130_fd_sc_hd__and3b_4
XTAP_2657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__256__B net252 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_372_ net321 net1682 net65 vssd vssd vccd vccd net524 sky130_fd_sc_hd__and3b_4
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2205_A net2206 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input392_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B net1330 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input86_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__272__A net1773 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output507_A net1120 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1040_A net750 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1138_A net568 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1305_A net949 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output876_A net1278 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] la_data_in_enable\[19\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[19\] sky130_fd_sc_hd__nand2_2
XFILLER_32_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[75\]_B la_data_in_enable\[75\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__182__A net1843 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1674_A net1675 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput502 net1144 vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__buf_8
XFILLER_44_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput513 net1143 vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__buf_8
XFILLER_48_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput524 net1142 vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__buf_8
Xoutput535 net1141 vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__buf_8
Xoutput546 net1140 vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__buf_8
XFILLER_44_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput557 net1139 vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__buf_8
XANTENNA_wire1841_A mprj_logic1\[350\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput568 net1138 vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__buf_8
XFILLER_25_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1939_A net1940 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput579 net1137 vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__buf_8
XFILLER_5_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__A net1711 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1964 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__092__A la_data_in_mprj_bar\[109\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3990 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1800 mprj_logic1\[423\] vssd vssd vccd vccd net1800 sky130_fd_sc_hd__buf_6
XANTENNA_input140_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1811 mprj_logic1\[3\] vssd vssd vccd vccd net1811 sky130_fd_sc_hd__buf_6
XANTENNA_wire2155_A mprj_logic1\[15\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1822 mprj_logic1\[371\] vssd vssd vccd vccd net1822 sky130_fd_sc_hd__buf_6
XANTENNA_input238_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1833 net1834 vssd vssd vccd vccd net1833 sky130_fd_sc_hd__buf_6
XFILLER_24_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1844 mprj_logic1\[348\] vssd vssd vccd vccd net1844 sky130_fd_sc_hd__buf_6
XFILLER_46_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1855 mprj_logic1\[341\] vssd vssd vccd vccd net1855 sky130_fd_sc_hd__buf_6
XFILLER_18_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1866 mprj_logic1\[333\] vssd vssd vccd vccd net1866 sky130_fd_sc_hd__buf_6
XTAP_3122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1877 net1878 vssd vssd vccd vccd net1877 sky130_fd_sc_hd__buf_6
XTAP_3133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1888 mprj_logic1\[325\] vssd vssd vccd vccd net1888 sky130_fd_sc_hd__buf_6
XFILLER_41_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1899 net1900 vssd vssd vccd vccd net1899 sky130_fd_sc_hd__buf_6
XTAP_3155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input405_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 mprj_logic1\[252\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__267__A net1782 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 mprj_logic1\[395\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1706 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 net1352 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_166 net1401 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_424_ net338 mprj_logic1\[129\] net82 vssd vssd vccd vccd net541 sky130_fd_sc_hd__and3b_1
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 net1811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_188 net1818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_199 net1837 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ net1713 net1376 vssd vssd vccd vccd net922 sky130_fd_sc_hd__and2_1
XFILLER_50_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_286_ net1744 net158 vssd vssd vccd vccd la_data_in_enable\[123\] sky130_fd_sc_hd__and2_4
XFILLER_13_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__433__C net92 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1255_A net862 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput6 la_data_out_mprj[101] vssd vssd vccd vccd net6 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1422_A net1423 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__177__A net1849 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1791_A net1792 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1889_A net1890 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__624__B net1872 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] la_data_in_enable\[0\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[0\] sky130_fd_sc_hd__nand2_2
XFILLER_40_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1107 net521 vssd vssd vccd vccd net1107 sky130_fd_sc_hd__buf_6
XFILLER_29_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1118 net509 vssd vssd vccd vccd net1118 sky130_fd_sc_hd__buf_6
Xwire1129 net497 vssd vssd vccd vccd net1129 sky130_fd_sc_hd__buf_6
XFILLER_25_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__087__A la_data_in_mprj_bar\[104\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_B la_data_in_enable\[39\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_140_ mprj_dat_i_core_bar\[26\] vssd vssd vccd vccd net899 sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[123\]_B net1313 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_071_ net969 vssd vssd vccd vccd net705 sky130_fd_sc_hd__clkinv_2
XFILLER_32_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input188_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__550__A net336 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input355_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__A_N net380 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input49_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1630 net103 vssd vssd vccd vccd net1630 sky130_fd_sc_hd__buf_6
Xwire1641 net1642 vssd vssd vccd vccd net1641 sky130_fd_sc_hd__buf_6
XFILLER_47_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1652 net1653 vssd vssd vccd vccd net1652 sky130_fd_sc_hd__buf_6
XFILLER_46_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1663 net1664 vssd vssd vccd vccd net1663 sky130_fd_sc_hd__buf_6
Xwire1674 net1675 vssd vssd vccd vccd net1674 sky130_fd_sc_hd__buf_6
XFILLER_19_4040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1685 mprj_logic1\[76\] vssd vssd vccd vccd net1685 sky130_fd_sc_hd__buf_6
XFILLER_47_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1696 net1697 vssd vssd vccd vccd net1696 sky130_fd_sc_hd__buf_6
XFILLER_38_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__428__C net86 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ net319 mprj_logic1\[112\] net63 vssd vssd vccd vccd net522 sky130_fd_sc_hd__and3b_4
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__444__B net2180 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_B net1314 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_338_ mprj_logic1\[43\] net1372 vssd vssd vccd vccd net924 sky130_fd_sc_hd__and2_4
XANTENNA_output574_A net574 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_269_ net1778 net139 vssd vssd vccd vccd la_data_in_enable\[106\] sky130_fd_sc_hd__and2_4
Xwire971 la_data_in_mprj_bar\[86\] vssd vssd vccd vccd net971 sky130_fd_sc_hd__buf_6
XFILLER_31_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire982 la_data_in_mprj_bar\[122\] vssd vssd vccd vccd net982 sky130_fd_sc_hd__buf_6
Xwire993 la_data_in_mprj_bar\[100\] vssd vssd vccd vccd net993 sky130_fd_sc_hd__buf_6
XANTENNA_output741_A net1041 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output839_A net839 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1372_A net1373 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] net1328 vssd vssd vccd vccd la_data_in_mprj_bar\[86\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1637_A net1638 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__619__B net1889 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[23\]_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_11 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_22 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_B la_data_in_enable\[105\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__354__B net1377 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_33 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_44 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_55 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_66 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_77 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_88 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_99 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__485__A_N net1590 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2020_A mprj_logic1\[266\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input103_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2118_A mprj_logic1\[183\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__545__A net1559 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__264__B net134 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_123_ mprj_dat_i_core_bar\[9\] vssd vssd vccd vccd net912 sky130_fd_sc_hd__clkinv_2
XFILLER_10_2421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_054_ la_data_in_mprj_bar\[71\] vssd vssd vccd vccd net687 sky130_fd_sc_hd__inv_2
XFILLER_10_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__280__A net1757 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2150 net2151 vssd vssd vccd vccd net2150 sky130_fd_sc_hd__buf_6
XFILLER_1_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2161 mprj_logic1\[158\] vssd vssd vccd vccd net2161 sky130_fd_sc_hd__buf_6
XFILLER_40_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2172 mprj_logic1\[153\] vssd vssd vccd vccd net2172 sky130_fd_sc_hd__buf_6
XFILLER_8_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2183 mprj_logic1\[148\] vssd vssd vccd vccd net2183 sky130_fd_sc_hd__buf_6
XFILLER_5_2780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2194 mprj_logic1\[140\] vssd vssd vccd vccd net2194 sky130_fd_sc_hd__buf_6
XFILLER_47_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1460 net1461 vssd vssd vccd vccd net1460 sky130_fd_sc_hd__buf_6
XFILLER_1_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1471 net404 vssd vssd vccd vccd net1471 sky130_fd_sc_hd__buf_6
XANTENNA__439__B net2189 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1482 net1483 vssd vssd vccd vccd net1482 sky130_fd_sc_hd__buf_6
XFILLER_21_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1493 net398 vssd vssd vccd vccd net1493 sky130_fd_sc_hd__buf_6
XFILLER_47_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1120_A net507 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1218_A net1219 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output691_A net691 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output789_A net789 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[14\]
+ sky130_fd_sc_hd__nand2_2
Xinput20 la_data_out_mprj[114] vssd vssd vccd vccd net20 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput31 la_data_out_mprj[124] vssd vssd vccd vccd net31 sky130_fd_sc_hd__buf_6
XFILLER_50_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput42 la_data_out_mprj[19] vssd vssd vccd vccd net42 sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_out_mprj[29] vssd vssd vccd vccd net53 sky130_fd_sc_hd__clkbuf_4
Xinput64 la_data_out_mprj[39] vssd vssd vccd vccd net64 sky130_fd_sc_hd__clkbuf_4
Xinput75 la_data_out_mprj[49] vssd vssd vccd vccd net75 sky130_fd_sc_hd__clkbuf_4
Xinput86 la_data_out_mprj[59] vssd vssd vccd vccd net86 sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__A net1830 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput97 la_data_out_mprj[69] vssd vssd vccd vccd net97 sky130_fd_sc_hd__buf_6
XFILLER_6_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1921_A mprj_logic1\[315\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] la_data_in_enable\[112\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[112\] sky130_fd_sc_hd__nand2_2
XANTENNA__349__B net1385 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__365__A net1696 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput402 mprj_adr_o_core[22] vssd vssd vccd vccd net402 sky130_fd_sc_hd__buf_6
XFILLER_7_1629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput413 mprj_adr_o_core[3] vssd vssd vccd vccd net413 sky130_fd_sc_hd__buf_6
XFILLER_9_2190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput424 mprj_dat_o_core[12] vssd vssd vccd vccd net424 sky130_fd_sc_hd__buf_6
XFILLER_6_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2068_A mprj_logic1\[201\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput435 mprj_dat_o_core[22] vssd vssd vccd vccd net435 sky130_fd_sc_hd__buf_6
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput446 mprj_dat_o_core[3] vssd vssd vccd vccd net446 sky130_fd_sc_hd__buf_6
XFILLER_2_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput457 mprj_sel_o_core[3] vssd vssd vccd vccd net457 sky130_fd_sc_hd__buf_4
XFILLER_22_3582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input220_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input318_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__A net1767 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_106_ net981 vssd vssd vccd vccd net617 sky130_fd_sc_hd__clkinv_2
XFILLER_51_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput909 net909 vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_8
X_037_ la_data_in_mprj_bar\[54\] vssd vssd vccd vccd net668 sky130_fd_sc_hd__inv_2
XFILLER_45_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__441__C net1632 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output537_A net1092 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1070_A net586 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1168_A net1169 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1290 net1291 vssd vssd vccd vccd net1290 sky130_fd_sc_hd__buf_8
XFILLER_39_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] la_data_in_enable\[49\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[49\] sky130_fd_sc_hd__nand2_2
XFILLER_34_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1502_A net1503 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__185__A net1839 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1871_A mprj_logic1\[330\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1969_A net1970 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__095__A net987 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__542__B mprj_logic1\[247\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input170_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input268_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input435_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput210 la_iena_mprj[55] vssd vssd vccd vccd net210 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input31_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput221 la_iena_mprj[65] vssd vssd vccd vccd net221 sky130_fd_sc_hd__buf_4
XFILLER_23_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput232 la_iena_mprj[75] vssd vssd vccd vccd net232 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput243 la_iena_mprj[85] vssd vssd vccd vccd net243 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput254 la_iena_mprj[95] vssd vssd vccd vccd net254 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput265 la_oenb_mprj[104] vssd vssd vccd vccd net265 sky130_fd_sc_hd__buf_6
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput276 la_oenb_mprj[114] vssd vssd vccd vccd net276 sky130_fd_sc_hd__buf_6
Xinput287 la_oenb_mprj[124] vssd vssd vccd vccd net287 sky130_fd_sc_hd__buf_6
XFILLER_18_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput298 la_oenb_mprj[19] vssd vssd vccd vccd net298 sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_586_ net375 net1976 vssd vssd vccd vccd net834 sky130_fd_sc_hd__and2_2
XFILLER_16_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__C net1337 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output487_A net487 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__452__B net2162 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output654_A net654 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput706 net706 vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_8
Xoutput717 net717 vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_8
XFILLER_29_2821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput728 net728 vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__buf_8
XANTENNA_wire1285_A net1286 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput739 net739 vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__buf_8
XFILLER_42_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output821_A net821 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output919_A net1208 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1452_A net1453 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__362__B net1366 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[6\]_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_440_ net1546 net2188 net1633 vssd vssd vccd vccd net559 sky130_fd_sc_hd__and3b_4
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__419__A_N net333 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_371_ net310 net1684 net54 vssd vssd vccd vccd net513 sky130_fd_sc_hd__and3b_4
XFILLER_18_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2100_A net2101 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__553__A net339 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input385_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__272__B net142 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input79_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__447__B net2173 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1033_A net757 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_569_ net1545 net2010 vssd vssd vccd vccd net816 sky130_fd_sc_hd__and2_4
XFILLER_31_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1200_A net1201 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output771_A net771 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output869_A net869 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput503 net1124 vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__buf_8
XFILLER_9_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput514 net1114 vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__buf_8
XFILLER_44_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1667_A mprj_logic1\[84\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput525 net1104 vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__buf_8
XFILLER_48_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput536 net1093 vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__buf_8
XFILLER_29_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput547 net1080 vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__buf_8
XFILLER_42_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput558 net558 vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__buf_8
Xoutput569 net569 vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1834_A mprj_logic1\[355\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__357__B net1371 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1801 mprj_logic1\[422\] vssd vssd vccd vccd net1801 sky130_fd_sc_hd__buf_4
XFILLER_1_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1812 mprj_logic1\[39\] vssd vssd vccd vccd net1812 sky130_fd_sc_hd__buf_6
Xwire1823 mprj_logic1\[36\] vssd vssd vccd vccd net1823 sky130_fd_sc_hd__buf_6
Xwire1834 mprj_logic1\[355\] vssd vssd vccd vccd net1834 sky130_fd_sc_hd__buf_6
Xwire1845 mprj_logic1\[347\] vssd vssd vccd vccd net1845 sky130_fd_sc_hd__buf_6
XFILLER_19_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input133_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2050_A mprj_logic1\[211\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1856 mprj_logic1\[340\] vssd vssd vccd vccd net1856 sky130_fd_sc_hd__buf_6
XTAP_3101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1867 net1868 vssd vssd vccd vccd net1867 sky130_fd_sc_hd__buf_6
XFILLER_45_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1878 mprj_logic1\[328\] vssd vssd vccd vccd net1878 sky130_fd_sc_hd__buf_6
XANTENNA__548__A net1558 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1889 net1890 vssd vssd vccd vccd net1889 sky130_fd_sc_hd__buf_6
XTAP_3145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_112 mprj_logic1\[261\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input300_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_123 mprj_logic1\[380\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__267__B net137 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 mprj_logic1\[395\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 net1368 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_167 net1512 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ net337 mprj_logic1\[128\] net81 vssd vssd vccd vccd net540 sky130_fd_sc_hd__and3b_4
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_178 net1811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__391__A_N net302 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 net1818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_354_ net1715 net1377 vssd vssd vccd vccd net921 sky130_fd_sc_hd__and2_4
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__283__A net1751 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_285_ net1746 net157 vssd vssd vccd vccd la_data_in_enable\[122\] sky130_fd_sc_hd__and2_4
XFILLER_13_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1246 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1150_A net1151 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput7 la_data_out_mprj[102] vssd vssd vccd vccd net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__177__B net165 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1415_A net1416 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] la_data_in_enable\[31\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[31\] sky130_fd_sc_hd__nand2_2
XFILLER_53_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_138 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__193__A net1826 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1784_A mprj_logic1\[433\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1951_A net1952 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2542 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1108 net520 vssd vssd vccd vccd net1108 sky130_fd_sc_hd__buf_6
XFILLER_5_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1119 net508 vssd vssd vccd vccd net1119 sky130_fd_sc_hd__buf_6
XFILLER_22_3978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__368__A net1690 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_070_ net970 vssd vssd vccd vccd net704 sky130_fd_sc_hd__inv_2
XFILLER_17_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2098_A mprj_logic1\[191\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__550__B mprj_logic1\[255\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input250_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input348_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1620 net114 vssd vssd vccd vccd net1620 sky130_fd_sc_hd__buf_6
XFILLER_1_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1631 net102 vssd vssd vccd vccd net1631 sky130_fd_sc_hd__buf_6
XFILLER_19_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1642 mprj_logic1\[96\] vssd vssd vccd vccd net1642 sky130_fd_sc_hd__buf_6
Xwire1653 mprj_logic1\[90\] vssd vssd vccd vccd net1653 sky130_fd_sc_hd__buf_6
XFILLER_47_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__278__A net1761 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1664 net1665 vssd vssd vccd vccd net1664 sky130_fd_sc_hd__buf_6
XFILLER_24_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1675 mprj_logic1\[80\] vssd vssd vccd vccd net1675 sky130_fd_sc_hd__buf_6
XFILLER_46_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1686 net1687 vssd vssd vccd vccd net1686 sky130_fd_sc_hd__buf_6
Xwire1697 mprj_logic1\[70\] vssd vssd vccd vccd net1697 sky130_fd_sc_hd__buf_6
XFILLER_47_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ net318 mprj_logic1\[111\] net62 vssd vssd vccd vccd net521 sky130_fd_sc_hd__and3b_4
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_337_ mprj_logic1\[42\] net1391 vssd vssd vccd vccd net913 sky130_fd_sc_hd__and2_4
XANTENNA__444__C net1629 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_268_ net1780 net138 vssd vssd vccd vccd la_data_in_enable\[105\] sky130_fd_sc_hd__and2_4
XANTENNA_output567_A net567 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire961 la_data_in_mprj_bar\[99\] vssd vssd vccd vccd net961 sky130_fd_sc_hd__buf_6
XFILLER_28_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire972 la_data_in_mprj_bar\[85\] vssd vssd vccd vccd net972 sky130_fd_sc_hd__buf_6
XFILLER_45_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire983 la_data_in_mprj_bar\[117\] vssd vssd vccd vccd net983 sky130_fd_sc_hd__buf_6
XFILLER_31_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire994 net836 vssd vssd vccd vccd net994 sky130_fd_sc_hd__buf_6
X_199_ mprj_logic1\[366\] net189 vssd vssd vccd vccd la_data_in_enable\[36\] sky130_fd_sc_hd__and2_4
XANTENNA_wire1198_A net1199 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__460__B net2143 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output734_A net734 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1365_A net439 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output901_A net901 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] net1333 vssd vssd vccd vccd la_data_in_mprj_bar\[79\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1532_A net371 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__188__A net1833 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[23\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1999_A net2000 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire985_A la_data_in_mprj_bar\[114\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_12 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_23 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_34 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_45 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_56 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_67 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_78 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_89 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__370__B net1686 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__098__A net984 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[14\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__545__B mprj_logic1\[250\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input298_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_122_ mprj_dat_i_core_bar\[8\] vssd vssd vccd vccd net911 sky130_fd_sc_hd__clkinv_2
XFILLER_11_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__561__A net1553 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_053_ la_data_in_mprj_bar\[70\] vssd vssd vccd vccd net686 sky130_fd_sc_hd__inv_2
XFILLER_27_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__280__B net151 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2140 mprj_logic1\[169\] vssd vssd vccd vccd net2140 sky130_fd_sc_hd__buf_6
Xwire2151 mprj_logic1\[161\] vssd vssd vccd vccd net2151 sky130_fd_sc_hd__buf_6
XFILLER_43_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2162 net2163 vssd vssd vccd vccd net2162 sky130_fd_sc_hd__buf_6
Xwire2173 net2174 vssd vssd vccd vccd net2173 sky130_fd_sc_hd__buf_6
XFILLER_1_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2184 net2185 vssd vssd vccd vccd net2184 sky130_fd_sc_hd__buf_6
Xwire1450 net1451 vssd vssd vccd vccd net1450 sky130_fd_sc_hd__buf_6
XFILLER_5_2792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2195 mprj_logic1\[13\] vssd vssd vccd vccd net2195 sky130_fd_sc_hd__buf_6
Xwire1461 net406 vssd vssd vccd vccd net1461 sky130_fd_sc_hd__buf_6
XFILLER_47_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1472 net1473 vssd vssd vccd vccd net1472 sky130_fd_sc_hd__buf_6
XANTENNA__439__C net1334 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1483 net1484 vssd vssd vccd vccd net1483 sky130_fd_sc_hd__buf_6
XFILLER_1_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1494 net1495 vssd vssd vccd vccd net1494 sky130_fd_sc_hd__buf_6
XFILLER_19_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__455__B net2152 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output684_A net684 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput10 la_data_out_mprj[105] vssd vssd vccd vccd net10 sky130_fd_sc_hd__clkbuf_4
XANTENNA_output851_A net1266 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput21 la_data_out_mprj[115] vssd vssd vccd vccd net21 sky130_fd_sc_hd__buf_4
XFILLER_28_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput32 la_data_out_mprj[125] vssd vssd vccd vccd net32 sky130_fd_sc_hd__buf_6
XFILLER_11_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output949_A net1303 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput43 la_data_out_mprj[1] vssd vssd vccd vccd net43 sky130_fd_sc_hd__clkbuf_4
Xinput54 la_data_out_mprj[2] vssd vssd vccd vccd net54 sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput65 la_data_out_mprj[3] vssd vssd vccd vccd net65 sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1482_A net1483 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput76 la_data_out_mprj[4] vssd vssd vccd vccd net76 sky130_fd_sc_hd__clkbuf_4
Xinput87 la_data_out_mprj[5] vssd vssd vccd vccd net87 sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__B net179 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput98 la_data_out_mprj[6] vssd vssd vccd vccd net98 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1747_A net1748 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] la_data_in_enable\[105\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[105\] sky130_fd_sc_hd__nand2_8
XFILLER_0_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj2_logic_high_inst net953 vccd2_uq0 vssd2_uq0 mprj2_logic_high
XFILLER_11_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__365__B net1363 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__452__A_N net1534 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput403 mprj_adr_o_core[23] vssd vssd vccd vccd net403 sky130_fd_sc_hd__buf_6
XFILLER_44_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput414 mprj_adr_o_core[4] vssd vssd vccd vccd net414 sky130_fd_sc_hd__buf_6
XFILLER_22_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput425 mprj_dat_o_core[13] vssd vssd vccd vccd net425 sky130_fd_sc_hd__buf_6
XFILLER_22_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput436 mprj_dat_o_core[23] vssd vssd vccd vccd net436 sky130_fd_sc_hd__buf_6
XFILLER_40_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput447 mprj_dat_o_core[4] vssd vssd vccd vccd net447 sky130_fd_sc_hd__buf_6
Xinput458 mprj_stb_o_core vssd vssd vccd vccd net458 sky130_fd_sc_hd__buf_6
XFILLER_25_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2130_A net2131 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input213_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_959 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__556__A net342 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__B net146 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__291__A net1732 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_105_ net982 vssd vssd vccd vccd net616 sky130_fd_sc_hd__inv_2
XFILLER_7_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_036_ la_data_in_mprj_bar\[53\] vssd vssd vccd vccd net667 sky130_fd_sc_hd__inv_2
XFILLER_45_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1063_A net467 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1280 net1281 vssd vssd vccd vccd net1280 sky130_fd_sc_hd__buf_8
Xwire1291 net1292 vssd vssd vccd vccd net1291 sky130_fd_sc_hd__buf_6
XANTENNA_wire1230_A net1231 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__475__A_N net1601 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1328_A la_data_in_enable\[86\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__185__B net174 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1697_A mprj_logic1\[70\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1864_A mprj_logic1\[334\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high_inst mprj_logic1\[0\] mprj_logic1\[100\] mprj_logic1\[101\] mprj_logic1\[102\]
+ mprj_logic1\[103\] mprj_logic1\[104\] mprj_logic1\[105\] mprj_logic1\[106\] mprj_logic1\[107\]
+ mprj_logic1\[108\] mprj_logic1\[109\] mprj_logic1\[10\] mprj_logic1\[110\] mprj_logic1\[111\]
+ mprj_logic1\[112\] mprj_logic1\[113\] mprj_logic1\[114\] mprj_logic1\[115\] mprj_logic1\[116\]
+ mprj_logic1\[117\] mprj_logic1\[118\] mprj_logic1\[119\] mprj_logic1\[11\] mprj_logic1\[120\]
+ mprj_logic1\[121\] mprj_logic1\[122\] mprj_logic1\[123\] mprj_logic1\[124\] mprj_logic1\[125\]
+ mprj_logic1\[126\] mprj_logic1\[127\] mprj_logic1\[128\] mprj_logic1\[129\] mprj_logic1\[12\]
+ mprj_logic1\[130\] mprj_logic1\[131\] mprj_logic1\[132\] mprj_logic1\[133\] mprj_logic1\[134\]
+ mprj_logic1\[135\] mprj_logic1\[136\] mprj_logic1\[137\] mprj_logic1\[138\] mprj_logic1\[139\]
+ mprj_logic1\[13\] mprj_logic1\[140\] mprj_logic1\[141\] mprj_logic1\[142\] mprj_logic1\[143\]
+ mprj_logic1\[144\] mprj_logic1\[145\] mprj_logic1\[146\] mprj_logic1\[147\] mprj_logic1\[148\]
+ mprj_logic1\[149\] mprj_logic1\[14\] mprj_logic1\[150\] mprj_logic1\[151\] mprj_logic1\[152\]
+ mprj_logic1\[153\] mprj_logic1\[154\] mprj_logic1\[155\] mprj_logic1\[156\] mprj_logic1\[157\]
+ mprj_logic1\[158\] mprj_logic1\[159\] mprj_logic1\[15\] mprj_logic1\[160\] mprj_logic1\[161\]
+ mprj_logic1\[162\] mprj_logic1\[163\] mprj_logic1\[164\] mprj_logic1\[165\] mprj_logic1\[166\]
+ mprj_logic1\[167\] mprj_logic1\[168\] mprj_logic1\[169\] mprj_logic1\[16\] mprj_logic1\[170\]
+ mprj_logic1\[171\] mprj_logic1\[172\] mprj_logic1\[173\] mprj_logic1\[174\] mprj_logic1\[175\]
+ mprj_logic1\[176\] mprj_logic1\[177\] mprj_logic1\[178\] mprj_logic1\[179\] mprj_logic1\[17\]
+ mprj_logic1\[180\] mprj_logic1\[181\] mprj_logic1\[182\] mprj_logic1\[183\] mprj_logic1\[184\]
+ mprj_logic1\[185\] mprj_logic1\[186\] mprj_logic1\[187\] mprj_logic1\[188\] mprj_logic1\[189\]
+ mprj_logic1\[18\] mprj_logic1\[190\] mprj_logic1\[191\] mprj_logic1\[192\] mprj_logic1\[193\]
+ mprj_logic1\[194\] mprj_logic1\[195\] mprj_logic1\[196\] mprj_logic1\[197\] mprj_logic1\[198\]
+ mprj_logic1\[199\] mprj_logic1\[19\] mprj_logic1\[1\] mprj_logic1\[200\] mprj_logic1\[201\]
+ mprj_logic1\[202\] mprj_logic1\[203\] mprj_logic1\[204\] mprj_logic1\[205\] mprj_logic1\[206\]
+ mprj_logic1\[207\] mprj_logic1\[208\] mprj_logic1\[209\] mprj_logic1\[20\] mprj_logic1\[210\]
+ mprj_logic1\[211\] mprj_logic1\[212\] mprj_logic1\[213\] mprj_logic1\[214\] mprj_logic1\[215\]
+ mprj_logic1\[216\] mprj_logic1\[217\] mprj_logic1\[218\] mprj_logic1\[219\] mprj_logic1\[21\]
+ mprj_logic1\[220\] mprj_logic1\[221\] mprj_logic1\[222\] mprj_logic1\[223\] mprj_logic1\[224\]
+ mprj_logic1\[225\] mprj_logic1\[226\] mprj_logic1\[227\] mprj_logic1\[228\] mprj_logic1\[229\]
+ mprj_logic1\[22\] mprj_logic1\[230\] mprj_logic1\[231\] mprj_logic1\[232\] mprj_logic1\[233\]
+ mprj_logic1\[234\] mprj_logic1\[235\] mprj_logic1\[236\] mprj_logic1\[237\] mprj_logic1\[238\]
+ mprj_logic1\[239\] mprj_logic1\[23\] mprj_logic1\[240\] mprj_logic1\[241\] mprj_logic1\[242\]
+ mprj_logic1\[243\] mprj_logic1\[244\] mprj_logic1\[245\] mprj_logic1\[246\] mprj_logic1\[247\]
+ mprj_logic1\[248\] mprj_logic1\[249\] mprj_logic1\[24\] mprj_logic1\[250\] mprj_logic1\[251\]
+ mprj_logic1\[252\] mprj_logic1\[253\] mprj_logic1\[254\] mprj_logic1\[255\] mprj_logic1\[256\]
+ mprj_logic1\[257\] mprj_logic1\[258\] mprj_logic1\[259\] mprj_logic1\[25\] mprj_logic1\[260\]
+ mprj_logic1\[261\] mprj_logic1\[262\] mprj_logic1\[263\] mprj_logic1\[264\] mprj_logic1\[265\]
+ mprj_logic1\[266\] mprj_logic1\[267\] mprj_logic1\[268\] mprj_logic1\[269\] mprj_logic1\[26\]
+ mprj_logic1\[270\] mprj_logic1\[271\] mprj_logic1\[272\] mprj_logic1\[273\] mprj_logic1\[274\]
+ mprj_logic1\[275\] mprj_logic1\[276\] mprj_logic1\[277\] mprj_logic1\[278\] mprj_logic1\[279\]
+ mprj_logic1\[27\] mprj_logic1\[280\] mprj_logic1\[281\] mprj_logic1\[282\] mprj_logic1\[283\]
+ mprj_logic1\[284\] mprj_logic1\[285\] mprj_logic1\[286\] mprj_logic1\[287\] mprj_logic1\[288\]
+ mprj_logic1\[289\] mprj_logic1\[28\] mprj_logic1\[290\] mprj_logic1\[291\] mprj_logic1\[292\]
+ mprj_logic1\[293\] mprj_logic1\[294\] mprj_logic1\[295\] mprj_logic1\[296\] mprj_logic1\[297\]
+ mprj_logic1\[298\] mprj_logic1\[299\] mprj_logic1\[29\] mprj_logic1\[2\] mprj_logic1\[300\]
+ mprj_logic1\[301\] mprj_logic1\[302\] mprj_logic1\[303\] mprj_logic1\[304\] mprj_logic1\[305\]
+ mprj_logic1\[306\] mprj_logic1\[307\] mprj_logic1\[308\] mprj_logic1\[309\] mprj_logic1\[30\]
+ mprj_logic1\[310\] mprj_logic1\[311\] mprj_logic1\[312\] mprj_logic1\[313\] mprj_logic1\[314\]
+ mprj_logic1\[315\] mprj_logic1\[316\] mprj_logic1\[317\] mprj_logic1\[318\] mprj_logic1\[319\]
+ mprj_logic1\[31\] mprj_logic1\[320\] mprj_logic1\[321\] mprj_logic1\[322\] mprj_logic1\[323\]
+ mprj_logic1\[324\] mprj_logic1\[325\] mprj_logic1\[326\] mprj_logic1\[327\] mprj_logic1\[328\]
+ mprj_logic1\[329\] mprj_logic1\[32\] mprj_logic1\[330\] mprj_logic1\[331\] mprj_logic1\[332\]
+ mprj_logic1\[333\] mprj_logic1\[334\] mprj_logic1\[335\] mprj_logic1\[336\] mprj_logic1\[337\]
+ mprj_logic1\[338\] mprj_logic1\[339\] mprj_logic1\[33\] mprj_logic1\[340\] mprj_logic1\[341\]
+ mprj_logic1\[342\] mprj_logic1\[343\] mprj_logic1\[344\] mprj_logic1\[345\] mprj_logic1\[346\]
+ mprj_logic1\[347\] mprj_logic1\[348\] mprj_logic1\[349\] mprj_logic1\[34\] mprj_logic1\[350\]
+ mprj_logic1\[351\] mprj_logic1\[352\] mprj_logic1\[353\] mprj_logic1\[354\] mprj_logic1\[355\]
+ mprj_logic1\[356\] mprj_logic1\[357\] mprj_logic1\[358\] mprj_logic1\[359\] mprj_logic1\[35\]
+ mprj_logic1\[360\] mprj_logic1\[361\] mprj_logic1\[362\] mprj_logic1\[363\] mprj_logic1\[364\]
+ mprj_logic1\[365\] mprj_logic1\[366\] mprj_logic1\[367\] mprj_logic1\[368\] mprj_logic1\[369\]
+ mprj_logic1\[36\] mprj_logic1\[370\] mprj_logic1\[371\] mprj_logic1\[372\] mprj_logic1\[373\]
+ mprj_logic1\[374\] mprj_logic1\[375\] mprj_logic1\[376\] mprj_logic1\[377\] mprj_logic1\[378\]
+ mprj_logic1\[379\] mprj_logic1\[37\] mprj_logic1\[380\] mprj_logic1\[381\] mprj_logic1\[382\]
+ mprj_logic1\[383\] mprj_logic1\[384\] mprj_logic1\[385\] mprj_logic1\[386\] mprj_logic1\[387\]
+ mprj_logic1\[388\] mprj_logic1\[389\] mprj_logic1\[38\] mprj_logic1\[390\] mprj_logic1\[391\]
+ mprj_logic1\[392\] mprj_logic1\[393\] mprj_logic1\[394\] mprj_logic1\[395\] mprj_logic1\[396\]
+ mprj_logic1\[397\] mprj_logic1\[398\] mprj_logic1\[399\] mprj_logic1\[39\] mprj_logic1\[3\]
+ mprj_logic1\[400\] mprj_logic1\[401\] mprj_logic1\[402\] mprj_logic1\[403\] mprj_logic1\[404\]
+ mprj_logic1\[405\] mprj_logic1\[406\] mprj_logic1\[407\] mprj_logic1\[408\] mprj_logic1\[409\]
+ mprj_logic1\[40\] mprj_logic1\[410\] mprj_logic1\[411\] mprj_logic1\[412\] mprj_logic1\[413\]
+ mprj_logic1\[414\] mprj_logic1\[415\] mprj_logic1\[416\] mprj_logic1\[417\] mprj_logic1\[418\]
+ mprj_logic1\[419\] mprj_logic1\[41\] mprj_logic1\[420\] mprj_logic1\[421\] mprj_logic1\[422\]
+ mprj_logic1\[423\] mprj_logic1\[424\] mprj_logic1\[425\] mprj_logic1\[426\] mprj_logic1\[427\]
+ mprj_logic1\[428\] mprj_logic1\[429\] mprj_logic1\[42\] mprj_logic1\[430\] mprj_logic1\[431\]
+ mprj_logic1\[432\] mprj_logic1\[433\] mprj_logic1\[434\] mprj_logic1\[435\] mprj_logic1\[436\]
+ mprj_logic1\[437\] mprj_logic1\[438\] mprj_logic1\[439\] mprj_logic1\[43\] mprj_logic1\[440\]
+ mprj_logic1\[441\] mprj_logic1\[442\] mprj_logic1\[443\] mprj_logic1\[444\] mprj_logic1\[445\]
+ mprj_logic1\[446\] mprj_logic1\[447\] mprj_logic1\[448\] mprj_logic1\[449\] mprj_logic1\[44\]
+ mprj_logic1\[450\] mprj_logic1\[451\] mprj_logic1\[452\] mprj_logic1\[453\] mprj_logic1\[454\]
+ mprj_logic1\[455\] mprj_logic1\[456\] mprj_logic1\[457\] mprj_logic1\[458\] mprj_logic1\[459\]
+ mprj_logic1\[45\] mprj_logic1\[460\] net951 mprj_logic1\[462\] mprj_logic1\[46\]
+ mprj_logic1\[47\] mprj_logic1\[48\] mprj_logic1\[49\] mprj_logic1\[4\] mprj_logic1\[50\]
+ mprj_logic1\[51\] mprj_logic1\[52\] mprj_logic1\[53\] mprj_logic1\[54\] mprj_logic1\[55\]
+ mprj_logic1\[56\] mprj_logic1\[57\] mprj_logic1\[58\] mprj_logic1\[59\] mprj_logic1\[5\]
+ mprj_logic1\[60\] mprj_logic1\[61\] mprj_logic1\[62\] mprj_logic1\[63\] mprj_logic1\[64\]
+ mprj_logic1\[65\] mprj_logic1\[66\] mprj_logic1\[67\] mprj_logic1\[68\] mprj_logic1\[69\]
+ mprj_logic1\[6\] mprj_logic1\[70\] mprj_logic1\[71\] mprj_logic1\[72\] mprj_logic1\[73\]
+ mprj_logic1\[74\] mprj_logic1\[75\] mprj_logic1\[76\] mprj_logic1\[77\] mprj_logic1\[78\]
+ mprj_logic1\[79\] mprj_logic1\[7\] mprj_logic1\[80\] mprj_logic1\[81\] mprj_logic1\[82\]
+ mprj_logic1\[83\] mprj_logic1\[84\] mprj_logic1\[85\] mprj_logic1\[86\] mprj_logic1\[87\]
+ mprj_logic1\[88\] mprj_logic1\[89\] mprj_logic1\[8\] mprj_logic1\[90\] mprj_logic1\[91\]
+ mprj_logic1\[92\] mprj_logic1\[93\] mprj_logic1\[94\] mprj_logic1\[95\] mprj_logic1\[96\]
+ mprj_logic1\[97\] mprj_logic1\[98\] mprj_logic1\[99\] mprj_logic1\[9\] vccd1_uq1
+ vssd1_uq1 mprj_logic_high
XTAP_3508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2080_A net2081 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input163_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2178_A mprj_logic1\[150\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput200 la_iena_mprj[46] vssd vssd vccd vccd net200 sky130_fd_sc_hd__buf_4
Xinput211 la_iena_mprj[56] vssd vssd vccd vccd net211 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput222 la_iena_mprj[66] vssd vssd vccd vccd net222 sky130_fd_sc_hd__buf_4
XFILLER_0_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput233 la_iena_mprj[76] vssd vssd vccd vccd net233 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input330_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput244 la_iena_mprj[86] vssd vssd vccd vccd net244 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input428_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput255 la_iena_mprj[96] vssd vssd vccd vccd net255 sky130_fd_sc_hd__clkbuf_4
Xinput266 la_oenb_mprj[105] vssd vssd vccd vccd net266 sky130_fd_sc_hd__buf_6
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input24_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput277 la_oenb_mprj[115] vssd vssd vccd vccd net277 sky130_fd_sc_hd__buf_6
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput288 la_oenb_mprj[125] vssd vssd vccd vccd net288 sky130_fd_sc_hd__buf_6
Xinput299 la_oenb_mprj[1] vssd vssd vccd vccd net299 sky130_fd_sc_hd__buf_4
XFILLER_18_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__286__A net1744 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_585_ net1529 net1977 vssd vssd vccd vccd net833 sky130_fd_sc_hd__and2_4
XFILLER_17_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__452__C net1621 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput707 net707 vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_8
Xoutput718 net718 vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_8
XFILLER_10_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput729 net729 vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__buf_8
XANTENNA_output647_A net647 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_019_ la_data_in_mprj_bar\[36\] vssd vssd vccd vccd net648 sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1180_A net1181 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1278_A net1279 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output814_A net814 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1445_A net1446 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] la_data_in_enable\[61\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[61\] sky130_fd_sc_hd__nand2_2
XFILLER_23_2498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__196__A mprj_logic1\[363\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1981_A net1982 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[6\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ net299 net1686 net43 vssd vssd vccd vccd net502 sky130_fd_sc_hd__and3b_4
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__553__B mprj_logic1\[258\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input280_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input378_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_542 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__447__C net1626 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_568_ net1546 net2012 vssd vssd vccd vccd net815 sky130_fd_sc_hd__and2_4
XANTENNA_wire1026_A net765 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output597_A net597 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2578 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_499_ net310 net2060 vssd vssd vccd vccd net769 sky130_fd_sc_hd__and2_4
XFILLER_31_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__B net2141 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output764_A net1027 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1395_A net1396 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput504 net1123 vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__buf_8
XANTENNA_output931_A net1166 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput515 net1113 vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__buf_8
XFILLER_44_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput526 net1103 vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__buf_8
Xoutput537 net1092 vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__buf_8
Xoutput548 net1079 vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__buf_8
XFILLER_47_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput559 net559 vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__buf_8
XFILLER_25_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1827_A mprj_logic1\[35\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__373__B net1680 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1802 mprj_logic1\[421\] vssd vssd vccd vccd net1802 sky130_fd_sc_hd__buf_6
XFILLER_5_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1813 mprj_logic1\[399\] vssd vssd vccd vccd net1813 sky130_fd_sc_hd__buf_6
Xwire1824 mprj_logic1\[362\] vssd vssd vccd vccd net1824 sky130_fd_sc_hd__buf_4
XFILLER_41_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1835 net1836 vssd vssd vccd vccd net1835 sky130_fd_sc_hd__buf_6
Xwire1846 mprj_logic1\[346\] vssd vssd vccd vccd net1846 sky130_fd_sc_hd__buf_6
XTAP_3102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1857 mprj_logic1\[339\] vssd vssd vccd vccd net1857 sky130_fd_sc_hd__buf_6
XFILLER_24_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1868 mprj_logic1\[332\] vssd vssd vccd vccd net1868 sky130_fd_sc_hd__buf_6
XFILLER_41_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1879 net1880 vssd vssd vccd vccd net1879 sky130_fd_sc_hd__buf_6
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__548__B mprj_logic1\[253\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2043_A mprj_logic1\[215\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_113 mprj_logic1\[261\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_124 mprj_logic1\[382\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_135 mprj_logic1\[395\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_422_ net336 mprj_logic1\[127\] net80 vssd vssd vccd vccd net539 sky130_fd_sc_hd__and3b_4
XANTENNA_157 net1368 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 net1555 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 net1811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__564__A net1550 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ net1716 net1378 vssd vssd vccd vccd net920 sky130_fd_sc_hd__and2_4
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input91_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_284_ net1749 net156 vssd vssd vccd vccd la_data_in_enable\[121\] sky130_fd_sc_hd__and2_4
XFILLER_52_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[7\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1258 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output512_A net1115 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput8 la_data_out_mprj[103] vssd vssd vccd vccd net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__458__B net2145 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1143_A net513 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1408_A net417 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_36_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] la_data_in_enable\[24\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[24\] sky130_fd_sc_hd__nand2_4
XFILLER_53_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__193__B net183 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1777_A mprj_logic1\[437\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1944_A mprj_logic1\[306\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__409__A_N net322 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1109 net519 vssd vssd vccd vccd net1109 sky130_fd_sc_hd__buf_6
XFILLER_5_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__368__B net1358 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_14_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput890 net890 vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_8
XFILLER_43_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2160_A net2161 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input243_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1610 net223 vssd vssd vccd vccd net1610 sky130_fd_sc_hd__buf_4
XANTENNA__559__A net1555 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1621 net113 vssd vssd vccd vccd net1621 sky130_fd_sc_hd__buf_6
XFILLER_4_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1632 net101 vssd vssd vccd vccd net1632 sky130_fd_sc_hd__buf_6
Xwire1643 net1644 vssd vssd vccd vccd net1643 sky130_fd_sc_hd__buf_6
XFILLER_46_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1654 mprj_logic1\[8\] vssd vssd vccd vccd net1654 sky130_fd_sc_hd__buf_6
XANTENNA_input410_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__278__B net149 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1665 mprj_logic1\[85\] vssd vssd vccd vccd net1665 sky130_fd_sc_hd__buf_6
Xwire1676 net1677 vssd vssd vccd vccd net1676 sky130_fd_sc_hd__buf_6
XFILLER_46_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1687 mprj_logic1\[75\] vssd vssd vccd vccd net1687 sky130_fd_sc_hd__buf_6
XFILLER_34_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1698 net1699 vssd vssd vccd vccd net1698 sky130_fd_sc_hd__buf_6
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__294__A net1720 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_405_ net317 mprj_logic1\[110\] net61 vssd vssd vccd vccd net520 sky130_fd_sc_hd__and3b_4
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_336_ net1803 net1427 vssd vssd vccd vccd net872 sky130_fd_sc_hd__and2_4
XFILLER_10_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_267_ net1782 net137 vssd vssd vccd vccd la_data_in_enable\[104\] sky130_fd_sc_hd__and2_4
Xwire962 la_data_in_mprj_bar\[95\] vssd vssd vccd vccd net962 sky130_fd_sc_hd__buf_6
XFILLER_10_3883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire973 la_data_in_mprj_bar\[84\] vssd vssd vccd vccd net973 sky130_fd_sc_hd__buf_6
X_198_ mprj_logic1\[365\] net188 vssd vssd vccd vccd la_data_in_enable\[35\] sky130_fd_sc_hd__and2_2
Xwire984 la_data_in_mprj_bar\[115\] vssd vssd vccd vccd net984 sky130_fd_sc_hd__buf_6
XFILLER_45_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire995 net834 vssd vssd vccd vccd net995 sky130_fd_sc_hd__buf_6
XFILLER_26_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__460__C net122 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1093_A net1094 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output727_A net727 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1358_A net445 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__188__B net1613 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1525_A net1526 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1894_A mprj_logic1\[323\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_13 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_24 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_35 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_46 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_57 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_68 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_79 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__C net43 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__381__A_N net291 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2006_A mprj_logic1\[277\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_121_ mprj_dat_i_core_bar\[7\] vssd vssd vccd vccd net910 sky130_fd_sc_hd__clkinv_2
XFILLER_49_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input193_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_052_ la_data_in_mprj_bar\[69\] vssd vssd vccd vccd net684 sky130_fd_sc_hd__inv_2
XANTENNA__561__B net2020 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input360_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input458_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input54_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2130 net2131 vssd vssd vccd vccd net2130 sky130_fd_sc_hd__buf_6
XFILLER_21_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2141 mprj_logic1\[168\] vssd vssd vccd vccd net2141 sky130_fd_sc_hd__buf_6
XANTENNA__289__A net1738 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2152 net2153 vssd vssd vccd vccd net2152 sky130_fd_sc_hd__buf_6
XFILLER_38_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2163 net2164 vssd vssd vccd vccd net2163 sky130_fd_sc_hd__buf_6
Xwire2174 mprj_logic1\[152\] vssd vssd vccd vccd net2174 sky130_fd_sc_hd__buf_6
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1440 net1441 vssd vssd vccd vccd net1440 sky130_fd_sc_hd__buf_6
Xwire2185 mprj_logic1\[147\] vssd vssd vccd vccd net2185 sky130_fd_sc_hd__buf_6
XFILLER_1_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1451 net408 vssd vssd vccd vccd net1451 sky130_fd_sc_hd__buf_6
XFILLER_21_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2196 mprj_logic1\[139\] vssd vssd vccd vccd net2196 sky130_fd_sc_hd__buf_6
XFILLER_4_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1462 net1463 vssd vssd vccd vccd net1462 sky130_fd_sc_hd__buf_8
XFILLER_21_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1473 net1474 vssd vssd vccd vccd net1473 sky130_fd_sc_hd__buf_6
XFILLER_1_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1484 net400 vssd vssd vccd vccd net1484 sky130_fd_sc_hd__buf_6
XFILLER_46_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1495 net1496 vssd vssd vccd vccd net1495 sky130_fd_sc_hd__buf_6
Xpowergood_check vccd vssd vdda1_uq0 vssa1_uq0 vdda2_uq0 vssa2_uq0 net954 net952 mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__455__C net1618 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1106_A net522 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_319_ mprj_logic1\[24\] net1509 vssd vssd vccd vccd net853 sky130_fd_sc_hd__and2_2
XFILLER_50_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput11 la_data_out_mprj[106] vssd vssd vccd vccd net11 sky130_fd_sc_hd__clkbuf_4
Xinput22 la_data_out_mprj[116] vssd vssd vccd vccd net22 sky130_fd_sc_hd__clkbuf_4
Xinput33 la_data_out_mprj[126] vssd vssd vccd vccd net33 sky130_fd_sc_hd__buf_6
XANTENNA__471__B net2130 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput44 la_data_out_mprj[20] vssd vssd vccd vccd net44 sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_out_mprj[30] vssd vssd vccd vccd net55 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output844_A net844 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput66 la_data_out_mprj[40] vssd vssd vccd vccd net66 sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_mprj[50] vssd vssd vccd vccd net77 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput88 la_data_out_mprj[60] vssd vssd vccd vccd net88 sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_mprj[70] vssd vssd vccd vccd net99 sky130_fd_sc_hd__buf_6
XFILLER_28_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1475_A net1476 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] net1323 vssd vssd vccd vccd la_data_in_mprj_bar\[91\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1642_A mprj_logic1\[96\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__199__A mprj_logic1\[366\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1907_A mprj_logic1\[319\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__B net1661 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput404 mprj_adr_o_core[24] vssd vssd vccd vccd net404 sky130_fd_sc_hd__buf_6
XFILLER_40_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput415 mprj_adr_o_core[5] vssd vssd vccd vccd net415 sky130_fd_sc_hd__buf_6
XFILLER_44_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput426 mprj_dat_o_core[14] vssd vssd vccd vccd net426 sky130_fd_sc_hd__buf_6
XFILLER_6_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput437 mprj_dat_o_core[24] vssd vssd vccd vccd net437 sky130_fd_sc_hd__buf_6
XFILLER_40_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput448 mprj_dat_o_core[5] vssd vssd vccd vccd net448 sky130_fd_sc_hd__buf_6
Xinput459 mprj_we_o_core vssd vssd vccd vccd net459 sky130_fd_sc_hd__buf_6
XFILLER_29_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_798 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2123_A mprj_logic1\[180\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input206_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__572__A net1542 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_104_ la_data_in_mprj_bar\[121\] vssd vssd vccd vccd net615 sky130_fd_sc_hd__clkinv_2
XFILLER_8_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__291__B net460 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_035_ la_data_in_mprj_bar\[52\] vssd vssd vccd vccd net666 sky130_fd_sc_hd__inv_2
XFILLER_10_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1056_A net475 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1270 net850 vssd vssd vccd vccd net1270 sky130_fd_sc_hd__buf_6
Xwire1281 net1282 vssd vssd vccd vccd net1281 sky130_fd_sc_hd__buf_6
XFILLER_19_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1292 net1293 vssd vssd vccd vccd net1292 sky130_fd_sc_hd__buf_6
XFILLER_19_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__466__B net2137 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1223_A net1224 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A net1007 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1857_A mprj_logic1\[339\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__376__B net1672 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B net1318 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2073_A net2074 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input156_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput201 la_iena_mprj[47] vssd vssd vccd vccd net201 sky130_fd_sc_hd__buf_4
XFILLER_27_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput212 la_iena_mprj[57] vssd vssd vccd vccd net212 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput223 la_iena_mprj[67] vssd vssd vccd vccd net223 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput234 la_iena_mprj[77] vssd vssd vccd vccd net234 sky130_fd_sc_hd__clkbuf_4
XTAP_4711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 la_iena_mprj[87] vssd vssd vccd vccd net245 sky130_fd_sc_hd__clkbuf_4
Xinput256 la_iena_mprj[97] vssd vssd vccd vccd net256 sky130_fd_sc_hd__buf_4
XFILLER_2_3453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput267 la_oenb_mprj[106] vssd vssd vccd vccd net267 sky130_fd_sc_hd__buf_6
XANTENNA_input323_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput278 la_oenb_mprj[116] vssd vssd vccd vccd net278 sky130_fd_sc_hd__buf_6
Xinput289 la_oenb_mprj[126] vssd vssd vccd vccd net289 sky130_fd_sc_hd__buf_6
XANTENNA__567__A net1547 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input17_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__286__B net158 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_584_ net1530 net1979 vssd vssd vccd vccd net832 sky130_fd_sc_hd__and2_4
XFILLER_16_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_B net1327 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput708 net708 vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_8
Xoutput719 net1053 vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__buf_8
X_018_ la_data_in_mprj_bar\[35\] vssd vssd vccd vccd net647 sky130_fd_sc_hd__inv_2
XANTENNA_output542_A net1085 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1173_A net930 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_B la_data_in_enable\[11\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_42_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__442__A_N net1544 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output807_A net807 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1438_A net1439 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] la_data_in_enable\[54\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[54\] sky130_fd_sc_hd__nand2_2
XFILLER_1_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_B la_data_in_enable\[78\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_53_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1974_A mprj_logic1\[293\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input9_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input273_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__465__A_N net383 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input440_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__297__A net1959 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_567_ net1547 net2014 vssd vssd vccd vccd net814 sky130_fd_sc_hd__and2_4
XFILLER_53_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_498_ net299 net2062 vssd vssd vccd vccd net758 sky130_fd_sc_hd__and2_4
XANTENNA_output492_A net492 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1019_A net779 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__C net125 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output757_A net1033 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1290_A net1291 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput505 net1122 vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__buf_8
Xoutput516 net1112 vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__buf_8
Xoutput527 net1102 vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__buf_8
XFILLER_29_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput538 net1091 vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__buf_8
XANTENNA_output924_A net1249 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput549 net1078 vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__buf_8
XFILLER_42_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1722_A mprj_logic1\[462\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__000__A la_data_in_mprj_bar\[17\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__488__A_N net1587 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1803 mprj_logic1\[41\] vssd vssd vccd vccd net1803 sky130_fd_sc_hd__buf_6
Xwire1814 mprj_logic1\[398\] vssd vssd vccd vccd net1814 sky130_fd_sc_hd__buf_6
XFILLER_4_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1825 mprj_logic1\[361\] vssd vssd vccd vccd net1825 sky130_fd_sc_hd__buf_6
Xwire1836 mprj_logic1\[354\] vssd vssd vccd vccd net1836 sky130_fd_sc_hd__buf_6
XFILLER_3_3570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1847 net1848 vssd vssd vccd vccd net1847 sky130_fd_sc_hd__buf_6
XTAP_3103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1858 mprj_logic1\[338\] vssd vssd vccd vccd net1858 sky130_fd_sc_hd__buf_6
XTAP_3114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1869 net1870 vssd vssd vccd vccd net1869 sky130_fd_sc_hd__buf_6
XFILLER_18_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 mprj_logic1\[383\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2036_A mprj_logic1\[219\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_421_ net335 mprj_logic1\[126\] net79 vssd vssd vccd vccd net538 sky130_fd_sc_hd__and3b_4
XANTENNA_136 mprj_logic1\[395\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_147 mprj_logic1\[46\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 net1368 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 net1575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__564__B net2017 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_352_ net1717 net1379 vssd vssd vccd vccd net919 sky130_fd_sc_hd__and2_4
XFILLER_32_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[126\]_B la_data_in_enable\[126\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2203_A net2204 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_283_ net1751 net155 vssd vssd vccd vccd la_data_in_enable\[120\] sky130_fd_sc_hd__and2_4
XFILLER_35_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input390_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input84_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__580__A net1534 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput9 la_data_out_mprj[104] vssd vssd vccd vccd net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__458__C net119 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output505_A net1122 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1136_A net590 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_619_ net1584 net1889 vssd vssd vccd vccd net744 sky130_fd_sc_hd__and2_4
XFILLER_17_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__B net2124 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[117\]_B la_data_in_enable\[117\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_wire1303_A net1304 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] la_data_in_enable\[17\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[17\] sky130_fd_sc_hd__nand2_4
XFILLER_11_3829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1672_A net1673 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1937_A net1938 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__B net1655 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B la_data_in_enable\[108\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput880 net1306 vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__buf_8
Xoutput891 net891 vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_8
XFILLER_5_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1600 net268 vssd vssd vccd vccd net1600 sky130_fd_sc_hd__buf_6
Xwire1611 net22 vssd vssd vccd vccd net1611 sky130_fd_sc_hd__buf_4
XFILLER_21_3446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__559__B net2022 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1622 net112 vssd vssd vccd vccd net1622 sky130_fd_sc_hd__buf_6
XANTENNA_input236_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2153_A net2154 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[17\]_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1633 net100 vssd vssd vccd vccd net1633 sky130_fd_sc_hd__buf_4
XFILLER_4_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1644 mprj_logic1\[95\] vssd vssd vccd vccd net1644 sky130_fd_sc_hd__buf_6
XFILLER_41_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1655 net1656 vssd vssd vccd vccd net1655 sky130_fd_sc_hd__buf_6
XFILLER_24_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1666 net1667 vssd vssd vccd vccd net1666 sky130_fd_sc_hd__buf_6
XFILLER_19_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1677 mprj_logic1\[7\] vssd vssd vccd vccd net1677 sky130_fd_sc_hd__buf_6
Xwire1688 net1689 vssd vssd vccd vccd net1688 sky130_fd_sc_hd__buf_6
XFILLER_41_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1699 mprj_logic1\[6\] vssd vssd vccd vccd net1699 sky130_fd_sc_hd__buf_6
XANTENNA_input403_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__A net1539 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__294__B net453 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_404_ net1569 mprj_logic1\[109\] net60 vssd vssd vccd vccd net519 sky130_fd_sc_hd__and3b_4
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_335_ net1809 net1432 vssd vssd vccd vccd net871 sky130_fd_sc_hd__and2_4
XFILLER_30_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_266_ net1784 net136 vssd vssd vccd vccd la_data_in_enable\[103\] sky130_fd_sc_hd__and2_2
XFILLER_10_3840 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire963 la_data_in_mprj_bar\[94\] vssd vssd vccd vccd net963 sky130_fd_sc_hd__buf_6
XFILLER_26_4003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_197_ mprj_logic1\[364\] net187 vssd vssd vccd vccd la_data_in_enable\[34\] sky130_fd_sc_hd__and2_2
Xwire974 la_data_in_mprj_bar\[83\] vssd vssd vccd vccd net974 sky130_fd_sc_hd__buf_6
Xwire985 la_data_in_mprj_bar\[114\] vssd vssd vccd vccd net985 sky130_fd_sc_hd__buf_6
XFILLER_48_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire996 net804 vssd vssd vccd vccd net996 sky130_fd_sc_hd__buf_6
XFILLER_26_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__B net2133 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1253_A net863 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_936 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1420_A net1421 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1518_A net1519 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_14 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_25 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1887_A net1888 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_36 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_47 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_58 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_69 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__379__B net1666 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_120_ mprj_dat_i_core_bar\[6\] vssd vssd vccd vccd net909 sky130_fd_sc_hd__clkinv_2
XFILLER_10_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_051_ la_data_in_mprj_bar\[68\] vssd vssd vccd vccd net683 sky130_fd_sc_hd__inv_2
XFILLER_49_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input186_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input353_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input47_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2120 mprj_logic1\[182\] vssd vssd vccd vccd net2120 sky130_fd_sc_hd__buf_6
XFILLER_1_4027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2131 mprj_logic1\[176\] vssd vssd vccd vccd net2131 sky130_fd_sc_hd__buf_6
XANTENNA__289__B net161 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2142 mprj_logic1\[166\] vssd vssd vccd vccd net2142 sky130_fd_sc_hd__buf_6
XFILLER_5_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2153 net2154 vssd vssd vccd vccd net2153 sky130_fd_sc_hd__buf_6
Xwire2164 mprj_logic1\[157\] vssd vssd vccd vccd net2164 sky130_fd_sc_hd__buf_6
Xwire1430 net1431 vssd vssd vccd vccd net1430 sky130_fd_sc_hd__buf_6
Xwire2175 net2176 vssd vssd vccd vccd net2175 sky130_fd_sc_hd__buf_6
Xwire1441 net410 vssd vssd vccd vccd net1441 sky130_fd_sc_hd__buf_6
XFILLER_1_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2186 net2187 vssd vssd vccd vccd net2186 sky130_fd_sc_hd__buf_6
Xwire1452 net1453 vssd vssd vccd vccd net1452 sky130_fd_sc_hd__buf_8
Xwire2197 mprj_logic1\[138\] vssd vssd vccd vccd net2197 sky130_fd_sc_hd__buf_6
XFILLER_46_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1463 net1464 vssd vssd vccd vccd net1463 sky130_fd_sc_hd__buf_6
Xwire1474 net403 vssd vssd vccd vccd net1474 sky130_fd_sc_hd__buf_6
Xwire1485 net1486 vssd vssd vccd vccd net1485 sky130_fd_sc_hd__buf_6
XFILLER_47_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1496 net1497 vssd vssd vccd vccd net1496 sky130_fd_sc_hd__buf_6
XFILLER_46_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_318_ mprj_logic1\[23\] net1512 vssd vssd vccd vccd net852 sky130_fd_sc_hd__and2_4
XANTENNA_wire1001_A net800 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output572_A net572 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_mprj[107] vssd vssd vccd vccd net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput23 la_data_out_mprj[117] vssd vssd vccd vccd net23 sky130_fd_sc_hd__clkbuf_4
Xinput34 la_data_out_mprj[127] vssd vssd vccd vccd net34 sky130_fd_sc_hd__clkbuf_4
Xinput45 la_data_out_mprj[21] vssd vssd vccd vccd net45 sky130_fd_sc_hd__clkbuf_4
XANTENNA__471__C net7 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_249_ net1806 net244 vssd vssd vccd vccd la_data_in_enable\[86\] sky130_fd_sc_hd__and2_4
XFILLER_45_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput56 la_data_out_mprj[31] vssd vssd vccd vccd net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput67 la_data_out_mprj[41] vssd vssd vccd vccd net67 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput78 la_data_out_mprj[51] vssd vssd vccd vccd net78 sky130_fd_sc_hd__clkbuf_4
Xinput89 la_data_out_mprj[61] vssd vssd vccd vccd net89 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output837_A net837 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1370_A net434 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1468_A net1469 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] net1330 vssd vssd vccd vccd la_data_in_mprj_bar\[84\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__199__B net189 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1635_A net1636 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__C net35 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput405 mprj_adr_o_core[25] vssd vssd vccd vccd net405 sky130_fd_sc_hd__buf_6
XFILLER_40_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput416 mprj_adr_o_core[6] vssd vssd vccd vccd net416 sky130_fd_sc_hd__buf_6
XFILLER_2_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput427 mprj_dat_o_core[15] vssd vssd vccd vccd net427 sky130_fd_sc_hd__buf_6
XFILLER_44_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput438 mprj_dat_o_core[25] vssd vssd vccd vccd net438 sky130_fd_sc_hd__buf_6
Xinput449 mprj_dat_o_core[6] vssd vssd vccd vccd net449 sky130_fd_sc_hd__buf_6
XFILLER_2_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input101_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__572__B net2005 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_103_ la_data_in_mprj_bar\[120\] vssd vssd vccd vccd net614 sky130_fd_sc_hd__inv_2
XFILLER_7_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_034_ la_data_in_mprj_bar\[51\] vssd vssd vccd vccd net665 sky130_fd_sc_hd__clkinv_2
XFILLER_7_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1260 net855 vssd vssd vccd vccd net1260 sky130_fd_sc_hd__buf_6
XFILLER_1_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1271 net1272 vssd vssd vccd vccd net1271 sky130_fd_sc_hd__buf_6
XFILLER_40_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1282 net1283 vssd vssd vccd vccd net1282 sky130_fd_sc_hd__buf_6
XFILLER_1_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1293 net946 vssd vssd vccd vccd net1293 sky130_fd_sc_hd__buf_6
XFILLER_47_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1049_A net791 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__466__C net128 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1216_A net917 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output787_A net787 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__371__A_N net310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__B net2108 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output954_A net954 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[12\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_12_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1752_A mprj_logic1\[450\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] la_data_in_enable\[110\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[110\] sky130_fd_sc_hd__nand2_2
XFILLER_27_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__B net1639 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput202 la_iena_mprj[48] vssd vssd vccd vccd net202 sky130_fd_sc_hd__clkbuf_4
Xinput213 la_iena_mprj[58] vssd vssd vccd vccd net213 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput224 la_iena_mprj[68] vssd vssd vccd vccd net224 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input149_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2066_A net2067 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput235 la_iena_mprj[78] vssd vssd vccd vccd net235 sky130_fd_sc_hd__clkbuf_4
XTAP_4712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 la_iena_mprj[88] vssd vssd vccd vccd net246 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput257 la_iena_mprj[98] vssd vssd vccd vccd net257 sky130_fd_sc_hd__buf_4
Xinput268 la_oenb_mprj[107] vssd vssd vccd vccd net268 sky130_fd_sc_hd__buf_6
XFILLER_40_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput279 la_oenb_mprj[117] vssd vssd vccd vccd net279 sky130_fd_sc_hd__buf_6
XFILLER_18_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__567__B net2014 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input316_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_583_ net1531 net1981 vssd vssd vccd vccd net831 sky130_fd_sc_hd__and2_4
XFILLER_35_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__A_N net305 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__A net1531 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput709 net709 vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_8
XFILLER_7_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_017_ la_data_in_mprj_bar\[34\] vssd vssd vccd vccd net646 sky130_fd_sc_hd__inv_2
XFILLER_46_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output535_A net1141 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1166_A net1167 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__477__B net2119 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1090 net539 vssd vssd vccd vccd net1090 sky130_fd_sc_hd__buf_6
XFILLER_47_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] la_data_in_enable\[47\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[47\] sky130_fd_sc_hd__nand2_2
XFILLER_1_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1967_A net1968 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] la_data_in_enable\[9\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[9\] sky130_fd_sc_hd__nand2_4
XFILLER_28_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__387__B net1648 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2183_A mprj_logic1\[148\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input266_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input433_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__578__A net1536 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_566_ net1548 net2015 vssd vssd vccd vccd net812 sky130_fd_sc_hd__and2_4
XFILLER_32_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_497_ net260 net2064 vssd vssd vccd vccd net719 sky130_fd_sc_hd__and2_4
XFILLER_32_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output485_A net1133 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput506 net1121 vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__buf_8
XFILLER_9_3427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput517 net1111 vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__buf_8
Xoutput528 net1101 vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__buf_8
XANTENNA_wire1283_A net948 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput539 net1090 vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__buf_8
XFILLER_10_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output917_A net1214 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1450_A net1451 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1715_A mprj_logic1\[59\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1804 mprj_logic1\[418\] vssd vssd vccd vccd net1804 sky130_fd_sc_hd__buf_6
Xwire1815 mprj_logic1\[397\] vssd vssd vccd vccd net1815 sky130_fd_sc_hd__buf_6
XFILLER_41_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1826 mprj_logic1\[360\] vssd vssd vccd vccd net1826 sky130_fd_sc_hd__buf_6
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1837 net1838 vssd vssd vccd vccd net1837 sky130_fd_sc_hd__buf_6
XFILLER_24_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1848 mprj_logic1\[345\] vssd vssd vccd vccd net1848 sky130_fd_sc_hd__buf_6
XTAP_3104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1859 net1860 vssd vssd vccd vccd net1859 sky130_fd_sc_hd__buf_6
XTAP_3115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_104 mprj_logic1\[232\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 mprj_logic1\[387\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ net334 mprj_logic1\[125\] net78 vssd vssd vccd vccd net537 sky130_fd_sc_hd__and3b_4
XANTENNA_137 mprj_logic1\[395\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 net18 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 net1370 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2029_A mprj_logic1\[226\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_351_ net1718 net1381 vssd vssd vccd vccd net918 sky130_fd_sc_hd__and2_4
XFILLER_42_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_282_ net1753 net153 vssd vssd vccd vccd la_data_in_enable\[119\] sky130_fd_sc_hd__and2_4
XANTENNA__432__A_N net1554 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input383_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__580__B net1988 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input77_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__101__A la_data_in_mprj_bar\[118\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ net1585 net1892 vssd vssd vccd vccd net743 sky130_fd_sc_hd__and2_4
XTAP_3693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1031_A net760 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1129_A net497 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ net335 mprj_logic1\[254\] vssd vssd vccd vccd net794 sky130_fd_sc_hd__and2_2
XFILLER_32_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output867_A net867 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1498_A net1499 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__B net2085 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1832_A mprj_logic1\[356\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[26\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__455__A_N net1531 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__C net38 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput870 net870 vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_5_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput881 net881 vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_8
XFILLER_1_4209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput892 net892 vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_8
XFILLER_21_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1601 net267 vssd vssd vccd vccd net1601 sky130_fd_sc_hd__buf_6
XFILLER_5_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1612 net178 vssd vssd vccd vccd net1612 sky130_fd_sc_hd__buf_6
XFILLER_21_3458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1623 net111 vssd vssd vccd vccd net1623 sky130_fd_sc_hd__buf_6
XFILLER_8_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[17\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1634 mprj_logic1\[9\] vssd vssd vccd vccd net1634 sky130_fd_sc_hd__buf_6
XFILLER_41_2161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1645 mprj_logic1\[94\] vssd vssd vccd vccd net1645 sky130_fd_sc_hd__buf_6
XANTENNA_input131_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1656 mprj_logic1\[89\] vssd vssd vccd vccd net1656 sky130_fd_sc_hd__buf_6
XANTENNA_wire2146_A net2147 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1667 mprj_logic1\[84\] vssd vssd vccd vccd net1667 sky130_fd_sc_hd__buf_6
XANTENNA_input229_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1678 net1679 vssd vssd vccd vccd net1678 sky130_fd_sc_hd__buf_6
Xwire1689 mprj_logic1\[74\] vssd vssd vccd vccd net1689 sky130_fd_sc_hd__buf_6
XFILLER_34_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__B net1998 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ net315 mprj_logic1\[108\] net59 vssd vssd vccd vccd net518 sky130_fd_sc_hd__and3b_4
XFILLER_26_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ net1812 net1442 vssd vssd vccd vccd net869 sky130_fd_sc_hd__and2_4
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__591__A net381 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_265_ net1785 net135 vssd vssd vccd vccd la_data_in_enable\[102\] sky130_fd_sc_hd__and2_4
XFILLER_10_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire964 la_data_in_mprj_bar\[93\] vssd vssd vccd vccd net964 sky130_fd_sc_hd__buf_6
X_196_ mprj_logic1\[363\] net186 vssd vssd vccd vccd la_data_in_enable\[33\] sky130_fd_sc_hd__and2_4
Xwire975 la_data_in_mprj_bar\[81\] vssd vssd vccd vccd net975 sky130_fd_sc_hd__buf_6
XFILLER_41_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire986 la_data_in_mprj_bar\[113\] vssd vssd vccd vccd net986 sky130_fd_sc_hd__buf_6
Xwire997 net998 vssd vssd vccd vccd net997 sky130_fd_sc_hd__buf_6
XFILLER_48_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1079_A net548 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__469__C net5 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1246_A net1247 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__478__A_N net270 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__485__B net2099 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1413_A net1414 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_15 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_26 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_37 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_48 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1782_A net1783 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_59 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__006__A la_data_in_mprj_bar\[23\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__379__C net15 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__395__B mprj_logic1\[100\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_050_ la_data_in_mprj_bar\[67\] vssd vssd vccd vccd net682 sky130_fd_sc_hd__clkinv_2
XFILLER_32_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2096_A mprj_logic1\[192\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input179_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input346_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2110 net2111 vssd vssd vccd vccd net2110 sky130_fd_sc_hd__buf_6
Xwire2121 net2122 vssd vssd vccd vccd net2121 sky130_fd_sc_hd__buf_6
Xwire2132 mprj_logic1\[175\] vssd vssd vccd vccd net2132 sky130_fd_sc_hd__buf_6
XFILLER_27_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2143 mprj_logic1\[165\] vssd vssd vccd vccd net2143 sky130_fd_sc_hd__buf_6
XFILLER_1_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2154 mprj_logic1\[160\] vssd vssd vccd vccd net2154 sky130_fd_sc_hd__buf_6
Xwire1420 net1421 vssd vssd vccd vccd net1420 sky130_fd_sc_hd__buf_6
Xwire2165 net2166 vssd vssd vccd vccd net2165 sky130_fd_sc_hd__buf_6
Xwire1431 net412 vssd vssd vccd vccd net1431 sky130_fd_sc_hd__buf_6
Xwire2176 mprj_logic1\[151\] vssd vssd vccd vccd net2176 sky130_fd_sc_hd__buf_6
XFILLER_5_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1442 net1443 vssd vssd vccd vccd net1442 sky130_fd_sc_hd__buf_8
Xwire2187 mprj_logic1\[146\] vssd vssd vccd vccd net2187 sky130_fd_sc_hd__buf_6
Xwire1453 net1454 vssd vssd vccd vccd net1453 sky130_fd_sc_hd__buf_6
Xwire2198 mprj_logic1\[137\] vssd vssd vccd vccd net2198 sky130_fd_sc_hd__buf_6
XFILLER_4_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__586__A net375 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1464 net1465 vssd vssd vccd vccd net1464 sky130_fd_sc_hd__buf_6
XFILLER_46_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1475 net1476 vssd vssd vccd vccd net1475 sky130_fd_sc_hd__buf_6
Xwire1486 net1487 vssd vssd vccd vccd net1486 sky130_fd_sc_hd__buf_6
Xwire1497 net397 vssd vssd vccd vccd net1497 sky130_fd_sc_hd__buf_6
XFILLER_46_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_317_ mprj_logic1\[22\] net1515 vssd vssd vccd vccd net851 sky130_fd_sc_hd__and2_1
XFILLER_50_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput13 la_data_out_mprj[108] vssd vssd vccd vccd net13 sky130_fd_sc_hd__clkbuf_4
Xinput24 la_data_out_mprj[118] vssd vssd vccd vccd net24 sky130_fd_sc_hd__buf_4
XFILLER_10_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_248_ mprj_logic1\[415\] net243 vssd vssd vccd vccd la_data_in_enable\[85\] sky130_fd_sc_hd__and2_4
XFILLER_7_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput35 la_data_out_mprj[12] vssd vssd vccd vccd net35 sky130_fd_sc_hd__clkbuf_4
Xinput46 la_data_out_mprj[22] vssd vssd vccd vccd net46 sky130_fd_sc_hd__clkbuf_4
XANTENNA_output565_A net565 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput57 la_data_out_mprj[32] vssd vssd vccd vccd net57 sky130_fd_sc_hd__clkbuf_4
Xinput68 la_data_out_mprj[42] vssd vssd vccd vccd net68 sky130_fd_sc_hd__clkbuf_4
Xinput79 la_data_out_mprj[52] vssd vssd vccd vccd net79 sky130_fd_sc_hd__clkbuf_4
X_179_ net1846 net167 vssd vssd vccd vccd la_data_in_enable\[16\] sky130_fd_sc_hd__and2_4
XANTENNA_wire1196_A net1197 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output732_A net732 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] la_data_in_enable\[77\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[77\] sky130_fd_sc_hd__nand2_8
XFILLER_38_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1530_A net373 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1628_A net105 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1997_A mprj_logic1\[281\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire983_A la_data_in_mprj_bar\[117\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput406 mprj_adr_o_core[26] vssd vssd vccd vccd net406 sky130_fd_sc_hd__buf_6
XFILLER_22_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput417 mprj_adr_o_core[7] vssd vssd vccd vccd net417 sky130_fd_sc_hd__buf_6
Xinput428 mprj_dat_o_core[16] vssd vssd vccd vccd net428 sky130_fd_sc_hd__buf_6
XFILLER_2_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput439 mprj_dat_o_core[26] vssd vssd vccd vccd net439 sky130_fd_sc_hd__buf_6
XFILLER_9_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2109_A mprj_logic1\[187\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input296_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_102_ la_data_in_mprj_bar\[119\] vssd vssd vccd vccd net612 sky130_fd_sc_hd__inv_2
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_033_ la_data_in_mprj_bar\[50\] vssd vssd vccd vccd net664 sky130_fd_sc_hd__clkinv_2
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3442 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1250 net924 vssd vssd vccd vccd net1250 sky130_fd_sc_hd__buf_6
Xwire1261 net854 vssd vssd vccd vccd net1261 sky130_fd_sc_hd__buf_6
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1272 net1273 vssd vssd vccd vccd net1272 sky130_fd_sc_hd__buf_6
XFILLER_47_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1283 net948 vssd vssd vccd vccd net1283 sky130_fd_sc_hd__buf_6
Xwire1294 net1295 vssd vssd vccd vccd net1294 sky130_fd_sc_hd__buf_8
XFILLER_38_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1209_A net1210 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output682_A net682 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__C net19 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output947_A net1284 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1480_A net1481 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1912_A net1913 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] net1316 vssd vssd vccd vccd la_data_in_mprj_bar\[103\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_26_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__392__C net47 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput203 la_iena_mprj[49] vssd vssd vccd vccd net203 sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[9\]_B la_data_in_enable\[9\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput214 la_iena_mprj[59] vssd vssd vccd vccd net214 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput225 la_iena_mprj[69] vssd vssd vccd vccd net225 sky130_fd_sc_hd__buf_4
XTAP_4702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 la_iena_mprj[79] vssd vssd vccd vccd net236 sky130_fd_sc_hd__clkbuf_4
XTAP_4713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput247 la_iena_mprj[89] vssd vssd vccd vccd net247 sky130_fd_sc_hd__clkbuf_4
Xinput258 la_iena_mprj[99] vssd vssd vccd vccd net258 sky130_fd_sc_hd__buf_4
XFILLER_5_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput269 la_oenb_mprj[108] vssd vssd vccd vccd net269 sky130_fd_sc_hd__buf_6
XFILLER_2_2721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2059_A mprj_logic1\[205\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input211_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_582_ net1532 net1984 vssd vssd vccd vccd net830 sky130_fd_sc_hd__and2_4
XFILLER_29_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input309_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__B net1981 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_016_ la_data_in_mprj_bar\[33\] vssd vssd vccd vccd net645 sky130_fd_sc_hd__inv_2
XFILLER_10_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__104__A la_data_in_mprj_bar\[121\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output528_A net1101 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1061_A net469 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1159_A net1160 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1080 net547 vssd vssd vccd vccd net1080 sky130_fd_sc_hd__buf_6
XFILLER_53_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1091 net538 vssd vssd vccd vccd net1091 sky130_fd_sc_hd__buf_6
XFILLER_1_2264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1326_A la_data_in_enable\[88\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__493__B net2076 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_740 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1695_A mprj_logic1\[71\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1738 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1862_A mprj_logic1\[335\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_length1562_A net329 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input161_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2176_A mprj_logic1\[151\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input259_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__578__B net1992 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input426_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input22_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__594__A net384 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_565_ net1549 net2016 vssd vssd vccd vccd net811 sky130_fd_sc_hd__and2_4
XFILLER_2_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_496_ net1579 net2066 net1557 vssd vssd vccd vccd net493 sky130_fd_sc_hd__and3b_4
XFILLER_35_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output478_A net478 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput507 net1120 vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__buf_8
XFILLER_29_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput518 net1110 vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__buf_8
XFILLER_9_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput529 net1100 vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__buf_8
XANTENNA_output645_A net645 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1276_A net878 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output812_A net812 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__488__B net2091 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1443_A net1444 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1708_A mprj_logic1\[65\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_max_length1310_A wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__384__A_N net294 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__398__B mprj_logic1\[103\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1805 mprj_logic1\[417\] vssd vssd vccd vccd net1805 sky130_fd_sc_hd__buf_4
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1816 mprj_logic1\[38\] vssd vssd vccd vccd net1816 sky130_fd_sc_hd__buf_6
XFILLER_28_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1827 mprj_logic1\[35\] vssd vssd vccd vccd net1827 sky130_fd_sc_hd__buf_6
XFILLER_24_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1838 mprj_logic1\[353\] vssd vssd vccd vccd net1838 sky130_fd_sc_hd__buf_6
XFILLER_41_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1849 mprj_logic1\[344\] vssd vssd vccd vccd net1849 sky130_fd_sc_hd__buf_6
XTAP_3105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_105 mprj_logic1\[232\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 mprj_logic1\[387\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 net26 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ net1719 net1383 vssd vssd vccd vccd net917 sky130_fd_sc_hd__and2_4
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_281_ net1755 net152 vssd vssd vccd vccd la_data_in_enable\[118\] sky130_fd_sc_hd__and2_4
XFILLER_14_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input376_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__589__A net379 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_617_ net1586 net1895 vssd vssd vccd vccd net742 sky130_fd_sc_hd__and2_4
XFILLER_45_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ net1558 mprj_logic1\[253\] vssd vssd vccd vccd net793 sky130_fd_sc_hd__and2_4
XTAP_2993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1024_A net773 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output595_A net595 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_479_ net272 net2115 net16 vssd vssd vccd vccd net475 sky130_fd_sc_hd__and3b_2
XFILLER_31_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output762_A net1029 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__C net28 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1393_A net421 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1658_A mprj_logic1\[88\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__499__A net310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput860 net1256 vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__buf_8
Xoutput871 net871 vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_5_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput882 net882 vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_8
XFILLER_8_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput893 net893 vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_8
XANTENNA__202__A mprj_logic1\[369\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1602 net266 vssd vssd vccd vccd net1602 sky130_fd_sc_hd__buf_6
XFILLER_8_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1613 net177 vssd vssd vccd vccd net1613 sky130_fd_sc_hd__buf_6
Xwire1624 net110 vssd vssd vccd vccd net1624 sky130_fd_sc_hd__buf_6
Xwire1635 net1636 vssd vssd vccd vccd net1635 sky130_fd_sc_hd__buf_6
Xwire1646 net1647 vssd vssd vccd vccd net1646 sky130_fd_sc_hd__buf_6
XFILLER_19_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1657 net1658 vssd vssd vccd vccd net1657 sky130_fd_sc_hd__buf_6
XFILLER_5_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1668 net1669 vssd vssd vccd vccd net1668 sky130_fd_sc_hd__buf_6
Xwire1679 mprj_logic1\[79\] vssd vssd vccd vccd net1679 sky130_fd_sc_hd__buf_6
XANTENNA_wire2041_A mprj_logic1\[216\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input124_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2139_A mprj_logic1\[170\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ net314 mprj_logic1\[107\] net58 vssd vssd vccd vccd net517 sky130_fd_sc_hd__and3b_2
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_333_ net1816 net1447 vssd vssd vccd vccd net868 sky130_fd_sc_hd__and2_4
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__591__B net1969 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_264_ net1787 net134 vssd vssd vccd vccd la_data_in_enable\[101\] sky130_fd_sc_hd__and2_2
XFILLER_10_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_195_ net1824 net185 vssd vssd vccd vccd la_data_in_enable\[32\] sky130_fd_sc_hd__and2_4
XFILLER_6_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire965 la_data_in_mprj_bar\[92\] vssd vssd vccd vccd net965 sky130_fd_sc_hd__buf_6
XFILLER_10_3875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire976 la_data_in_mprj_bar\[80\] vssd vssd vccd vccd net976 sky130_fd_sc_hd__buf_6
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[5\]
+ sky130_fd_sc_hd__nand2_4
Xwire987 la_data_in_mprj_bar\[112\] vssd vssd vccd vccd net987 sky130_fd_sc_hd__buf_6
Xwire998 net803 vssd vssd vccd vccd net998 sky130_fd_sc_hd__buf_6
XFILLER_48_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output510_A net1117 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output608_A net608 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1141_A net535 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1239_A net1240 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__485__C net1611 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1406_A net1407 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] la_data_in_enable\[22\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[22\] sky130_fd_sc_hd__nand2_4
XFILLER_32_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_16 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_27 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_38 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_49 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1775_A net1776 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1942_A mprj_logic1\[307\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__422__A_N net336 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__395__C net50 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2089_A net2090 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2100 net2101 vssd vssd vccd vccd net2100 sky130_fd_sc_hd__buf_6
Xoutput690 net690 vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_8
Xwire2111 mprj_logic1\[186\] vssd vssd vccd vccd net2111 sky130_fd_sc_hd__buf_6
XFILLER_40_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input241_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2122 mprj_logic1\[181\] vssd vssd vccd vccd net2122 sky130_fd_sc_hd__buf_6
XFILLER_8_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2133 net2134 vssd vssd vccd vccd net2133 sky130_fd_sc_hd__buf_6
XANTENNA_input339_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2144 mprj_logic1\[164\] vssd vssd vccd vccd net2144 sky130_fd_sc_hd__buf_6
XFILLER_21_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1410 net1411 vssd vssd vccd vccd net1410 sky130_fd_sc_hd__buf_6
Xwire2155 mprj_logic1\[15\] vssd vssd vccd vccd net2155 sky130_fd_sc_hd__buf_6
Xwire1421 net414 vssd vssd vccd vccd net1421 sky130_fd_sc_hd__buf_6
Xwire2166 mprj_logic1\[156\] vssd vssd vccd vccd net2166 sky130_fd_sc_hd__buf_6
XFILLER_4_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1432 net1433 vssd vssd vccd vccd net1432 sky130_fd_sc_hd__buf_8
Xwire2177 net2178 vssd vssd vccd vccd net2177 sky130_fd_sc_hd__buf_6
XFILLER_38_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1443 net1444 vssd vssd vccd vccd net1443 sky130_fd_sc_hd__buf_6
XFILLER_21_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2188 mprj_logic1\[145\] vssd vssd vccd vccd net2188 sky130_fd_sc_hd__buf_6
Xwire1454 net1455 vssd vssd vccd vccd net1454 sky130_fd_sc_hd__buf_6
Xwire2199 mprj_logic1\[12\] vssd vssd vccd vccd net2199 sky130_fd_sc_hd__buf_6
Xwire1465 net1466 vssd vssd vccd vccd net1465 sky130_fd_sc_hd__buf_6
XFILLER_1_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1476 net402 vssd vssd vccd vccd net1476 sky130_fd_sc_hd__buf_6
XANTENNA__586__B net1976 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1487 net1488 vssd vssd vccd vccd net1487 sky130_fd_sc_hd__buf_6
Xwire1498 net1499 vssd vssd vccd vccd net1498 sky130_fd_sc_hd__buf_6
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_316_ mprj_logic1\[21\] net1518 vssd vssd vccd vccd net850 sky130_fd_sc_hd__and2_2
XFILLER_10_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__107__A la_data_in_mprj_bar\[124\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput14 la_data_out_mprj[109] vssd vssd vccd vccd net14 sky130_fd_sc_hd__clkbuf_4
X_247_ mprj_logic1\[414\] net242 vssd vssd vccd vccd la_data_in_enable\[84\] sky130_fd_sc_hd__and2_4
XFILLER_32_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput25 la_data_out_mprj[119] vssd vssd vccd vccd net25 sky130_fd_sc_hd__buf_6
Xinput36 la_data_out_mprj[13] vssd vssd vccd vccd net36 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput47 la_data_out_mprj[23] vssd vssd vccd vccd net47 sky130_fd_sc_hd__clkbuf_4
Xinput58 la_data_out_mprj[33] vssd vssd vccd vccd net58 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput69 la_data_out_mprj[43] vssd vssd vccd vccd net69 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_178_ net1847 net166 vssd vssd vccd vccd la_data_in_enable\[15\] sky130_fd_sc_hd__and2_4
XFILLER_7_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output558_A net558 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1091_A net538 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__445__A_N net1541 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output725_A net725 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1356_A net1357 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__496__B net2066 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1523_A net1524 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1892_A net1893 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire976_A la_data_in_mprj_bar\[80\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_B la_data_in_enable\[32\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_40_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput407 mprj_adr_o_core[27] vssd vssd vccd vccd net407 sky130_fd_sc_hd__buf_6
XFILLER_6_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput418 mprj_adr_o_core[8] vssd vssd vccd vccd net418 sky130_fd_sc_hd__buf_6
Xinput429 mprj_dat_o_core[17] vssd vssd vccd vccd net429 sky130_fd_sc_hd__buf_6
XFILLER_22_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[99\]_B net1317 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2004_A mprj_logic1\[278\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_101_ la_data_in_mprj_bar\[118\] vssd vssd vccd vccd net611 sky130_fd_sc_hd__inv_2
XFILLER_36_1393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input191_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input289_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_032_ la_data_in_mprj_bar\[49\] vssd vssd vccd vccd net662 sky130_fd_sc_hd__inv_2
XANTENNA__468__A_N net1527 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input456_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input52_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__597__A net1607 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1240 net940 vssd vssd vccd vccd net1240 sky130_fd_sc_hd__buf_6
Xwire1251 net1252 vssd vssd vccd vccd net1251 sky130_fd_sc_hd__buf_6
XFILLER_21_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1262 net1263 vssd vssd vccd vccd net1262 sky130_fd_sc_hd__buf_6
XFILLER_40_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1273 net849 vssd vssd vccd vccd net1273 sky130_fd_sc_hd__buf_6
Xwire1284 net1285 vssd vssd vccd vccd net1284 sky130_fd_sc_hd__buf_8
XFILLER_1_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1295 net1296 vssd vssd vccd vccd net1295 sky130_fd_sc_hd__buf_8
XFILLER_47_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1104_A net525 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output842_A net842 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1473_A net1474 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B la_data_in_enable\[14\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_45_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1640_A mprj_logic1\[97\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1738_A net1739 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__300__A net1714 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1905_A net1906 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput204 la_iena_mprj[4] vssd vssd vccd vccd net204 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput215 la_iena_mprj[5] vssd vssd vccd vccd net215 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput226 la_iena_mprj[6] vssd vssd vccd vccd net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 la_iena_mprj[7] vssd vssd vccd vccd net237 sky130_fd_sc_hd__clkbuf_4
XTAP_4714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput248 la_iena_mprj[8] vssd vssd vccd vccd net248 sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput259 la_iena_mprj[9] vssd vssd vccd vccd net259 sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__210__A mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_581_ net1533 net1986 vssd vssd vccd vccd net829 sky130_fd_sc_hd__and2_4
XFILLER_44_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input204_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2121_A net2122 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_015_ la_data_in_mprj_bar\[32\] vssd vssd vccd vccd net644 sky130_fd_sc_hd__clkinv_4
XFILLER_10_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__120__A mprj_dat_i_core_bar\[6\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1070 net586 vssd vssd vccd vccd net1070 sky130_fd_sc_hd__buf_6
Xwire1081 net545 vssd vssd vccd vccd net1081 sky130_fd_sc_hd__buf_6
XFILLER_47_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1092 net537 vssd vssd vccd vccd net1092 sky130_fd_sc_hd__buf_6
XFILLER_53_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1221_A net1222 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output792_A net1009 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1319_A la_data_in_enable\[95\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__493__C net1573 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3586 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1688_A net1689 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1855_A mprj_logic1\[341\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__205__A net1821 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input154_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2071_A net2072 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2169_A net2170 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input321_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input419_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__594__B net1963 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_564_ net1550 net2017 vssd vssd vccd vccd net810 sky130_fd_sc_hd__and2_4
XTAP_3898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_495_ net1580 net2069 net1560 vssd vssd vccd vccd net492 sky130_fd_sc_hd__and3b_4
XFILLER_35_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2874 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput508 net1119 vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__buf_8
XFILLER_5_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput519 net1109 vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__buf_8
XFILLER_49_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output540_A net1089 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output638_A net638 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1171_A net1172 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_ack_gate mprj_ack_i_user net1310 vssd vssd vccd vccd mprj_ack_i_core_bar
+ sky130_fd_sc_hd__nand2_1
XANTENNA_wire1269_A net1270 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__488__C net1608 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output805_A net805 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1436_A net411 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] la_data_in_enable\[52\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[52\] sky130_fd_sc_hd__nand2_4
XFILLER_48_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3784 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1972_A mprj_logic1\[294\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__025__A la_data_in_mprj_bar\[42\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[29\]_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1806 mprj_logic1\[416\] vssd vssd vccd vccd net1806 sky130_fd_sc_hd__buf_4
XFILLER_41_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input7_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__398__C net53 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1817 mprj_logic1\[37\] vssd vssd vccd vccd net1817 sky130_fd_sc_hd__buf_6
XFILLER_24_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1828 mprj_logic1\[359\] vssd vssd vccd vccd net1828 sky130_fd_sc_hd__buf_6
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1839 mprj_logic1\[352\] vssd vssd vccd vccd net1839 sky130_fd_sc_hd__buf_6
XFILLER_41_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_106 mprj_logic1\[252\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_128 mprj_logic1\[388\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_139 mprj_logic1\[396\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_280_ net1757 net151 vssd vssd vccd vccd la_data_in_enable\[117\] sky130_fd_sc_hd__and2_4
XFILLER_30_4140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input271_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input369_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__589__B net1972 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ net1587 net1898 vssd vssd vccd vccd net740 sky130_fd_sc_hd__and2_4
XTAP_3673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_547_ net333 mprj_logic1\[252\] vssd vssd vccd vccd net792 sky130_fd_sc_hd__and2_2
XFILLER_35_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_478_ net270 net2117 net14 vssd vssd vccd vccd net473 sky130_fd_sc_hd__and3b_4
XANTENNA_output490_A net490 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output588_A net1068 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output755_A net1035 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2442 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output922_A net1198 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__499__B net2060 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1720_A net1721 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput850 net1268 vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_25_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput861 net861 vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__buf_8
XFILLER_47_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput872 net872 vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_5_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput883 net883 vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_8
XFILLER_5_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput894 net894 vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_8
XFILLER_43_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1603 net265 vssd vssd vccd vccd net1603 sky130_fd_sc_hd__buf_6
XFILLER_3_4071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1614 net176 vssd vssd vccd vccd net1614 sky130_fd_sc_hd__buf_6
Xwire1625 net108 vssd vssd vccd vccd net1625 sky130_fd_sc_hd__buf_6
XFILLER_8_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1636 mprj_logic1\[99\] vssd vssd vccd vccd net1636 sky130_fd_sc_hd__buf_6
Xwire1647 mprj_logic1\[93\] vssd vssd vccd vccd net1647 sky130_fd_sc_hd__buf_6
XFILLER_41_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1658 mprj_logic1\[88\] vssd vssd vccd vccd net1658 sky130_fd_sc_hd__buf_6
Xwire1669 mprj_logic1\[83\] vssd vssd vccd vccd net1669 sky130_fd_sc_hd__buf_6
XFILLER_19_4046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2034_A mprj_logic1\[221\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_401_ net1570 mprj_logic1\[106\] net57 vssd vssd vccd vccd net516 sky130_fd_sc_hd__and3b_2
XFILLER_15_3209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_332_ net1817 net1452 vssd vssd vccd vccd net867 sky130_fd_sc_hd__and2_4
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2201_A net2202 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_263_ net1789 net133 vssd vssd vccd vccd la_data_in_enable\[100\] sky130_fd_sc_hd__and2_4
XFILLER_6_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input82_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_194_ net1825 net184 vssd vssd vccd vccd la_data_in_enable\[31\] sky130_fd_sc_hd__and2_4
XFILLER_10_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire966 la_data_in_mprj_bar\[91\] vssd vssd vccd vccd net966 sky130_fd_sc_hd__buf_6
XFILLER_6_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire977 la_data_in_mprj_bar\[79\] vssd vssd vccd vccd net977 sky130_fd_sc_hd__buf_6
XFILLER_48_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire988 la_data_in_mprj_bar\[111\] vssd vssd vccd vccd net988 sky130_fd_sc_hd__buf_6
Xwire999 net801 vssd vssd vccd vccd net999 sky130_fd_sc_hd__buf_6
XFILLER_6_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output503_A net1124 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__374__A_N net343 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1301_A net1302 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output872_A net872 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_17 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[28\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_33_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_28 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] la_data_in_enable\[15\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[15\] sky130_fd_sc_hd__nand2_4
XANTENNA_39 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1670_A net1671 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1768_A mprj_logic1\[442\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__303__A net1654 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1935_A net1936 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] la_data_in_enable\[126\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[126\] sky130_fd_sc_hd__nand2_2
XFILLER_0_4244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__213__A mprj_logic1\[380\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput680 net680 vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_8
Xwire2101 mprj_logic1\[190\] vssd vssd vccd vccd net2101 sky130_fd_sc_hd__buf_6
Xwire2112 net2113 vssd vssd vccd vccd net2112 sky130_fd_sc_hd__buf_6
Xoutput691 net691 vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_8
XFILLER_43_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2123 mprj_logic1\[180\] vssd vssd vccd vccd net2123 sky130_fd_sc_hd__buf_6
XFILLER_5_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2134 mprj_logic1\[174\] vssd vssd vccd vccd net2134 sky130_fd_sc_hd__buf_6
XFILLER_47_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1400 net419 vssd vssd vccd vccd net1400 sky130_fd_sc_hd__buf_6
Xwire2145 mprj_logic1\[163\] vssd vssd vccd vccd net2145 sky130_fd_sc_hd__buf_6
Xwire1411 net416 vssd vssd vccd vccd net1411 sky130_fd_sc_hd__buf_6
Xwire2156 net2157 vssd vssd vccd vccd net2156 sky130_fd_sc_hd__buf_6
Xwire1422 net1423 vssd vssd vccd vccd net1422 sky130_fd_sc_hd__buf_6
Xwire2167 net2168 vssd vssd vccd vccd net2167 sky130_fd_sc_hd__buf_6
XFILLER_21_3268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input234_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1433 net1434 vssd vssd vccd vccd net1433 sky130_fd_sc_hd__buf_6
XFILLER_19_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2178 mprj_logic1\[150\] vssd vssd vccd vccd net2178 sky130_fd_sc_hd__buf_6
XFILLER_4_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1444 net1445 vssd vssd vccd vccd net1444 sky130_fd_sc_hd__buf_6
XFILLER_38_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2189 net2190 vssd vssd vccd vccd net2189 sky130_fd_sc_hd__buf_6
Xwire1455 net1456 vssd vssd vccd vccd net1455 sky130_fd_sc_hd__buf_6
Xwire1466 net405 vssd vssd vccd vccd net1466 sky130_fd_sc_hd__buf_6
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1477 net1478 vssd vssd vccd vccd net1477 sky130_fd_sc_hd__buf_6
XFILLER_19_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__397__A_N net308 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1488 net1489 vssd vssd vccd vccd net1488 sky130_fd_sc_hd__buf_6
XFILLER_41_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1499 net1500 vssd vssd vccd vccd net1499 sky130_fd_sc_hd__buf_6
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input401_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_315_ mprj_logic1\[20\] net1520 vssd vssd vccd vccd net849 sky130_fd_sc_hd__and2_2
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_246_ mprj_logic1\[413\] net241 vssd vssd vccd vccd la_data_in_enable\[83\] sky130_fd_sc_hd__and2_4
Xinput15 la_data_out_mprj[10] vssd vssd vccd vccd net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput26 la_data_out_mprj[11] vssd vssd vccd vccd net26 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput37 la_data_out_mprj[14] vssd vssd vccd vccd net37 sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput48 la_data_out_mprj[24] vssd vssd vccd vccd net48 sky130_fd_sc_hd__clkbuf_4
Xinput59 la_data_out_mprj[34] vssd vssd vccd vccd net59 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_177_ net1849 net165 vssd vssd vccd vccd la_data_in_enable\[14\] sky130_fd_sc_hd__and2_4
XFILLER_13_1372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1084_A net543 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1251_A net1252 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1349_A net450 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__496__C net1557 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1516_A net1517 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1885_A mprj_logic1\[326\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire969_A la_data_in_mprj_bar\[88\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__033__A la_data_in_mprj_bar\[50\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput408 mprj_adr_o_core[28] vssd vssd vccd vccd net408 sky130_fd_sc_hd__buf_6
XFILLER_44_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vssd vccd vccd net419 sky130_fd_sc_hd__buf_6
XFILLER_6_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__208__A net1818 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_100_ net983 vssd vssd vccd vccd net610 sky130_fd_sc_hd__inv_2
XFILLER_51_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_031_ la_data_in_mprj_bar\[48\] vssd vssd vccd vccd net661 sky130_fd_sc_hd__inv_2
XFILLER_10_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input184_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2199_A mprj_logic1\[12\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input351_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input449_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input45_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__597__B net1953 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1230 net1231 vssd vssd vccd vccd net1230 sky130_fd_sc_hd__buf_6
XFILLER_1_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1241 net1242 vssd vssd vccd vccd net1241 sky130_fd_sc_hd__buf_6
XFILLER_40_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1252 net913 vssd vssd vccd vccd net1252 sky130_fd_sc_hd__buf_6
XFILLER_21_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1263 net853 vssd vssd vccd vccd net1263 sky130_fd_sc_hd__buf_6
XFILLER_19_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1274 net1275 vssd vssd vccd vccd net1274 sky130_fd_sc_hd__buf_6
Xwire1285 net1286 vssd vssd vccd vccd net1285 sky130_fd_sc_hd__buf_8
Xwire1296 net1297 vssd vssd vccd vccd net1296 sky130_fd_sc_hd__buf_6
XFILLER_1_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__118__A mprj_dat_i_core_bar\[4\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__A_N net325 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output570_A net570 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_229_ mprj_logic1\[396\] net222 vssd vssd vccd vccd la_data_in_enable\[66\] sky130_fd_sc_hd__and2_2
XANTENNA_wire1299_A net1300 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output835_A net1045 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1466_A net405 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] la_data_in_enable\[82\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[82\] sky130_fd_sc_hd__nand2_8
XFILLER_44_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__B net1341 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3814 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput205 la_iena_mprj[50] vssd vssd vccd vccd net205 sky130_fd_sc_hd__clkbuf_4
Xinput216 la_iena_mprj[60] vssd vssd vccd vccd net216 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput227 la_iena_mprj[70] vssd vssd vccd vccd net227 sky130_fd_sc_hd__buf_4
XTAP_4704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput238 la_iena_mprj[80] vssd vssd vccd vccd net238 sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 la_iena_mprj[90] vssd vssd vccd vccd net249 sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__210__B net201 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_580_ net1534 net1988 vssd vssd vccd vccd net828 sky130_fd_sc_hd__and2_4
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__435__A_N net1551 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input399_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_786 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_014_ la_data_in_mprj_bar\[31\] vssd vssd vccd vccd net643 sky130_fd_sc_hd__clkinv_4
XFILLER_29_2805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1060 net470 vssd vssd vccd vccd net1060 sky130_fd_sc_hd__buf_6
Xwire1071 net585 vssd vssd vccd vccd net1071 sky130_fd_sc_hd__buf_6
Xwire1082 net1083 vssd vssd vccd vccd net1082 sky130_fd_sc_hd__buf_6
XFILLER_35_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1093 net1094 vssd vssd vccd vccd net1093 sky130_fd_sc_hd__buf_6
XFILLER_1_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1047_A net813 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1214_A net1215 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output785_A net1015 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output952_A net952 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[10\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_12_3598 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1750_A mprj_logic1\[451\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__458__A_N net375 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__205__B net196 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2064_A net2065 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input147_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input314_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_563_ net1551 net2018 vssd vssd vccd vccd net809 sky130_fd_sc_hd__and2_4
XTAP_3888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_494_ net1581 net2073 net1566 vssd vssd vccd vccd net491 sky130_fd_sc_hd__and3b_4
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2886 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput509 net1118 vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__buf_8
XFILLER_29_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output533_A net1096 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__131__A mprj_dat_i_core_bar\[17\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1164_A net1165 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1331_A la_data_in_enable\[83\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1429_A net1430 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] la_data_in_enable\[45\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[45\] sky130_fd_sc_hd__nand2_2
XFILLER_53_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1798_A mprj_logic1\[425\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__306__A net2200 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1965_A net1966 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] la_data_in_enable\[7\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[7\] sky130_fd_sc_hd__nand2_2
XFILLER_9_3986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1807 mprj_logic1\[412\] vssd vssd vccd vccd net1807 sky130_fd_sc_hd__buf_6
XFILLER_41_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1818 mprj_logic1\[375\] vssd vssd vccd vccd net1818 sky130_fd_sc_hd__buf_4
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1829 mprj_logic1\[358\] vssd vssd vccd vccd net1829 sky130_fd_sc_hd__buf_6
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 mprj_logic1\[252\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_129 mprj_logic1\[388\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__216__A mprj_logic1\[383\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2181_A mprj_logic1\[149\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input264_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2598 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ net1588 net1902 vssd vssd vccd vccd net739 sky130_fd_sc_hd__and2_4
XTAP_3663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ net331 net2023 vssd vssd vccd vccd net790 sky130_fd_sc_hd__and2_2
XFILLER_45_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_477_ net269 net2119 net13 vssd vssd vccd vccd net472 sky130_fd_sc_hd__and3b_4
XFILLER_50_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output483_A net483 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__126__A mprj_dat_i_core_bar\[12\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output650_A net650 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output748_A net748 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1281_A net1282 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1379_A net1380 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output915_A net1220 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1713_A mprj_logic1\[60\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire999_A net801 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__036__A la_data_in_mprj_bar\[53\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput840 net840 vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__buf_8
XFILLER_5_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput851 net1266 vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_43_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput862 net1254 vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_8_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput873 net873 vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__buf_8
Xoutput884 net884 vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_8
XFILLER_21_3406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput895 net895 vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_8
XFILLER_43_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1604 net264 vssd vssd vccd vccd net1604 sky130_fd_sc_hd__buf_6
XFILLER_28_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1615 net175 vssd vssd vccd vccd net1615 sky130_fd_sc_hd__buf_6
XFILLER_3_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1626 net107 vssd vssd vccd vccd net1626 sky130_fd_sc_hd__buf_6
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1637 net1638 vssd vssd vccd vccd net1637 sky130_fd_sc_hd__buf_6
XFILLER_24_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1648 net1649 vssd vssd vccd vccd net1648 sky130_fd_sc_hd__buf_6
Xwire1659 net1660 vssd vssd vccd vccd net1659 sky130_fd_sc_hd__buf_6
XFILLER_19_4036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ net312 mprj_logic1\[105\] net56 vssd vssd vccd vccd net515 sky130_fd_sc_hd__and3b_2
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2027_A mprj_logic1\[230\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ net1823 net1457 vssd vssd vccd vccd net866 sky130_fd_sc_hd__and2_4
XFILLER_19_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_262_ net1791 net258 vssd vssd vccd vccd la_data_in_enable\[99\] sky130_fd_sc_hd__and2_1
XFILLER_52_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input381_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_193_ net1826 net183 vssd vssd vccd vccd la_data_in_enable\[30\] sky130_fd_sc_hd__and2_4
XFILLER_6_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire967 la_data_in_mprj_bar\[90\] vssd vssd vccd vccd net967 sky130_fd_sc_hd__buf_6
XANTENNA_input75_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire978 la_data_in_mprj_bar\[78\] vssd vssd vccd vccd net978 sky130_fd_sc_hd__buf_6
XFILLER_6_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire989 la_data_in_mprj_bar\[110\] vssd vssd vccd vccd net989 sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1127_A net499 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_529_ net1570 mprj_logic1\[234\] vssd vssd vccd vccd net772 sky130_fd_sc_hd__and2_4
XTAP_2792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_18 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_29 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output865_A net865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1496_A net1497 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1663_A net1664 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__303__B net456 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1830_A mprj_logic1\[357\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1928_A net1929 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] la_data_in_enable\[119\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[119\] sky130_fd_sc_hd__nand2_4
XFILLER_0_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__213__B net205 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput670 net670 vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_8
XFILLER_27_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput681 net681 vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_8
XFILLER_5_4178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2102 net2103 vssd vssd vccd vccd net2102 sky130_fd_sc_hd__buf_6
Xoutput692 net692 vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_8
XFILLER_21_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2113 net2114 vssd vssd vccd vccd net2113 sky130_fd_sc_hd__buf_6
Xwire2124 net2125 vssd vssd vccd vccd net2124 sky130_fd_sc_hd__buf_6
XFILLER_25_3394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2135 mprj_logic1\[173\] vssd vssd vccd vccd net2135 sky130_fd_sc_hd__buf_6
XFILLER_8_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1401 net1402 vssd vssd vccd vccd net1401 sky130_fd_sc_hd__buf_6
Xwire2146 net2147 vssd vssd vccd vccd net2146 sky130_fd_sc_hd__buf_6
XFILLER_5_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1412 net1413 vssd vssd vccd vccd net1412 sky130_fd_sc_hd__buf_6
Xwire2157 net2158 vssd vssd vccd vccd net2157 sky130_fd_sc_hd__buf_6
XFILLER_28_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1423 net1424 vssd vssd vccd vccd net1423 sky130_fd_sc_hd__buf_6
Xwire2168 mprj_logic1\[155\] vssd vssd vccd vccd net2168 sky130_fd_sc_hd__buf_6
XFILLER_43_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1434 net1435 vssd vssd vccd vccd net1434 sky130_fd_sc_hd__buf_6
Xwire2179 mprj_logic1\[14\] vssd vssd vccd vccd net2179 sky130_fd_sc_hd__buf_6
Xwire1445 net1446 vssd vssd vccd vccd net1445 sky130_fd_sc_hd__buf_6
XFILLER_4_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1456 net407 vssd vssd vccd vccd net1456 sky130_fd_sc_hd__buf_6
XFILLER_38_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1467 net1468 vssd vssd vccd vccd net1467 sky130_fd_sc_hd__buf_8
XANTENNA_input227_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1478 net1479 vssd vssd vccd vccd net1478 sky130_fd_sc_hd__buf_6
Xwire1489 net399 vssd vssd vccd vccd net1489 sky130_fd_sc_hd__buf_6
XFILLER_28_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ mprj_logic1\[19\] net1398 vssd vssd vccd vccd net879 sky130_fd_sc_hd__and2_4
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_245_ net1807 net240 vssd vssd vccd vccd la_data_in_enable\[82\] sky130_fd_sc_hd__and2_4
XFILLER_32_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput16 la_data_out_mprj[110] vssd vssd vccd vccd net16 sky130_fd_sc_hd__clkbuf_4
Xinput27 la_data_out_mprj[120] vssd vssd vccd vccd net27 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput38 la_data_out_mprj[15] vssd vssd vccd vccd net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput49 la_data_out_mprj[25] vssd vssd vccd vccd net49 sky130_fd_sc_hd__clkbuf_4
X_176_ net1850 net164 vssd vssd vccd vccd la_data_in_enable\[13\] sky130_fd_sc_hd__and2_2
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1077_A net578 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1244_A net1245 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1990 net1991 vssd vssd vccd vccd net1990 sky130_fd_sc_hd__buf_6
XFILLER_18_450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1411_A net416 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__491__A_N net1584 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1509_A net1510 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1780_A net1781 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1878_A mprj_logic1\[328\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_6_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput409 mprj_adr_o_core[29] vssd vssd vccd vccd net409 sky130_fd_sc_hd__buf_6
XFILLER_25_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__208__B net199 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_030_ la_data_in_mprj_bar\[47\] vssd vssd vccd vccd net660 sky130_fd_sc_hd__inv_2
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__224__A mprj_logic1\[391\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input177_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2094_A net2095 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input344_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input38_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1220 net1221 vssd vssd vccd vccd net1220 sky130_fd_sc_hd__buf_6
XFILLER_1_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1231 net943 vssd vssd vccd vccd net1231 sky130_fd_sc_hd__buf_6
Xwire1242 net1243 vssd vssd vccd vccd net1242 sky130_fd_sc_hd__buf_6
XFILLER_5_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1253 net863 vssd vssd vccd vccd net1253 sky130_fd_sc_hd__buf_6
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1264 net1265 vssd vssd vccd vccd net1264 sky130_fd_sc_hd__buf_6
XFILLER_21_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1275 net879 vssd vssd vccd vccd net1275 sky130_fd_sc_hd__buf_6
Xwire1286 net1287 vssd vssd vccd vccd net1286 sky130_fd_sc_hd__buf_6
XFILLER_1_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1297 net1298 vssd vssd vccd vccd net1297 sky130_fd_sc_hd__buf_6
XFILLER_35_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_228_ mprj_logic1\[395\] net221 vssd vssd vccd vccd la_data_in_enable\[65\] sky130_fd_sc_hd__and2_2
XFILLER_7_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_159_ la_data_in_mprj_bar\[12\] vssd vssd vccd vccd net622 sky130_fd_sc_hd__inv_2
XFILLER_7_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1194_A net1195 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output730_A net1042 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output828_A net828 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1361_A net443 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1459_A net1460 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] la_data_in_enable\[75\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[75\] sky130_fd_sc_hd__nand2_4
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1626_A net107 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__309__A net2179 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1995_A mprj_logic1\[282\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__044__A la_data_in_mprj_bar\[61\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__387__A_N net297 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput206 la_iena_mprj[51] vssd vssd vccd vccd net206 sky130_fd_sc_hd__clkbuf_4
Xinput217 la_iena_mprj[61] vssd vssd vccd vccd net217 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput228 la_iena_mprj[71] vssd vssd vccd vccd net228 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput239 la_iena_mprj[81] vssd vssd vccd vccd net239 sky130_fd_sc_hd__clkbuf_4
XTAP_4716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2107_A mprj_logic1\[188\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_798 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input294_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_013_ la_data_in_mprj_bar\[30\] vssd vssd vccd vccd net642 sky130_fd_sc_hd__clkinv_4
XFILLER_29_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input461_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1050 net780 vssd vssd vccd vccd net1050 sky130_fd_sc_hd__buf_6
XFILLER_2_3981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1061 net469 vssd vssd vccd vccd net1061 sky130_fd_sc_hd__buf_6
XFILLER_40_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1072 net584 vssd vssd vccd vccd net1072 sky130_fd_sc_hd__buf_6
XFILLER_38_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1083 net544 vssd vssd vccd vccd net1083 sky130_fd_sc_hd__buf_6
Xwire1094 net536 vssd vssd vccd vccd net1094 sky130_fd_sc_hd__buf_6
XFILLER_53_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__129__A mprj_dat_i_core_bar\[15\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1207_A net920 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output778_A net1020 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output945_A net1294 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1576_A net1577 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__311__B net1409 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1910_A mprj_logic1\[318\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] la_data_in_enable\[101\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[101\] sky130_fd_sc_hd__nand2_2
XFILLER_53_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__502__A net343 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2057_A mprj_logic1\[206\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__402__A_N net314 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_562_ net1552 net2019 vssd vssd vccd vccd net808 sky130_fd_sc_hd__and2_4
XTAP_3878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input307_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_493_ net1582 net2076 net1573 vssd vssd vccd vccd net490 sky130_fd_sc_hd__and3b_4
XFILLER_44_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2898 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output526_A net1103 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1157_A net934 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1324_A la_data_in_enable\[90\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output895_A net895 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] la_data_in_enable\[38\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[38\] sky130_fd_sc_hd__nand2_2
XFILLER_53_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1693_A mprj_logic1\[72\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__306__B net1485 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1860_A mprj_logic1\[337\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1958_A mprj_logic1\[300\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__322__A mprj_logic1\[27\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__425__A_N net339 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1808 mprj_logic1\[411\] vssd vssd vccd vccd net1808 sky130_fd_sc_hd__buf_6
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1819 mprj_logic1\[374\] vssd vssd vccd vccd net1819 sky130_fd_sc_hd__buf_4
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_108 mprj_logic1\[252\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_119 mprj_logic1\[377\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__216__B net208 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_728 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_B net1332 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__232__A net1813 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input257_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2174_A mprj_logic1\[152\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input424_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_614_ net1589 net1905 vssd vssd vccd vccd net738 sky130_fd_sc_hd__and2_4
XTAP_4398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_545_ net1559 mprj_logic1\[250\] vssd vssd vccd vccd net789 sky130_fd_sc_hd__and2_4
XFILLER_35_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_476_ net1600 net2121 net12 vssd vssd vccd vccd net471 sky130_fd_sc_hd__and3b_4
XFILLER_53_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output476_A net1055 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B la_data_in_enable\[71\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__448__A_N net1538 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output643_A net643 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__142__A mprj_dat_i_core_bar\[28\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1274_A net1275 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output810_A net810 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1441_A net410 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1539_A net363 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_4251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1706_A net1707 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput830 net830 vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__buf_8
XANTENNA__052__A la_data_in_mprj_bar\[69\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput841 net841 vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__buf_8
XFILLER_25_3521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput852 net1264 vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput863 net1253 vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__buf_8
Xoutput874 net874 vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_28_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput885 net885 vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_8
Xoutput896 net896 vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_8
XFILLER_43_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1605 net263 vssd vssd vccd vccd net1605 sky130_fd_sc_hd__buf_6
XFILLER_8_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1616 net118 vssd vssd vccd vccd net1616 sky130_fd_sc_hd__buf_6
XFILLER_5_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1627 net106 vssd vssd vccd vccd net1627 sky130_fd_sc_hd__buf_6
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1638 mprj_logic1\[98\] vssd vssd vccd vccd net1638 sky130_fd_sc_hd__buf_6
XFILLER_19_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1649 mprj_logic1\[92\] vssd vssd vccd vccd net1649 sky130_fd_sc_hd__buf_6
XFILLER_6_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ net1827 net1462 vssd vssd vccd vccd net865 sky130_fd_sc_hd__and2_4
XFILLER_26_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__227__A mprj_logic1\[394\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_261_ net1793 net257 vssd vssd vccd vccd la_data_in_enable\[98\] sky130_fd_sc_hd__and2_4
XFILLER_17_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_192_ net1828 net181 vssd vssd vccd vccd la_data_in_enable\[29\] sky130_fd_sc_hd__and2_2
XFILLER_48_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_2289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire968 la_data_in_mprj_bar\[89\] vssd vssd vccd vccd net968 sky130_fd_sc_hd__buf_6
Xwire979 la_data_in_mprj_bar\[127\] vssd vssd vccd vccd net979 sky130_fd_sc_hd__buf_6
XANTENNA_input374_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input68_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_528_ net1571 mprj_logic1\[233\] vssd vssd vccd vccd net771 sky130_fd_sc_hd__and2_4
XFILLER_50_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1022_A net1023 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output593_A net593 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__137__A mprj_dat_i_core_bar\[23\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_459_ net377 net2144 net121 vssd vssd vccd vccd net580 sky130_fd_sc_hd__and3b_4
XANTENNA_19 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output760_A net1031 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output858_A net1257 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1391_A net1392 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1656_A mprj_logic1\[89\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__600__A net1604 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1823_A mprj_logic1\[36\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__047__A la_data_in_mprj_bar\[64\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[35\]_B la_data_in_enable\[35\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_49_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput660 net660 vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_8
XFILLER_40_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput671 net671 vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_8
Xoutput682 net682 vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_8
Xwire2103 net2104 vssd vssd vccd vccd net2103 sky130_fd_sc_hd__buf_6
Xoutput693 net693 vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_8
XFILLER_8_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2114 mprj_logic1\[185\] vssd vssd vccd vccd net2114 sky130_fd_sc_hd__buf_6
Xwire2125 mprj_logic1\[179\] vssd vssd vccd vccd net2125 sky130_fd_sc_hd__buf_6
XANTENNA__510__A net292 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2136 mprj_logic1\[172\] vssd vssd vccd vccd net2136 sky130_fd_sc_hd__buf_6
XFILLER_8_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1402 net1403 vssd vssd vccd vccd net1402 sky130_fd_sc_hd__buf_6
XFILLER_21_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2147 net2148 vssd vssd vccd vccd net2147 sky130_fd_sc_hd__buf_6
Xwire1413 net1414 vssd vssd vccd vccd net1413 sky130_fd_sc_hd__buf_6
Xwire2158 mprj_logic1\[159\] vssd vssd vccd vccd net2158 sky130_fd_sc_hd__buf_6
XFILLER_25_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1424 net1425 vssd vssd vccd vccd net1424 sky130_fd_sc_hd__buf_6
Xwire2169 net2170 vssd vssd vccd vccd net2169 sky130_fd_sc_hd__buf_6
Xwire1435 net1436 vssd vssd vccd vccd net1435 sky130_fd_sc_hd__buf_6
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1446 net409 vssd vssd vccd vccd net1446 sky130_fd_sc_hd__buf_6
Xwire1457 net1458 vssd vssd vccd vccd net1457 sky130_fd_sc_hd__buf_8
Xwire1468 net1469 vssd vssd vccd vccd net1468 sky130_fd_sc_hd__buf_6
Xwire1479 net1480 vssd vssd vccd vccd net1479 sky130_fd_sc_hd__buf_6
XFILLER_38_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input122_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2137_A net2138 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_313_ mprj_logic1\[18\] net1401 vssd vssd vccd vccd net878 sky130_fd_sc_hd__and2_2
XFILLER_35_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_244_ net1808 net239 vssd vssd vccd vccd la_data_in_enable\[81\] sky130_fd_sc_hd__and2_4
XFILLER_10_340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput17 la_data_out_mprj[111] vssd vssd vccd vccd net17 sky130_fd_sc_hd__clkbuf_4
Xinput28 la_data_out_mprj[121] vssd vssd vccd vccd net28 sky130_fd_sc_hd__buf_4
XFILLER_10_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput39 la_data_out_mprj[16] vssd vssd vccd vccd net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_175_ net1852 net163 vssd vssd vccd vccd la_data_in_enable\[12\] sky130_fd_sc_hd__and2_1
XFILLER_6_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[3\]
+ sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[110\]_B la_data_in_enable\[110\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_6_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output606_A net606 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1980 mprj_logic1\[289\] vssd vssd vccd vccd net1980 sky130_fd_sc_hd__buf_6
Xwire1991 mprj_logic1\[284\] vssd vssd vccd vccd net1991 sky130_fd_sc_hd__buf_6
XFILLER_4_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1404_A net418 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] la_data_in_enable\[20\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[20\] sky130_fd_sc_hd__nand2_1
XFILLER_53_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1773_A net1774 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[17\]_B la_data_in_enable\[17\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__314__B net1398 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1940_A mprj_logic1\[308\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__330__A net1827 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__505__A net376 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2087_A mprj_logic1\[195\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__A mprj_logic1\[407\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput490 net490 vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__buf_8
XFILLER_43_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input337_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1210 net919 vssd vssd vccd vccd net1210 sky130_fd_sc_hd__buf_6
XFILLER_43_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1221 net1222 vssd vssd vccd vccd net1221 sky130_fd_sc_hd__buf_6
Xwire1232 net1233 vssd vssd vccd vccd net1232 sky130_fd_sc_hd__buf_6
XFILLER_38_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1243 net939 vssd vssd vccd vccd net1243 sky130_fd_sc_hd__buf_6
Xwire1254 net1255 vssd vssd vccd vccd net1254 sky130_fd_sc_hd__buf_6
XFILLER_19_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1265 net852 vssd vssd vccd vccd net1265 sky130_fd_sc_hd__buf_6
XFILLER_5_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1276 net878 vssd vssd vccd vccd net1276 sky130_fd_sc_hd__buf_6
XFILLER_38_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1287 net1288 vssd vssd vccd vccd net1287 sky130_fd_sc_hd__buf_6
Xwire1298 net945 vssd vssd vccd vccd net1298 sky130_fd_sc_hd__buf_6
XFILLER_34_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_227_ mprj_logic1\[394\] net220 vssd vssd vccd vccd la_data_in_enable\[64\] sky130_fd_sc_hd__and2_2
XFILLER_45_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_158_ la_data_in_mprj_bar\[11\] vssd vssd vccd vccd net613 sky130_fd_sc_hd__inv_2
XFILLER_13_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output556_A net556 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_089_ la_data_in_mprj_bar\[106\] vssd vssd vccd vccd net598 sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1187_A net1188 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output723_A net723 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1354_A net1355 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] la_data_in_enable\[68\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[68\] sky130_fd_sc_hd__nand2_4
XFILLER_22_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1521_A net389 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1619_A net115 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__309__B net1417 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1890_A net1891 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1988_A net1989 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire974_A la_data_in_mprj_bar\[83\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3859 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__060__A la_data_in_mprj_bar\[77\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput207 la_iena_mprj[52] vssd vssd vccd vccd net207 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput218 la_iena_mprj[62] vssd vssd vccd vccd net218 sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vssd vccd vccd net229 sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_958 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2002_A mprj_logic1\[279\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__235__A mprj_logic1\[402\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input287_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_012_ la_data_in_mprj_bar\[29\] vssd vssd vccd vccd net640 sky130_fd_sc_hd__clkinv_4
XFILLER_4_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input454_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input50_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__481__A_N net1594 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__401__C net57 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1040 net750 vssd vssd vccd vccd net1040 sky130_fd_sc_hd__buf_6
Xwire1051 net769 vssd vssd vccd vccd net1051 sky130_fd_sc_hd__buf_6
Xwire1062 net468 vssd vssd vccd vccd net1062 sky130_fd_sc_hd__buf_6
Xwire1073 net583 vssd vssd vccd vccd net1073 sky130_fd_sc_hd__buf_6
XFILLER_40_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1084 net543 vssd vssd vccd vccd net1084 sky130_fd_sc_hd__buf_6
XFILLER_35_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1095 net534 vssd vssd vccd vccd net1095 sky130_fd_sc_hd__buf_6
XFILLER_18_3913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1102_A net527 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__145__A mprj_dat_i_core_bar\[31\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output840_A net840 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output938_A net1244 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1471_A net404 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1736_A net1737 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1903_A net1904 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__055__A la_data_in_mprj_bar\[72\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__502__B net2055 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_561_ net1553 net2020 vssd vssd vccd vccd net807 sky130_fd_sc_hd__and2_4
XTAP_3868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input202_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_492_ net1583 net2079 net30 vssd vssd vccd vccd net489 sky130_fd_sc_hd__and3b_4
XFILLER_44_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input98_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__B mprj_logic1\[117\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output519_A net1109 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1052_A net758 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__377__A_N net376 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3754 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output790_A net1011 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1686_A net1687 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__603__A net1601 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1853_A mprj_logic1\[342\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__322__B net1498 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1809 mprj_logic1\[40\] vssd vssd vccd vccd net1809 sky130_fd_sc_hd__buf_6
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_109 mprj_logic1\[252\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__513__A net295 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__232__B net225 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input152_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2167_A net2168 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input417_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_613_ net1590 net1908 vssd vssd vccd vccd net737 sky130_fd_sc_hd__and2_4
XTAP_4388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_544_ net1561 mprj_logic1\[249\] vssd vssd vccd vccd net788 sky130_fd_sc_hd__and2_4
XTAP_3698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_475_ net1601 net2123 net11 vssd vssd vccd vccd net470 sky130_fd_sc_hd__and3b_4
XFILLER_15_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__407__B mprj_logic1\[112\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output469_A net1061 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output636_A net636 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output803_A net997 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1434_A net1435 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput390 mprj_adr_o_core[11] vssd vssd vccd vccd net390 sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] la_data_in_enable\[50\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[50\] sky130_fd_sc_hd__nand2_4
XFILLER_53_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__317__B net1515 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1970_A mprj_logic1\[296\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__A net1816 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput820 net820 vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__buf_8
XFILLER_47_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput831 net831 vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__buf_8
XFILLER_9_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput842 net842 vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__buf_8
XFILLER_8_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput853 net1262 vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__buf_8
XFILLER_25_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput864 net864 vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__buf_8
XFILLER_43_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput875 net875 vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__buf_8
Xoutput886 net886 vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_8
Xoutput897 net897 vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_8
XFILLER_25_3577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1606 net262 vssd vssd vccd vccd net1606 sky130_fd_sc_hd__buf_6
XANTENNA_input5_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1617 net117 vssd vssd vccd vccd net1617 sky130_fd_sc_hd__buf_6
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1628 net105 vssd vssd vccd vccd net1628 sky130_fd_sc_hd__buf_6
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1639 net1640 vssd vssd vccd vccd net1639 sky130_fd_sc_hd__buf_6
XFILLER_3_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__508__A net282 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__227__B net220 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_260_ net1795 net256 vssd vssd vccd vccd la_data_in_enable\[97\] sky130_fd_sc_hd__and2_4
XFILLER_23_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_191_ net1829 net180 vssd vssd vccd vccd la_data_in_enable\[28\] sky130_fd_sc_hd__and2_2
XFILLER_32_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire969 la_data_in_mprj_bar\[88\] vssd vssd vccd vccd net969 sky130_fd_sc_hd__buf_6
XFILLER_10_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__243__A mprj_logic1\[410\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input367_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_irq_gates\[2\] user_irq_core[2] user_irq_enable\[2\] vssd vssd vccd vccd user_irq_bar\[2\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_43_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_527_ net1572 mprj_logic1\[232\] vssd vssd vccd vccd net770 sky130_fd_sc_hd__and2_2
XFILLER_15_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_458_ net375 net2145 net119 vssd vssd vccd vccd net578 sky130_fd_sc_hd__and3b_4
XANTENNA__415__A_N net328 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output586_A net1070 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_389_ net300 net1645 net44 vssd vssd vccd vccd net503 sky130_fd_sc_hd__and3b_4
XFILLER_31_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output753_A net1037 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output920_A net1205 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] la_data_in_enable\[98\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[98\] sky130_fd_sc_hd__nand2_8
XFILLER_29_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1649_A mprj_logic1\[92\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__600__B net1945 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1816_A mprj_logic1\[38\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__063__A net976 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput650 net650 vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_8
Xoutput661 net661 vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_8
XFILLER_9_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput672 net672 vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_8
XFILLER_40_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput683 net683 vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_8
XFILLER_44_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2104 mprj_logic1\[189\] vssd vssd vccd vccd net2104 sky130_fd_sc_hd__buf_6
Xwire2115 net2116 vssd vssd vccd vccd net2115 sky130_fd_sc_hd__buf_6
Xoutput694 net694 vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_8
XFILLER_8_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2126 net2127 vssd vssd vccd vccd net2126 sky130_fd_sc_hd__buf_6
XANTENNA__510__B net2042 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2137 net2138 vssd vssd vccd vccd net2137 sky130_fd_sc_hd__buf_6
Xwire1403 net1404 vssd vssd vccd vccd net1403 sky130_fd_sc_hd__buf_6
Xwire2148 mprj_logic1\[162\] vssd vssd vccd vccd net2148 sky130_fd_sc_hd__buf_6
XFILLER_5_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1414 net1415 vssd vssd vccd vccd net1414 sky130_fd_sc_hd__buf_6
Xwire2159 net2160 vssd vssd vccd vccd net2159 sky130_fd_sc_hd__buf_6
Xwire1425 net1426 vssd vssd vccd vccd net1425 sky130_fd_sc_hd__buf_6
XFILLER_25_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1436 net411 vssd vssd vccd vccd net1436 sky130_fd_sc_hd__buf_6
Xwire1447 net1448 vssd vssd vccd vccd net1447 sky130_fd_sc_hd__buf_8
Xwire1458 net1459 vssd vssd vccd vccd net1458 sky130_fd_sc_hd__buf_6
Xwire1469 net1470 vssd vssd vccd vccd net1469 sky130_fd_sc_hd__buf_6
XFILLER_28_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2032_A mprj_logic1\[223\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input115_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__438__A_N net1548 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__238__A mprj_logic1\[405\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ mprj_logic1\[17\] net1405 vssd vssd vccd vccd net877 sky130_fd_sc_hd__and2_2
XFILLER_51_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_2488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_243_ mprj_logic1\[410\] net238 vssd vssd vccd vccd la_data_in_enable\[80\] sky130_fd_sc_hd__and2_2
XFILLER_32_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput18 la_data_out_mprj[112] vssd vssd vccd vccd net18 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input80_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput29 la_data_out_mprj[122] vssd vssd vccd vccd net29 sky130_fd_sc_hd__clkbuf_4
X_174_ net1854 net154 vssd vssd vccd vccd la_data_in_enable\[11\] sky130_fd_sc_hd__and2_2
XFILLER_6_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__404__C net60 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__420__B mprj_logic1\[125\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1690 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1970 mprj_logic1\[296\] vssd vssd vccd vccd net1970 sky130_fd_sc_hd__buf_6
XFILLER_19_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output501_A net1125 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1981 net1982 vssd vssd vccd vccd net1981 sky130_fd_sc_hd__buf_6
XFILLER_37_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1992 net1993 vssd vssd vccd vccd net1992 sky130_fd_sc_hd__buf_6
XFILLER_15_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1132_A net494 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] la_data_in_enable\[13\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[13\] sky130_fd_sc_hd__nand2_2
XFILLER_53_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[26\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_14_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1599_A net269 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1766_A mprj_logic1\[443\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__611__A net1592 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__330__B net1462 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] net1312 vssd vssd vccd vccd la_data_in_mprj_bar\[124\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__058__A la_data_in_mprj_bar\[75\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[10\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__505__B net2051 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__521__A net304 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput480 net480 vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__buf_8
Xoutput491 net491 vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__buf_8
XFILLER_40_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__B net234 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1200 net1201 vssd vssd vccd vccd net1200 sky130_fd_sc_hd__buf_6
Xwire1211 net1212 vssd vssd vccd vccd net1211 sky130_fd_sc_hd__buf_6
XFILLER_43_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1222 net915 vssd vssd vccd vccd net1222 sky130_fd_sc_hd__buf_6
Xwire1233 net1234 vssd vssd vccd vccd net1233 sky130_fd_sc_hd__buf_6
XANTENNA_input232_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1244 net1245 vssd vssd vccd vccd net1244 sky130_fd_sc_hd__buf_6
XFILLER_5_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1255 net862 vssd vssd vccd vccd net1255 sky130_fd_sc_hd__buf_6
Xwire1266 net1267 vssd vssd vccd vccd net1266 sky130_fd_sc_hd__buf_6
Xwire1277 net877 vssd vssd vccd vccd net1277 sky130_fd_sc_hd__buf_6
XFILLER_35_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1288 net947 vssd vssd vccd vccd net1288 sky130_fd_sc_hd__buf_6
Xwire1299 net1300 vssd vssd vccd vccd net1299 sky130_fd_sc_hd__buf_8
XFILLER_38_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_226_ mprj_logic1\[393\] net219 vssd vssd vccd vccd la_data_in_enable\[63\] sky130_fd_sc_hd__and2_2
XANTENNA__415__B mprj_logic1\[120\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_157_ la_data_in_mprj_bar\[10\] vssd vssd vccd vccd net602 sky130_fd_sc_hd__clkinv_2
XFILLER_6_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_088_ la_data_in_mprj_bar\[105\] vssd vssd vccd vccd net597 sky130_fd_sc_hd__clkinv_4
XFILLER_45_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output549_A net1078 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1082_A net1083 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output716_A net716 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1347_A net451 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__606__A net1597 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1883_A net1884 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__325__B net1482 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire967_A la_data_in_mprj_bar\[90\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__341__A mprj_logic1\[46\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4034 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput208 la_iena_mprj[53] vssd vssd vccd vccd net208 sky130_fd_sc_hd__clkbuf_4
Xinput219 la_iena_mprj[63] vssd vssd vccd vccd net219 sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__516__A net298 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__235__B net229 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_011_ la_data_in_mprj_bar\[28\] vssd vssd vccd vccd net639 sky130_fd_sc_hd__clkinv_4
XFILLER_46_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input182_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2197_A mprj_logic1\[138\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__251__A net1804 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input447_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1030 net761 vssd vssd vccd vccd net1030 sky130_fd_sc_hd__buf_6
XFILLER_7_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1041 net741 vssd vssd vccd vccd net1041 sky130_fd_sc_hd__buf_6
XFILLER_2_3961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1052 net758 vssd vssd vccd vccd net1052 sky130_fd_sc_hd__buf_6
XFILLER_38_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1063 net467 vssd vssd vccd vccd net1063 sky130_fd_sc_hd__buf_6
Xwire1074 net582 vssd vssd vccd vccd net1074 sky130_fd_sc_hd__buf_6
Xwire1085 net1086 vssd vssd vccd vccd net1085 sky130_fd_sc_hd__buf_6
XFILLER_1_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1096 net533 vssd vssd vccd vccd net1096 sky130_fd_sc_hd__buf_6
XFILLER_1_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output499_A net1127 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_209_ mprj_logic1\[376\] net200 vssd vssd vccd vccd la_data_in_enable\[46\] sky130_fd_sc_hd__and2_1
XFILLER_32_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1297_A net1298 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output833_A net833 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__161__A la_data_in_mprj_bar\[14\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1464_A net1465 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] net1332 vssd vssd vccd vccd la_data_in_mprj_bar\[80\]
+ sky130_fd_sc_hd__nand2_4
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1806 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1631_A net102 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1729_A net1730 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__336__A net1803 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__071__A net969 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_560_ net1554 net2021 vssd vssd vccd vccd net806 sky130_fd_sc_hd__and2_4
XTAP_3858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_491_ net1584 net2082 net29 vssd vssd vccd vccd net488 sky130_fd_sc_hd__and3b_4
XFILLER_35_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2112_A net2113 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__246__A mprj_logic1\[413\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input397_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__C net69 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1045_A net835 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3766 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1212_A net1213 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output783_A net1016 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__156__A la_data_in_mprj_bar\[9\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output950_A net1299 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1679_A mprj_logic1\[79\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__603__B net1939 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1846_A mprj_logic1\[346\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[2\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__471__A_N net1605 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__066__A net974 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__513__B net2037 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2062_A net2063 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input145_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_612_ net1591 net1911 vssd vssd vccd vccd net736 sky130_fd_sc_hd__and2_4
XTAP_4378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input312_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_543_ net1563 mprj_logic1\[248\] vssd vssd vccd vccd net787 sky130_fd_sc_hd__and2_4
XTAP_2932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_474_ net1602 net2124 net10 vssd vssd vccd vccd net469 sky130_fd_sc_hd__and3b_4
XFILLER_13_4320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__423__B mprj_logic1\[128\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output531_A net1098 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1162_A net1163 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput380 la_oenb_mprj[93] vssd vssd vccd vccd net380 sky130_fd_sc_hd__buf_8
XFILLER_42_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput391 mprj_adr_o_core[12] vssd vssd vccd vccd net391 sky130_fd_sc_hd__buf_6
XFILLER_36_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1427_A net1428 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__494__A_N net1581 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] la_data_in_enable\[43\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[43\] sky130_fd_sc_hd__nand2_2
XFILLER_18_3530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1090 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A net1589 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1963_A net1964 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__B net1447 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput810 net810 vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__buf_8
Xoutput821 net821 vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__buf_8
Xoutput832 net832 vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__buf_8
XFILLER_47_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput843 net843 vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__buf_8
XFILLER_9_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput854 net1261 vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__buf_8
Xoutput865 net865 vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] la_data_in_enable\[5\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[5\] sky130_fd_sc_hd__nand2_2
Xoutput876 net1278 vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__buf_8
XFILLER_8_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput887 net887 vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_8
XFILLER_28_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput898 net898 vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_8
XFILLER_25_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1607 net261 vssd vssd vccd vccd net1607 sky130_fd_sc_hd__buf_6
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1618 net116 vssd vssd vccd vccd net1618 sky130_fd_sc_hd__buf_6
XFILLER_3_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1629 net104 vssd vssd vccd vccd net1629 sky130_fd_sc_hd__buf_6
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__508__B net2045 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_190_ net1830 net179 vssd vssd vccd vccd la_data_in_enable\[27\] sky130_fd_sc_hd__and2_1
XFILLER_10_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__524__A net1575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__243__B net238 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input262_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__418__B mprj_logic1\[123\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_526_ net1574 mprj_logic1\[231\] vssd vssd vccd vccd net768 sky130_fd_sc_hd__and2_4
XFILLER_50_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_457_ net1529 net2146 net1616 vssd vssd vccd vccd net577 sky130_fd_sc_hd__and3b_4
XFILLER_53_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_388_ net298 net1646 net42 vssd vssd vccd vccd net501 sky130_fd_sc_hd__and3b_4
XANTENNA_output481_A net481 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output579_A net1137 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output746_A net746 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1377_A net429 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output913_A net1251 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1544_A net358 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1711_A mprj_logic1\[62\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1809_A mprj_logic1\[40\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__609__A net1594 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__328__B net1472 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire997_A net998 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__344__A mprj_logic1\[49\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_10_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput640 net640 vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_8
XFILLER_5_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput651 net651 vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_8
XFILLER_25_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput662 net662 vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_8
XFILLER_25_3353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput673 net673 vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_8
Xoutput684 net684 vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_8
Xwire2105 net2106 vssd vssd vccd vccd net2105 sky130_fd_sc_hd__buf_6
XFILLER_40_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput695 net695 vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_8
Xwire2116 mprj_logic1\[184\] vssd vssd vccd vccd net2116 sky130_fd_sc_hd__buf_6
XFILLER_47_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2127 mprj_logic1\[178\] vssd vssd vccd vccd net2127 sky130_fd_sc_hd__buf_6
Xwire2138 mprj_logic1\[171\] vssd vssd vccd vccd net2138 sky130_fd_sc_hd__buf_6
Xwire1404 net418 vssd vssd vccd vccd net1404 sky130_fd_sc_hd__buf_6
XFILLER_21_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2149 net2150 vssd vssd vccd vccd net2149 sky130_fd_sc_hd__buf_6
Xwire1415 net1416 vssd vssd vccd vccd net1415 sky130_fd_sc_hd__buf_6
Xwire1426 net413 vssd vssd vccd vccd net1426 sky130_fd_sc_hd__buf_6
XFILLER_3_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1437 net1438 vssd vssd vccd vccd net1437 sky130_fd_sc_hd__buf_8
XFILLER_47_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1448 net1449 vssd vssd vccd vccd net1448 sky130_fd_sc_hd__buf_6
Xwire1459 net1460 vssd vssd vccd vccd net1459 sky130_fd_sc_hd__buf_6
XFILLER_28_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__519__A net302 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__238__B net232 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input108_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_311_ mprj_logic1\[16\] net1409 vssd vssd vccd vccd net876 sky130_fd_sc_hd__and2_4
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_242_ mprj_logic1\[409\] net236 vssd vssd vccd vccd la_data_in_enable\[79\] sky130_fd_sc_hd__and2_2
XFILLER_52_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__254__A net1802 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput19 la_data_out_mprj[113] vssd vssd vccd vccd net19 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_173_ net1856 net143 vssd vssd vccd vccd la_data_in_enable\[10\] sky130_fd_sc_hd__and2_1
XFILLER_32_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input73_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__420__C net78 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1960 net1961 vssd vssd vccd vccd net1960 sky130_fd_sc_hd__buf_6
Xwire1971 mprj_logic1\[295\] vssd vssd vccd vccd net1971 sky130_fd_sc_hd__buf_6
XFILLER_20_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1982 net1983 vssd vssd vccd vccd net1982 sky130_fd_sc_hd__buf_6
XFILLER_4_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1993 mprj_logic1\[283\] vssd vssd vccd vccd net1993 sky130_fd_sc_hd__buf_6
XTAP_3260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1125_A net501 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_509_ net291 net2044 vssd vssd vccd vccd net750 sky130_fd_sc_hd__and2_4
XFILLER_37_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output863_A net1253 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__164__A net1869 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[19\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1494_A net1495 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1661_A net1662 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1759_A net1760 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__611__B net1915 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1926_A net1927 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] la_data_in_enable\[117\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[117\] sky130_fd_sc_hd__nand2_4
XFILLER_0_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__074__A net966 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3986 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__521__B net2029 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput470 net1060 vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__buf_8
XFILLER_44_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput481 net481 vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__buf_8
XFILLER_47_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput492 net492 vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__buf_8
XFILLER_40_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__405__A_N net317 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1201 net922 vssd vssd vccd vccd net1201 sky130_fd_sc_hd__buf_6
XFILLER_25_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1212 net1213 vssd vssd vccd vccd net1212 sky130_fd_sc_hd__buf_6
Xwire1223 net1224 vssd vssd vccd vccd net1223 sky130_fd_sc_hd__buf_6
XFILLER_43_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1234 net942 vssd vssd vccd vccd net1234 sky130_fd_sc_hd__buf_6
Xwire1245 net938 vssd vssd vccd vccd net1245 sky130_fd_sc_hd__buf_6
XFILLER_1_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1256 net860 vssd vssd vccd vccd net1256 sky130_fd_sc_hd__buf_6
XFILLER_21_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2142_A mprj_logic1\[166\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input225_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1267 net851 vssd vssd vccd vccd net1267 sky130_fd_sc_hd__buf_6
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1278 net1279 vssd vssd vccd vccd net1278 sky130_fd_sc_hd__buf_6
XFILLER_21_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1289 net1290 vssd vssd vccd vccd net1289 sky130_fd_sc_hd__buf_8
XFILLER_34_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__249__A net1806 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_225_ mprj_logic1\[392\] net218 vssd vssd vccd vccd la_data_in_enable\[62\] sky130_fd_sc_hd__and2_2
XFILLER_11_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__415__C net72 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_156_ la_data_in_mprj_bar\[9\] vssd vssd vccd vccd net718 sky130_fd_sc_hd__inv_2
XFILLER_32_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_087_ la_data_in_mprj_bar\[104\] vssd vssd vccd vccd net596 sky130_fd_sc_hd__clkinv_4
XFILLER_49_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__B mprj_logic1\[136\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1075_A net581 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output611_A net611 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output709_A net709 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1242_A net1243 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1790 mprj_logic1\[430\] vssd vssd vccd vccd net1790 sky130_fd_sc_hd__buf_6
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1507_A net1508 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__606__B net1931 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1876_A net1877 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__622__A net1581 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__341__B net1354 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__428__A_N net342 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput209 la_iena_mprj[54] vssd vssd vccd vccd net209 sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__069__A net971 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__516__B net2034 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_010_ la_data_in_mprj_bar\[27\] vssd vssd vccd vccd net638 sky130_fd_sc_hd__inv_4
XFILLER_10_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__532__A net1569 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2092_A net2093 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input175_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3278 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input342_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input36_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1020 net1021 vssd vssd vccd vccd net1020 sky130_fd_sc_hd__buf_6
XFILLER_0_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1031 net760 vssd vssd vccd vccd net1031 sky130_fd_sc_hd__buf_6
XFILLER_1_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1042 net1043 vssd vssd vccd vccd net1042 sky130_fd_sc_hd__buf_6
Xwire1053 net719 vssd vssd vccd vccd net1053 sky130_fd_sc_hd__buf_6
XFILLER_5_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1064 net466 vssd vssd vccd vccd net1064 sky130_fd_sc_hd__buf_6
XFILLER_53_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1075 net581 vssd vssd vccd vccd net1075 sky130_fd_sc_hd__buf_6
Xwire1086 net542 vssd vssd vccd vccd net1086 sky130_fd_sc_hd__buf_6
Xwire1097 net532 vssd vssd vccd vccd net1097 sky130_fd_sc_hd__buf_6
XFILLER_35_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_208_ net1818 net199 vssd vssd vccd vccd la_data_in_enable\[45\] sky130_fd_sc_hd__and2_1
XFILLER_45_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output561_A net561 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output659_A net659 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_139_ mprj_dat_i_core_bar\[25\] vssd vssd vccd vccd net898 sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1192_A net1193 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output826_A net826 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1457_A net1458 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] la_data_in_enable\[73\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[73\] sky130_fd_sc_hd__nand2_4
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1624_A net110 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__617__A net1586 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1993_A mprj_logic1\[283\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__336__B net1427 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2924 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_B net1322 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__352__A net1717 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_490_ net1585 net2085 net28 vssd vssd vccd vccd net487 sky130_fd_sc_hd__and3b_4
XANTENNA__527__A net1572 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2105_A net2106 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input292_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_B net1331 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__262__A net1791 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xmax_length1562 net329 vssd vssd vccd vccd net1562 sky130_fd_sc_hd__buf_6
XFILLER_4_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1038_A net752 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1205_A net1206 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output776_A net776 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[74\]_B la_data_in_enable\[74\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output943_A net1229 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__172__A net1857 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1741_A mprj_logic1\[455\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1839_A mprj_logic1\[352\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1058 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__347__A mprj_logic1\[52\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__082__A net961 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input138_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2055_A net2056 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_611_ net1592 net1915 vssd vssd vccd vccd net735 sky130_fd_sc_hd__and2_4
XFILLER_29_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_542_ net327 mprj_logic1\[247\] vssd vssd vccd vccd net786 sky130_fd_sc_hd__and2_2
XTAP_3678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input305_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__257__A net1799 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_473_ net1603 net2126 net9 vssd vssd vccd vccd net468 sky130_fd_sc_hd__and3b_4
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__423__C net81 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3810 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output524_A net1142 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1155_A net1156 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput370 la_oenb_mprj[84] vssd vssd vccd vccd net370 sky130_fd_sc_hd__buf_6
Xinput381 la_oenb_mprj[94] vssd vssd vccd vccd net381 sky130_fd_sc_hd__buf_6
XFILLER_7_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput392 mprj_adr_o_core[13] vssd vssd vccd vccd net392 sky130_fd_sc_hd__buf_6
XFILLER_40_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1322_A la_data_in_enable\[92\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__167__A net1863 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] la_data_in_enable\[36\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[36\] sky130_fd_sc_hd__nand2_4
XFILLER_36_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1691_A mprj_logic1\[73\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1789_A net1790 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__614__B net1905 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1956_A mprj_logic1\[301\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput800 net1000 vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__buf_8
Xoutput811 net811 vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__buf_8
XFILLER_9_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput822 net822 vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__buf_8
Xoutput833 net833 vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__buf_8
Xoutput844 net844 vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__buf_8
Xoutput855 net1260 vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_47_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput866 net866 vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__buf_8
XFILLER_25_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput877 net1277 vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__buf_8
XFILLER_5_3629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput888 net888 vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_8
XFILLER_28_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput899 net899 vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_8
XFILLER_25_2834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1608 net25 vssd vssd vccd vccd net1608 sky130_fd_sc_hd__buf_6
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1619 net115 vssd vssd vccd vccd net1619 sky130_fd_sc_hd__buf_6
XFILLER_3_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__077__A net963 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_B la_data_in_enable\[38\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_10_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__524__B mprj_logic1\[229\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_B la_data_in_enable\[122\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__540__A net1564 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2172_A mprj_logic1\[153\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input255_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input422_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_525_ net308 net2027 vssd vssd vccd vccd net767 sky130_fd_sc_hd__and2_4
XTAP_2752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__418__C net75 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_456_ net1530 net2149 net1617 vssd vssd vccd vccd net576 sky130_fd_sc_hd__and3b_4
XFILLER_31_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_387_ net297 net1648 net41 vssd vssd vccd vccd net500 sky130_fd_sc_hd__and3b_4
XFILLER_35_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[29\]_B la_data_in_enable\[29\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__434__B net2196 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_B la_data_in_enable\[113\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output474_A net1135 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output739_A net739 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1272_A net1273 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__461__A_N net379 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1537_A net366 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__609__B net1922 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1704_A net1705 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[22\]_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__625__A net1871 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__344__B net1348 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[104\]_B la_data_in_enable\[104\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_14_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput630 net630 vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_8
XANTENNA__360__A net1708 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput641 net641 vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_8
Xoutput652 net652 vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_8
XFILLER_47_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput663 net663 vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_8
XFILLER_9_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput674 net674 vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_8
XFILLER_25_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput685 net685 vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_8
Xwire2106 net2107 vssd vssd vccd vccd net2106 sky130_fd_sc_hd__buf_6
Xoutput696 net696 vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_8
Xwire2117 net2118 vssd vssd vccd vccd net2117 sky130_fd_sc_hd__buf_6
Xwire2128 net2129 vssd vssd vccd vccd net2128 sky130_fd_sc_hd__buf_6
XFILLER_5_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2139 mprj_logic1\[170\] vssd vssd vccd vccd net2139 sky130_fd_sc_hd__buf_6
XFILLER_25_2664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1405 net1406 vssd vssd vccd vccd net1405 sky130_fd_sc_hd__buf_6
Xwire1416 net415 vssd vssd vccd vccd net1416 sky130_fd_sc_hd__buf_6
Xwire1427 net1428 vssd vssd vccd vccd net1427 sky130_fd_sc_hd__buf_6
Xwire1438 net1439 vssd vssd vccd vccd net1438 sky130_fd_sc_hd__buf_6
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1449 net1450 vssd vssd vccd vccd net1449 sky130_fd_sc_hd__buf_6
XFILLER_19_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__519__B net2031 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ net2155 net1412 vssd vssd vccd vccd net875 sky130_fd_sc_hd__and2_4
XFILLER_42_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2018_A mprj_logic1\[268\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__535__A net319 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_241_ mprj_logic1\[408\] net235 vssd vssd vccd vccd la_data_in_enable\[78\] sky130_fd_sc_hd__and2_4
XFILLER_51_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__254__B net250 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_172_ net1857 net259 vssd vssd vccd vccd la_data_in_enable\[9\] sky130_fd_sc_hd__and2_4
XFILLER_49_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input372_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__A_N net1591 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__270__A net1777 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1950 net1951 vssd vssd vccd vccd net1950 sky130_fd_sc_hd__buf_6
XFILLER_19_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1961 net1962 vssd vssd vccd vccd net1961 sky130_fd_sc_hd__buf_6
Xwire1972 mprj_logic1\[294\] vssd vssd vccd vccd net1972 sky130_fd_sc_hd__buf_6
XFILLER_18_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1983 mprj_logic1\[288\] vssd vssd vccd vccd net1983 sky130_fd_sc_hd__buf_6
XFILLER_18_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1994 net1995 vssd vssd vccd vccd net1994 sky130_fd_sc_hd__buf_6
XTAP_3250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_250 net1381 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_508_ net282 net2045 vssd vssd vccd vccd net741 sky130_fd_sc_hd__and2_4
XTAP_2582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1020_A net1021 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1118_A net509 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output689_A net689 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ net1547 net2189 net1334 vssd vssd vccd vccd net558 sky130_fd_sc_hd__and3b_4
XFILLER_31_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output856_A net1258 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1487_A net1488 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__180__A net1845 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1654_A mprj_logic1\[8\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1919_A net1920 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__339__B net1360 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__355__A net1713 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__090__A net991 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput471 net1059 vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__buf_8
XFILLER_9_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput482 net482 vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__buf_8
Xoutput493 net493 vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__buf_8
XFILLER_5_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1202 net1203 vssd vssd vccd vccd net1202 sky130_fd_sc_hd__buf_6
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1213 net918 vssd vssd vccd vccd net1213 sky130_fd_sc_hd__buf_6
XFILLER_47_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1224 net1225 vssd vssd vccd vccd net1224 sky130_fd_sc_hd__buf_6
Xwire1235 net1236 vssd vssd vccd vccd net1235 sky130_fd_sc_hd__buf_6
Xwire1246 net1247 vssd vssd vccd vccd net1246 sky130_fd_sc_hd__buf_6
XFILLER_5_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1257 net858 vssd vssd vccd vccd net1257 sky130_fd_sc_hd__buf_6
Xwire1268 net1269 vssd vssd vccd vccd net1268 sky130_fd_sc_hd__buf_6
XFILLER_38_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1279 net876 vssd vssd vccd vccd net1279 sky130_fd_sc_hd__buf_6
XFILLER_1_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input120_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2135_A mprj_logic1\[173\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input218_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__265__A net1785 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_224_ mprj_logic1\[391\] net217 vssd vssd vccd vccd la_data_in_enable\[61\] sky130_fd_sc_hd__and2_2
XFILLER_7_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_155_ la_data_in_mprj_bar\[8\] vssd vssd vccd vccd net707 sky130_fd_sc_hd__inv_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[1\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_45_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_086_ net992 vssd vssd vccd vccd net595 sky130_fd_sc_hd__inv_2
XFILLER_6_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__C net90 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1068_A net588 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output604_A net604 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1780 net1781 vssd vssd vccd vccd net1780 sky130_fd_sc_hd__buf_6
XANTENNA_wire1235_A net1236 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1791 net1792 vssd vssd vccd vccd net1791 sky130_fd_sc_hd__buf_6
XFILLER_18_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1402_A net1403 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__175__A net1852 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[31\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_37_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1771_A net1772 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1869_A net1870 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__622__B net1879 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__085__A la_data_in_mprj_bar\[102\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2730 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2085_A net2086 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input168_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input335_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1010 net792 vssd vssd vccd vccd net1010 sky130_fd_sc_hd__buf_6
Xwire1021 net778 vssd vssd vccd vccd net1021 sky130_fd_sc_hd__buf_6
Xwire1032 net759 vssd vssd vccd vccd net1032 sky130_fd_sc_hd__buf_6
Xwire1043 net730 vssd vssd vccd vccd net1043 sky130_fd_sc_hd__buf_6
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input29_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1054 net477 vssd vssd vccd vccd net1054 sky130_fd_sc_hd__buf_6
Xwire1065 net465 vssd vssd vccd vccd net1065 sky130_fd_sc_hd__buf_6
XFILLER_1_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1076 net580 vssd vssd vccd vccd net1076 sky130_fd_sc_hd__buf_6
Xwire1087 net1088 vssd vssd vccd vccd net1087 sky130_fd_sc_hd__buf_6
XFILLER_5_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1098 net531 vssd vssd vccd vccd net1098 sky130_fd_sc_hd__buf_6
XFILLER_18_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__426__C net84 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_207_ net1819 net198 vssd vssd vccd vccd la_data_in_enable\[44\] sky130_fd_sc_hd__and2_1
XFILLER_50_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_138_ mprj_dat_i_core_bar\[24\] vssd vssd vccd vccd net897 sky130_fd_sc_hd__clkinv_2
XANTENNA__442__B net2184 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output554_A net554 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_069_ net971 vssd vssd vccd vccd net703 sky130_fd_sc_hd__inv_2
XFILLER_45_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output721_A net721 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output819_A net819 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1352_A net1353 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] la_data_in_enable\[66\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[66\] sky130_fd_sc_hd__nand2_4
XFILLER_1_3440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1617_A net117 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__617__B net1895 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1986_A net1987 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire972_A la_data_in_mprj_bar\[85\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__352__B net1379 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[5\]_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__543__A net1563 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input285_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__262__B net258 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input452_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__437__B net2192 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__418__A_N net331 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1100_A net529 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output769_A net1051 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4418 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output936_A net1150 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1567_A net318 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1734_A mprj_logic1\[458\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1901_A mprj_logic1\[321\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__347__B net1389 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__A net1702 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_610_ net1593 net1919 vssd vssd vccd vccd net734 sky130_fd_sc_hd__and2_4
XTAP_4358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2048_A mprj_logic1\[212\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__A net323 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ net326 mprj_logic1\[246\] vssd vssd vccd vccd net785 sky130_fd_sc_hd__and2_2
XTAP_2912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input200_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__257__B net253 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_472_ net264 net2128 net8 vssd vssd vccd vccd net467 sky130_fd_sc_hd__and3b_4
XTAP_2978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input96_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__273__A net1771 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3866 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output517_A net1111 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput360 la_oenb_mprj[75] vssd vssd vccd vccd net360 sky130_fd_sc_hd__buf_6
XFILLER_42_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput371 la_oenb_mprj[85] vssd vssd vccd vccd net371 sky130_fd_sc_hd__buf_6
XFILLER_23_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput382 la_oenb_mprj[95] vssd vssd vccd vccd net382 sky130_fd_sc_hd__buf_8
XANTENNA_wire1050_A net780 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1148_A net1149 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput393 mprj_adr_o_core[14] vssd vssd vccd vccd net393 sky130_fd_sc_hd__buf_6
XFILLER_36_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] la_data_in_enable\[29\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[29\] sky130_fd_sc_hd__nand2_2
XANTENNA__390__A_N net301 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__183__A net1841 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1684_A net1685 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput801 net999 vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__buf_8
Xoutput812 net812 vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__buf_8
XANTENNA_wire1851_A mprj_logic1\[343\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput823 net823 vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__buf_8
XFILLER_9_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1949_A mprj_logic1\[304\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput834 net995 vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__buf_8
Xoutput845 net845 vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__buf_8
XFILLER_8_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput856 net1258 vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__buf_8
Xoutput867 net867 vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__buf_8
XFILLER_9_3788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput878 net1276 vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput889 net889 vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_8
XFILLER_3_4033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1609 net224 vssd vssd vccd vccd net1609 sky130_fd_sc_hd__buf_4
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__358__A net1710 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3930 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__093__A net989 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input150_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2165_A net2166 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input248_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input415_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__268__A net1780 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ net1575 mprj_logic1\[229\] vssd vssd vccd vccd net766 sky130_fd_sc_hd__and2_4
XTAP_2742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ net1531 net2152 net1618 vssd vssd vccd vccd net575 sky130_fd_sc_hd__and3b_4
XTAP_2797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_386_ net296 net1650 net40 vssd vssd vccd vccd net499 sky130_fd_sc_hd__and3b_4
XFILLER_50_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__434__C net1339 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output467_A net1063 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1098_A net531 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__450__B net2167 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output634_A net634 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1265_A net852 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output801_A net999 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1432_A net1433 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput190 la_iena_mprj[37] vssd vssd vccd vccd net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__178__A net1847 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1899_A net1900 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput620 net620 vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_8
XFILLER_47_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput631 net631 vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_8
XFILLER_9_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__360__B net1368 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput642 net642 vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_8
XFILLER_47_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput653 net653 vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_8
XFILLER_47_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput664 net664 vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_8
XFILLER_28_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput675 net675 vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_8
XFILLER_9_3596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput686 net686 vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_8
Xwire2107 mprj_logic1\[188\] vssd vssd vccd vccd net2107 sky130_fd_sc_hd__buf_6
Xoutput697 net697 vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_8
Xwire2118 mprj_logic1\[183\] vssd vssd vccd vccd net2118 sky130_fd_sc_hd__buf_6
XFILLER_25_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2129 mprj_logic1\[177\] vssd vssd vccd vccd net2129 sky130_fd_sc_hd__buf_6
XFILLER_28_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1406 net1407 vssd vssd vccd vccd net1406 sky130_fd_sc_hd__buf_6
Xwire1417 net1418 vssd vssd vccd vccd net1417 sky130_fd_sc_hd__buf_8
XFILLER_47_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1428 net1429 vssd vssd vccd vccd net1428 sky130_fd_sc_hd__buf_6
Xwire1439 net1440 vssd vssd vccd vccd net1439 sky130_fd_sc_hd__buf_6
XFILLER_3_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__088__A la_data_in_mprj_bar\[105\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_240_ mprj_logic1\[407\] net234 vssd vssd vccd vccd la_data_in_enable\[77\] sky130_fd_sc_hd__and2_4
XANTENNA__535__B net2025 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_171_ net1858 net248 vssd vssd vccd vccd la_data_in_enable\[8\] sky130_fd_sc_hd__and2_2
XFILLER_10_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input198_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__A net337 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input365_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_510 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_irq_gates\[0\] user_irq_core[0] user_irq_enable\[0\] vssd vssd vccd vccd user_irq_bar\[0\]
+ sky130_fd_sc_hd__nand2_1
XANTENNA_input59_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1940 mprj_logic1\[308\] vssd vssd vccd vccd net1940 sky130_fd_sc_hd__buf_6
XFILLER_4_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1951 net1952 vssd vssd vccd vccd net1951 sky130_fd_sc_hd__buf_6
XFILLER_19_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1962 mprj_logic1\[2\] vssd vssd vccd vccd net1962 sky130_fd_sc_hd__buf_6
Xwire1973 net1974 vssd vssd vccd vccd net1973 sky130_fd_sc_hd__buf_6
Xwire1984 net1985 vssd vssd vccd vccd net1984 sky130_fd_sc_hd__buf_6
XTAP_3240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__429__C net88 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1995 mprj_logic1\[282\] vssd vssd vccd vccd net1995 sky130_fd_sc_hd__buf_6
XFILLER_19_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_240 net1754 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 net1575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ net271 net2047 vssd vssd vccd vccd net730 sky130_fd_sc_hd__and2_2
XFILLER_19_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__445__B net2177 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1013_A net1014 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ net1548 net2191 net1335 vssd vssd vccd vccd net556 sky130_fd_sc_hd__and3b_4
XANTENNA_output584_A net1072 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_369_ net260 net1688 net4 vssd vssd vccd vccd net463 sky130_fd_sc_hd__and3b_4
XFILLER_18_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output751_A net1039 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output849_A net1271 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] net1318 vssd vssd vccd vccd la_data_in_mprj_bar\[96\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1647_A mprj_logic1\[93\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__355__B net1376 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput472 net1058 vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__buf_8
XFILLER_47_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput483 net483 vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__buf_8
Xoutput494 net1132 vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__buf_8
XFILLER_5_3257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1203 net1204 vssd vssd vccd vccd net1203 sky130_fd_sc_hd__buf_6
Xwire1214 net1215 vssd vssd vccd vccd net1214 sky130_fd_sc_hd__buf_6
XFILLER_5_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1225 net914 vssd vssd vccd vccd net1225 sky130_fd_sc_hd__buf_6
XFILLER_47_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1236 net1237 vssd vssd vccd vccd net1236 sky130_fd_sc_hd__buf_6
XFILLER_1_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1247 net1248 vssd vssd vccd vccd net1247 sky130_fd_sc_hd__buf_6
XFILLER_5_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1258 net1259 vssd vssd vccd vccd net1258 sky130_fd_sc_hd__buf_6
XFILLER_21_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1269 net1270 vssd vssd vccd vccd net1269 sky130_fd_sc_hd__buf_6
XFILLER_38_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2030_A mprj_logic1\[225\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input113_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2128_A net2129 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__A net331 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__265__B net135 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__451__A_N net1535 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_223_ mprj_logic1\[390\] net216 vssd vssd vccd vccd la_data_in_enable\[60\] sky130_fd_sc_hd__and2_2
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_154_ la_data_in_mprj_bar\[7\] vssd vssd vccd vccd net696 sky130_fd_sc_hd__clkinv_2
XFILLER_13_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__281__A net1755 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_085_ la_data_in_mprj_bar\[102\] vssd vssd vccd vccd net594 sky130_fd_sc_hd__inv_2
XFILLER_49_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1770 mprj_logic1\[441\] vssd vssd vccd vccd net1770 sky130_fd_sc_hd__buf_6
XFILLER_4_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1781 mprj_logic1\[435\] vssd vssd vccd vccd net1781 sky130_fd_sc_hd__buf_6
XFILLER_53_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1792 mprj_logic1\[429\] vssd vssd vccd vccd net1792 sky130_fd_sc_hd__buf_6
XFILLER_15_4000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1130_A net496 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1228_A net944 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output799_A net799 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] la_data_in_enable\[11\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[11\] sky130_fd_sc_hd__nand2_2
XFILLER_15_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] wb_in_enable vssd vssd vccd vccd mprj_dat_i_core_bar\[24\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_50_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1597_A net270 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__191__A net1829 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1764_A mprj_logic1\[444\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1931_A net1932 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] la_data_in_enable\[122\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[122\] sky130_fd_sc_hd__nand2_2
XFILLER_6_2876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__A_N net1602 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__366__A net1694 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2078_A mprj_logic1\[198\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1000 net1001 vssd vssd vccd vccd net1000 sky130_fd_sc_hd__buf_6
Xwire1011 net1012 vssd vssd vccd vccd net1011 sky130_fd_sc_hd__buf_6
XFILLER_40_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1022 net1023 vssd vssd vccd vccd net1022 sky130_fd_sc_hd__buf_6
XANTENNA_input230_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1033 net757 vssd vssd vccd vccd net1033 sky130_fd_sc_hd__buf_6
XANTENNA_input328_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1044 net846 vssd vssd vccd vccd net1044 sky130_fd_sc_hd__buf_6
XFILLER_2_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1055 net476 vssd vssd vccd vccd net1055 sky130_fd_sc_hd__buf_6
XFILLER_53_4509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1066 net464 vssd vssd vccd vccd net1066 sky130_fd_sc_hd__buf_6
XFILLER_2_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1077 net578 vssd vssd vccd vccd net1077 sky130_fd_sc_hd__buf_6
Xwire1088 net541 vssd vssd vccd vccd net1088 sky130_fd_sc_hd__buf_6
Xwire1099 net530 vssd vssd vccd vccd net1099 sky130_fd_sc_hd__buf_6
XFILLER_28_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__276__A net1765 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_206_ net1820 net197 vssd vssd vccd vccd la_data_in_enable\[43\] sky130_fd_sc_hd__and2_1
XFILLER_10_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_137_ mprj_dat_i_core_bar\[23\] vssd vssd vccd vccd net896 sky130_fd_sc_hd__clkinv_2
XFILLER_8_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__442__C net1631 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_068_ net972 vssd vssd vccd vccd net702 sky130_fd_sc_hd__inv_2
XFILLER_45_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output547_A net1080 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1080_A net547 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1178_A net1179 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output714_A net714 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1345_A net452 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] la_data_in_enable\[59\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[59\] sky130_fd_sc_hd__nand2_2
XFILLER_1_2740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1512_A net1513 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1716 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__A net1837 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1881_A net1882 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1979_A net1980 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__096__A net986 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__543__B mprj_logic1\[248\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input180_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2195_A mprj_logic1\[13\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input445_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input41_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__437__C net1336 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output497_A net1129 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__B net2159 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1295_A net1296 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output831_A net831 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output929_A net1174 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1462_A net1463 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1727_A net1728 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__B net1365 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__B mprj_logic1\[243\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_540_ net1564 mprj_logic1\[245\] vssd vssd vccd vccd net784 sky130_fd_sc_hd__and2_4
XTAP_2913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ net1605 net2130 net7 vssd vssd vccd vccd net466 sky130_fd_sc_hd__and3b_4
XFILLER_32_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2110_A net2111 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2208_A net2209 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__A net340 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input395_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__273__B net144 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input89_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput350 la_oenb_mprj[66] vssd vssd vccd vccd net350 sky130_fd_sc_hd__buf_6
Xinput361 la_oenb_mprj[76] vssd vssd vccd vccd net361 sky130_fd_sc_hd__buf_6
Xinput372 la_oenb_mprj[86] vssd vssd vccd vccd net372 sky130_fd_sc_hd__buf_6
XFILLER_40_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput383 la_oenb_mprj[96] vssd vssd vccd vccd net383 sky130_fd_sc_hd__buf_6
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput394 mprj_adr_o_core[15] vssd vssd vccd vccd net394 sky130_fd_sc_hd__buf_6
XFILLER_53_4103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__448__B net2171 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1210_A net919 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output781_A net781 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1308_A net1309 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output879_A net1274 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput802 net1048 vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__buf_8
Xoutput813 net1047 vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__buf_8
Xoutput824 net1046 vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__buf_8
XFILLER_25_4249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput835 net1045 vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__buf_8
XFILLER_6_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput846 net1044 vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__buf_8
XFILLER_29_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput857 net857 vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__buf_8
XFILLER_5_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1844_A mprj_logic1\[348\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput868 net868 vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__buf_8
XFILLER_42_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput879 net1274 vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__buf_8
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__358__B net1370 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_2244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input143_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2060_A net2061 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2158_A mprj_logic1\[159\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1886 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__549__A net335 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__268__B net138 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input310_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input408_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_523_ net306 net2028 vssd vssd vccd vccd net765 sky130_fd_sc_hd__and2_4
XFILLER_22_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_454_ net1532 net2156 net1619 vssd vssd vccd vccd net574 sky130_fd_sc_hd__and3b_4
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__284__A net1749 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_385_ net295 net1652 net39 vssd vssd vccd vccd net498 sky130_fd_sc_hd__and3b_4
XFILLER_9_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__450__C net1623 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1160_A net1161 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1258_A net1259 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput180 la_iena_mprj[28] vssd vssd vccd vccd net180 sky130_fd_sc_hd__buf_4
XFILLER_42_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput191 la_iena_mprj[38] vssd vssd vccd vccd net191 sky130_fd_sc_hd__clkbuf_4
XANTENNA__178__B net166 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1425_A net1426 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] la_data_in_enable\[41\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[41\] sky130_fd_sc_hd__nand2_2
XFILLER_18_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__194__A net1825 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1961_A net1962 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput610 net610 vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_8
Xoutput621 net621 vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_8
Xoutput632 net632 vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_8
Xoutput643 net643 vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_8
XFILLER_9_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput654 net654 vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_8
XFILLER_5_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput665 net665 vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] la_data_in_enable\[3\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[3\] sky130_fd_sc_hd__nand2_1
XFILLER_47_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput676 net676 vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_8
XFILLER_28_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2108 net2109 vssd vssd vccd vccd net2108 sky130_fd_sc_hd__buf_6
Xoutput687 net687 vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_8
Xoutput698 net698 vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_8
Xwire2119 net2120 vssd vssd vccd vccd net2119 sky130_fd_sc_hd__buf_6
XFILLER_42_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1407 net1408 vssd vssd vccd vccd net1407 sky130_fd_sc_hd__buf_6
XFILLER_25_2677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1418 net1419 vssd vssd vccd vccd net1418 sky130_fd_sc_hd__buf_6
Xwire1429 net1430 vssd vssd vccd vccd net1429 sky130_fd_sc_hd__buf_6
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_170_ net1859 net237 vssd vssd vccd vccd la_data_in_enable\[7\] sky130_fd_sc_hd__and2_2
XFILLER_32_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__B mprj_logic1\[256\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input260_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input358_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_566 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__380__A_N net282 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__279__A net1759 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1930 mprj_logic1\[312\] vssd vssd vccd vccd net1930 sky130_fd_sc_hd__buf_6
Xwire1941 net1942 vssd vssd vccd vccd net1941 sky130_fd_sc_hd__buf_6
XFILLER_4_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1952 mprj_logic1\[303\] vssd vssd vccd vccd net1952 sky130_fd_sc_hd__buf_6
XFILLER_18_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1963 net1964 vssd vssd vccd vccd net1963 sky130_fd_sc_hd__buf_6
Xwire1974 mprj_logic1\[293\] vssd vssd vccd vccd net1974 sky130_fd_sc_hd__buf_6
XFILLER_20_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1985 mprj_logic1\[287\] vssd vssd vccd vccd net1985 sky130_fd_sc_hd__buf_6
XFILLER_19_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1996 net1997 vssd vssd vccd vccd net1996 sky130_fd_sc_hd__buf_6
XFILLER_34_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_230 mprj_logic1\[84\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_241 net1762 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_506_ net387 net2049 vssd vssd vccd vccd net846 sky130_fd_sc_hd__and2_4
XANTENNA_252 mprj_logic1\[78\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3558 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ net1549 net2192 net1336 vssd vssd vccd vccd net555 sky130_fd_sc_hd__and3b_4
XFILLER_50_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__445__C net1628 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_368_ net1690 net1358 vssd vssd vccd vccd net937 sky130_fd_sc_hd__and2_2
XFILLER_31_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output577_A net577 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_299_ mprj_logic1\[4\] net1342 vssd vssd vccd vccd net949 sky130_fd_sc_hd__and2_4
XFILLER_31_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__461__B net2142 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output744_A net744 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1375_A net431 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] net1325 vssd vssd vccd vccd la_data_in_mprj_bar\[89\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1542_A net360 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__189__A net1831 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1807_A mprj_logic1\[412\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire995_A net834 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__B net1684 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput473 net1057 vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__buf_8
Xoutput484 net484 vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__buf_8
XFILLER_47_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput495 net1131 vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__buf_8
XFILLER_5_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1204 net921 vssd vssd vccd vccd net1204 sky130_fd_sc_hd__buf_6
XFILLER_9_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1215 net1216 vssd vssd vccd vccd net1215 sky130_fd_sc_hd__buf_6
XFILLER_9_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__099__A la_data_in_mprj_bar\[116\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1226 net1227 vssd vssd vccd vccd net1226 sky130_fd_sc_hd__buf_6
XFILLER_19_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1237 net941 vssd vssd vccd vccd net1237 sky130_fd_sc_hd__buf_6
XFILLER_47_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1248 net935 vssd vssd vccd vccd net1248 sky130_fd_sc_hd__buf_6
XFILLER_47_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1259 net856 vssd vssd vccd vccd net1259 sky130_fd_sc_hd__buf_6
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__B net2023 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_222_ mprj_logic1\[389\] net214 vssd vssd vccd vccd la_data_in_enable\[59\] sky130_fd_sc_hd__and2_2
XFILLER_10_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__562__A net1552 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_153_ la_data_in_mprj_bar\[6\] vssd vssd vccd vccd net685 sky130_fd_sc_hd__clkinv_2
XFILLER_7_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input71_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_084_ la_data_in_mprj_bar\[101\] vssd vssd vccd vccd net593 sky130_fd_sc_hd__inv_4
XFILLER_45_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1760 mprj_logic1\[446\] vssd vssd vccd vccd net1760 sky130_fd_sc_hd__buf_6
XFILLER_20_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1771 net1772 vssd vssd vccd vccd net1771 sky130_fd_sc_hd__buf_6
XFILLER_19_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1782 net1783 vssd vssd vccd vccd net1782 sky130_fd_sc_hd__buf_6
Xwire1793 net1794 vssd vssd vccd vccd net1793 sky130_fd_sc_hd__buf_6
XFILLER_19_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__456__B net2149 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1123_A net504 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output861_A net861 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[17\]
+ sky130_fd_sc_hd__nand2_4
XANTENNA_wire1492_A net1493 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__191__B net180 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1757_A net1758 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1924_A mprj_logic1\[314\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] la_data_in_enable\[115\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[115\] sky130_fd_sc_hd__nand2_2
XFILLER_39_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__366__B net1362 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_B net1319 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1001 net800 vssd vssd vccd vccd net1001 sky130_fd_sc_hd__buf_6
XFILLER_5_2332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1012 net790 vssd vssd vccd vccd net1012 sky130_fd_sc_hd__buf_6
Xwire1023 net774 vssd vssd vccd vccd net1023 sky130_fd_sc_hd__buf_6
XFILLER_25_2282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1034 net756 vssd vssd vccd vccd net1034 sky130_fd_sc_hd__buf_6
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1045 net835 vssd vssd vccd vccd net1045 sky130_fd_sc_hd__buf_6
XFILLER_47_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1056 net475 vssd vssd vccd vccd net1056 sky130_fd_sc_hd__buf_6
XANTENNA_wire2140_A mprj_logic1\[169\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1067 net589 vssd vssd vccd vccd net1067 sky130_fd_sc_hd__buf_6
XANTENNA_input223_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1078 net549 vssd vssd vccd vccd net1078 sky130_fd_sc_hd__buf_6
XFILLER_38_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1089 net540 vssd vssd vccd vccd net1089 sky130_fd_sc_hd__buf_6
XANTENNA__557__A net344 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__276__B net147 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[86\]_B net1328 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__292__A net1729 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_205_ net1821 net196 vssd vssd vccd vccd la_data_in_enable\[42\] sky130_fd_sc_hd__and2_1
XFILLER_11_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_136_ mprj_dat_i_core_bar\[22\] vssd vssd vccd vccd net895 sky130_fd_sc_hd__clkinv_2
XFILLER_10_2540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_067_ net973 vssd vssd vccd vccd net701 sky130_fd_sc_hd__inv_2
XFILLER_45_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1073_A net583 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_4071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1590 net278 vssd vssd vccd vccd net1590 sky130_fd_sc_hd__buf_8
XFILLER_0_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__B net1615 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1505_A net1506 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[77\]_B la_data_in_enable\[77\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_50_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1874_A net1875 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__441__A_N net1545 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input173_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2188_A mprj_logic1\[145\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input340_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input438_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input34_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__287__A net1742 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__C net1620 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output657_A net657 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_119_ mprj_dat_i_core_bar\[5\] vssd vssd vccd vccd net908 sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1190_A net1191 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__A_N net382 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output824_A net1046 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1455_A net1456 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] la_data_in_enable\[71\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[71\] sky130_fd_sc_hd__nand2_4
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1622_A net112 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__197__A mprj_logic1\[364\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1991_A mprj_logic1\[284\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_470_ net1606 net2132 net6 vssd vssd vccd vccd net465 sky130_fd_sc_hd__and3b_4
XTAP_2958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[125\]_B la_data_in_enable\[125\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__B mprj_logic1\[259\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2103_A net2104 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input290_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input388_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__487__A_N net1588 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A net1544 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3982 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput340 la_oenb_mprj[57] vssd vssd vccd vccd net340 sky130_fd_sc_hd__buf_6
XFILLER_2_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput351 la_oenb_mprj[67] vssd vssd vccd vccd net351 sky130_fd_sc_hd__buf_6
Xinput362 la_oenb_mprj[77] vssd vssd vccd vccd net362 sky130_fd_sc_hd__buf_6
XFILLER_3_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput373 la_oenb_mprj[87] vssd vssd vccd vccd net373 sky130_fd_sc_hd__buf_6
Xinput384 la_oenb_mprj[97] vssd vssd vccd vccd net384 sky130_fd_sc_hd__buf_4
Xinput395 mprj_adr_o_core[16] vssd vssd vccd vccd net395 sky130_fd_sc_hd__buf_6
XFILLER_53_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__448__C net1625 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1036_A net754 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_599_ net1605 net1948 vssd vssd vccd vccd net722 sky130_fd_sc_hd__and2_4
XFILLER_43_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__B net2140 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_B la_data_in_enable\[116\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_4468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1203_A net1204 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output774_A net1022 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output941_A net1235 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput803 net997 vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__buf_8
Xoutput814 net814 vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__buf_8
Xoutput825 net825 vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput836 net994 vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__buf_8
Xoutput847 net847 vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_8
Xoutput858 net1257 vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_3_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput869 net869 vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1837_A net1838 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[25\]_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1366 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[107\]_B net1315 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__374__B net1678 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2522 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__549__B mprj_logic1\[254\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2053_A net2054 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input136_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[16\]_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_522_ net305 mprj_logic1\[227\] vssd vssd vccd vccd net764 sky130_fd_sc_hd__and2_1
XFILLER_22_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input303_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__565__A net1549 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_453_ net1533 net2159 net1620 vssd vssd vccd vccd net573 sky130_fd_sc_hd__and3b_4
XTAP_2777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_384_ net294 net1655 net38 vssd vssd vccd vccd net497 sky130_fd_sc_hd__and3b_4
XFILLER_35_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output522_A net1106 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__459__B net2144 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1153_A net936 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput170 la_iena_mprj[19] vssd vssd vccd vccd net170 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput181 la_iena_mprj[29] vssd vssd vccd vccd net181 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput192 la_iena_mprj[39] vssd vssd vccd vccd net192 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1320_A la_data_in_enable\[94\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1418_A net1419 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] la_data_in_enable\[34\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[34\] sky130_fd_sc_hd__nand2_1
XFILLER_53_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__194__B net184 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1787_A net1788 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1954_A mprj_logic1\[302\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput600 net600 vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_8
XFILLER_29_4194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput611 net611 vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_8
Xoutput622 net622 vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput633 net633 vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_8
XFILLER_44_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput644 net644 vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_8
Xoutput655 net655 vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_8
XFILLER_9_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput666 net666 vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_8
XFILLER_29_2770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput677 net677 vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_8
Xoutput688 net688 vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_8
Xwire2109 mprj_logic1\[187\] vssd vssd vccd vccd net2109 sky130_fd_sc_hd__buf_6
XFILLER_47_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput699 net699 vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_8
Xwire1408 net417 vssd vssd vccd vccd net1408 sky130_fd_sc_hd__buf_6
XFILLER_42_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1419 net1420 vssd vssd vccd vccd net1419 sky130_fd_sc_hd__buf_6
XFILLER_25_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__369__B net1688 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2170_A mprj_logic1\[154\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input253_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input420_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__279__B net150 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1920 net1921 vssd vssd vccd vccd net1920 sky130_fd_sc_hd__buf_6
XFILLER_19_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1931 net1932 vssd vssd vccd vccd net1931 sky130_fd_sc_hd__buf_6
XFILLER_1_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1942 mprj_logic1\[307\] vssd vssd vccd vccd net1942 sky130_fd_sc_hd__buf_6
Xwire1953 net1954 vssd vssd vccd vccd net1953 sky130_fd_sc_hd__buf_6
XFILLER_19_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1964 mprj_logic1\[299\] vssd vssd vccd vccd net1964 sky130_fd_sc_hd__buf_6
XFILLER_18_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1975 mprj_logic1\[292\] vssd vssd vccd vccd net1975 sky130_fd_sc_hd__buf_6
XFILLER_19_4330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1986 net1987 vssd vssd vccd vccd net1986 sky130_fd_sc_hd__buf_6
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1997 mprj_logic1\[281\] vssd vssd vccd vccd net1997 sky130_fd_sc_hd__buf_6
XFILLER_19_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_220 net2133 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_231 mprj_logic1\[94\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ net376 net2051 vssd vssd vccd vccd net835 sky130_fd_sc_hd__and2_2
XTAP_2552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_242 net1764 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 net1381 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_436_ net1550 net2193 net1337 vssd vssd vccd vccd net554 sky130_fd_sc_hd__and3b_4
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_367_ net1692 net1359 vssd vssd vccd vccd net936 sky130_fd_sc_hd__and2_2
XFILLER_32_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_298_ net1811 net1394 vssd vssd vccd vccd net880 sky130_fd_sc_hd__and2_2
XANTENNA_output472_A net1058 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__461__C net123 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output737_A net737 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1270_A net850 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1368_A net436 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__189__B net1612 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1535_A net368 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1702_A net1703 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__C net54 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput463 net1145 vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__buf_8
Xoutput474 net1135 vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__buf_8
Xoutput485 net1133 vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__buf_8
Xoutput496 net1130 vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__buf_8
XFILLER_9_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1205 net1206 vssd vssd vccd vccd net1205 sky130_fd_sc_hd__buf_6
XFILLER_9_1960 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1216 net917 vssd vssd vccd vccd net1216 sky130_fd_sc_hd__buf_6
Xwire1227 net1228 vssd vssd vccd vccd net1227 sky130_fd_sc_hd__buf_6
XFILLER_21_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1238 net1239 vssd vssd vccd vccd net1238 sky130_fd_sc_hd__buf_6
Xwire1249 net1250 vssd vssd vccd vccd net1249 sky130_fd_sc_hd__buf_6
XFILLER_38_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2016_A mprj_logic1\[270\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_221_ mprj_logic1\[388\] net213 vssd vssd vccd vccd la_data_in_enable\[58\] sky130_fd_sc_hd__and2_1
XFILLER_10_4146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_152_ la_data_in_mprj_bar\[5\] vssd vssd vccd vccd net674 sky130_fd_sc_hd__clkinv_2
XANTENNA__562__B net2019 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_083_ net993 vssd vssd vccd vccd net592 sky130_fd_sc_hd__clkinv_4
XANTENNA_input370_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input64_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1750 mprj_logic1\[451\] vssd vssd vccd vccd net1750 sky130_fd_sc_hd__buf_6
Xwire1761 net1762 vssd vssd vccd vccd net1761 sky130_fd_sc_hd__buf_6
Xwire1772 mprj_logic1\[440\] vssd vssd vccd vccd net1772 sky130_fd_sc_hd__buf_6
XFILLER_18_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1783 mprj_logic1\[434\] vssd vssd vccd vccd net1783 sky130_fd_sc_hd__buf_6
XFILLER_37_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1794 mprj_logic1\[428\] vssd vssd vccd vccd net1794 sky130_fd_sc_hd__buf_6
XTAP_3050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__456__C net1617 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1116_A net511 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output687_A net687 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ net333 mprj_logic1\[124\] net77 vssd vssd vccd vccd net536 sky130_fd_sc_hd__and3b_2
XFILLER_50_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__B net2128 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output854_A net1261 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1485_A net1486 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1652_A net1653 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1917_A net1918 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] la_data_in_enable\[108\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[108\] sky130_fd_sc_hd__nand2_2
XFILLER_17_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__A_N net299 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__382__B net1659 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[8\]_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1002 net1003 vssd vssd vccd vccd net1002 sky130_fd_sc_hd__buf_6
XFILLER_40_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1013 net1014 vssd vssd vccd vccd net1013 sky130_fd_sc_hd__buf_6
XFILLER_2_3933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1024 net773 vssd vssd vccd vccd net1024 sky130_fd_sc_hd__buf_6
Xwire1035 net755 vssd vssd vccd vccd net1035 sky130_fd_sc_hd__buf_6
XFILLER_5_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1046 net824 vssd vssd vccd vccd net1046 sky130_fd_sc_hd__buf_6
XFILLER_38_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1057 net473 vssd vssd vccd vccd net1057 sky130_fd_sc_hd__buf_6
XFILLER_47_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1068 net588 vssd vssd vccd vccd net1068 sky130_fd_sc_hd__buf_6
XFILLER_0_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1079 net548 vssd vssd vccd vccd net1079 sky130_fd_sc_hd__buf_6
XFILLER_38_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2133_A net2134 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input216_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__573__A net1541 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_204_ net1822 net195 vssd vssd vccd vccd la_data_in_enable\[41\] sky130_fd_sc_hd__and2_1
XFILLER_12_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__292__B net461 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_135_ mprj_dat_i_core_bar\[21\] vssd vssd vccd vccd net894 sky130_fd_sc_hd__inv_2
XFILLER_49_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_066_ net974 vssd vssd vccd vccd net700 sky130_fd_sc_hd__inv_2
XFILLER_10_2596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__467__B net2136 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1580 net289 vssd vssd vccd vccd net1580 sky130_fd_sc_hd__buf_6
XFILLER_21_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1591 net277 vssd vssd vccd vccd net1591 sky130_fd_sc_hd__buf_8
XANTENNA_wire1233_A net1234 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__393__A_N net304 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1400_A net419 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1867_A net1868 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__B net1670 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input166_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2083_A net2084 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input333_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__A net1546 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input27_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__287__B net159 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_118_ mprj_dat_i_core_bar\[4\] vssd vssd vccd vccd net907 sky130_fd_sc_hd__clkinv_2
XFILLER_29_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output552_A net552 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_049_ la_data_in_mprj_bar\[66\] vssd vssd vccd vccd net681 sky130_fd_sc_hd__clkinv_2
XFILLER_7_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1183_A net1184 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output817_A net817 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1350_A net1351 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1448_A net1449 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] la_data_in_enable\[64\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[64\] sky130_fd_sc_hd__nand2_4
XFILLER_1_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1984_A net1985 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire970_A la_data_in_mprj_bar\[87\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input283_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__B net2009 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput330 la_oenb_mprj[48] vssd vssd vccd vccd net330 sky130_fd_sc_hd__buf_6
XFILLER_2_4261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__298__A net1811 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput341 la_oenb_mprj[58] vssd vssd vccd vccd net341 sky130_fd_sc_hd__buf_6
XFILLER_48_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput352 la_oenb_mprj[68] vssd vssd vccd vccd net352 sky130_fd_sc_hd__buf_6
Xinput363 la_oenb_mprj[78] vssd vssd vccd vccd net363 sky130_fd_sc_hd__buf_6
Xinput374 la_oenb_mprj[88] vssd vssd vccd vccd net374 sky130_fd_sc_hd__buf_6
XFILLER_29_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput385 la_oenb_mprj[98] vssd vssd vccd vccd net385 sky130_fd_sc_hd__buf_6
XFILLER_48_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput396 mprj_adr_o_core[17] vssd vssd vccd vccd net396 sky130_fd_sc_hd__buf_6
XFILLER_18_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1029_A net762 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_598_ net1606 net1950 vssd vssd vccd vccd net721 sky130_fd_sc_hd__and2_4
XFILLER_38_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__C net126 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__A_N net1555 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output767_A net1025 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1398_A net1399 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__480__B net2112 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1 la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput804 net996 vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__buf_8
XANTENNA_output934_A net1154 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput815 net815 vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__buf_8
Xoutput826 net826 vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__buf_8
XFILLER_42_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput837 net837 vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__buf_8
XFILLER_6_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1565_A net322 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput848 net848 vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__buf_8
XFILLER_28_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput859 net859 vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_42_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_2985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1732_A net1733 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[25\]_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__390__B net1643 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[16\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2046_A mprj_logic1\[213\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input129_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1994 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_521_ net304 net2029 vssd vssd vccd vccd net763 sky130_fd_sc_hd__and2_2
XTAP_2723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__565__B net2016 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_452_ net1534 net2162 net1621 vssd vssd vccd vccd net572 sky130_fd_sc_hd__and3b_4
XFILLER_17_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__454__A_N net1532 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_383_ net293 net1657 net37 vssd vssd vccd vccd net496 sky130_fd_sc_hd__and3b_4
XFILLER_25_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input94_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__A net1533 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__459__C net121 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output515_A net1113 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput160 la_iena_mprj[125] vssd vssd vccd vccd net160 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput171 la_iena_mprj[1] vssd vssd vccd vccd net171 sky130_fd_sc_hd__clkbuf_4
Xinput182 la_iena_mprj[2] vssd vssd vccd vccd net182 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput193 la_iena_mprj[3] vssd vssd vccd vccd net193 sky130_fd_sc_hd__clkbuf_4
XTAP_4670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1146_A net1147 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__475__B net2123 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1313_A la_data_in_enable\[123\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] la_data_in_enable\[27\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[27\] sky130_fd_sc_hd__nand2_2
XFILLER_18_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1682_A net1683 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput601 net601 vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_8
XFILLER_25_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput612 net612 vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_8
XFILLER_47_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput623 net623 vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_8
Xoutput634 net634 vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_8
Xoutput645 net645 vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_8
XFILLER_47_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput656 net656 vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_8
XFILLER_25_3336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput667 net667 vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_8
XFILLER_29_2782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput678 net678 vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_8
Xoutput689 net689 vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_8
XFILLER_42_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1409 net1410 vssd vssd vccd vccd net1409 sky130_fd_sc_hd__buf_6
XFILLER_41_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__369__C net4 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__477__A_N net269 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__385__B net1652 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input246_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2163_A net2164 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1910 mprj_logic1\[318\] vssd vssd vccd vccd net1910 sky130_fd_sc_hd__buf_6
Xwire1921 mprj_logic1\[315\] vssd vssd vccd vccd net1921 sky130_fd_sc_hd__buf_6
XFILLER_41_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1932 net1933 vssd vssd vccd vccd net1932 sky130_fd_sc_hd__buf_6
XFILLER_46_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1943 net1944 vssd vssd vccd vccd net1943 sky130_fd_sc_hd__buf_6
Xwire1954 mprj_logic1\[302\] vssd vssd vccd vccd net1954 sky130_fd_sc_hd__buf_6
XTAP_3210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1965 net1966 vssd vssd vccd vccd net1965 sky130_fd_sc_hd__buf_6
XFILLER_19_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1976 mprj_logic1\[291\] vssd vssd vccd vccd net1976 sky130_fd_sc_hd__buf_6
XANTENNA_input413_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1987 mprj_logic1\[286\] vssd vssd vccd vccd net1987 sky130_fd_sc_hd__buf_6
XANTENNA__576__A net1538 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1998 net1999 vssd vssd vccd vccd net1998 sky130_fd_sc_hd__buf_6
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 net1960 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_221 net2134 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_504_ net365 net2052 vssd vssd vccd vccd net824 sky130_fd_sc_hd__and2_4
XANTENNA_232 net26 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__295__B net2203 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 net1790 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 net1575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ net1551 net2194 net1338 vssd vssd vccd vccd net553 sky130_fd_sc_hd__and3b_4
XFILLER_37_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_366_ net1694 net1362 vssd vssd vccd vccd net934 sky130_fd_sc_hd__and2_2
XFILLER_31_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_297_ net1959 net2 vssd vssd vccd vccd net956 sky130_fd_sc_hd__and2_2
XFILLER_35_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output465_A net1065 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1096_A net533 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1263_A net853 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1430_A net1431 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1897_A mprj_logic1\[322\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput464 net1066 vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput475 net1056 vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__buf_8
XFILLER_9_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput486 net486 vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__buf_8
Xoutput497 net1129 vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__buf_8
XFILLER_5_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1206 net1207 vssd vssd vccd vccd net1206 sky130_fd_sc_hd__buf_6
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1217 net1218 vssd vssd vccd vccd net1217 sky130_fd_sc_hd__buf_6
XFILLER_47_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1228 net944 vssd vssd vccd vccd net1228 sky130_fd_sc_hd__buf_6
XFILLER_41_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1239 net1240 vssd vssd vccd vccd net1239 sky130_fd_sc_hd__buf_6
XFILLER_28_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_220_ mprj_logic1\[387\] net212 vssd vssd vccd vccd la_data_in_enable\[57\] sky130_fd_sc_hd__and2_2
XFILLER_10_4125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2009_A mprj_logic1\[275\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_151_ la_data_in_mprj_bar\[4\] vssd vssd vccd vccd net663 sky130_fd_sc_hd__clkinv_2
XANTENNA_input196_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_082_ net961 vssd vssd vccd vccd net717 sky130_fd_sc_hd__clkinv_4
XFILLER_49_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input363_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input57_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1740 net1741 vssd vssd vccd vccd net1740 sky130_fd_sc_hd__buf_6
XFILLER_1_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1751 net1752 vssd vssd vccd vccd net1751 sky130_fd_sc_hd__buf_6
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1762 mprj_logic1\[445\] vssd vssd vccd vccd net1762 sky130_fd_sc_hd__buf_6
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1773 net1774 vssd vssd vccd vccd net1773 sky130_fd_sc_hd__buf_6
XFILLER_1_2946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1784 mprj_logic1\[433\] vssd vssd vccd vccd net1784 sky130_fd_sc_hd__buf_6
XTAP_3040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1795 net1796 vssd vssd vccd vccd net1795 sky130_fd_sc_hd__buf_6
XTAP_3051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_418_ net331 mprj_logic1\[123\] net75 vssd vssd vccd vccd net534 sky130_fd_sc_hd__and3b_4
XFILLER_42_792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1011_A net1012 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output582_A net1074 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1109_A net519 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_349_ mprj_logic1\[54\] net1385 vssd vssd vccd vccd net916 sky130_fd_sc_hd__and2_4
XFILLER_35_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1478_A net1479 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] net1320 vssd vssd vccd vccd la_data_in_mprj_bar\[94\]
+ sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1645_A mprj_logic1\[94\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1812_A mprj_logic1\[39\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__382__C net36 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[8\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1003 net798 vssd vssd vccd vccd net1003 sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[8\]_B la_data_in_enable\[8\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1014 net786 vssd vssd vccd vccd net1014 sky130_fd_sc_hd__buf_6
XFILLER_38_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1025 net767 vssd vssd vccd vccd net1025 sky130_fd_sc_hd__buf_6
XFILLER_9_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1036 net754 vssd vssd vccd vccd net1036 sky130_fd_sc_hd__buf_6
Xwire1047 net813 vssd vssd vccd vccd net1047 sky130_fd_sc_hd__buf_6
Xwire1058 net472 vssd vssd vccd vccd net1058 sky130_fd_sc_hd__buf_6
Xwire1069 net587 vssd vssd vccd vccd net1069 sky130_fd_sc_hd__buf_6
XFILLER_38_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input111_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input209_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2126_A net2127 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__573__B net2003 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_203_ mprj_logic1\[370\] net194 vssd vssd vccd vccd la_data_in_enable\[40\] sky130_fd_sc_hd__and2_2
XFILLER_10_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_134_ mprj_dat_i_core_bar\[20\] vssd vssd vccd vccd net893 sky130_fd_sc_hd__inv_2
XFILLER_10_2520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_065_ la_data_in_mprj_bar\[82\] vssd vssd vccd vccd net699 sky130_fd_sc_hd__clkinv_2
XFILLER_49_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1059_A net471 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1570 net313 vssd vssd vccd vccd net1570 sky130_fd_sc_hd__buf_6
XFILLER_39_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1581 net288 vssd vssd vccd vccd net1581 sky130_fd_sc_hd__buf_6
Xwire1592 net276 vssd vssd vccd vccd net1592 sky130_fd_sc_hd__buf_8
XFILLER_0_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1226_A net1227 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output797_A net1004 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__B net2105 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] net1310 vssd vssd vccd vccd mprj_dat_i_core_bar\[22\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_50_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1762_A mprj_logic1\[445\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] la_data_in_enable\[120\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[120\] sky130_fd_sc_hd__nand2_4
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__C net120 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__393__B net1637 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2076_A net2077 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input159_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__B net2012 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input326_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__584__A net1530 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_117_ mprj_dat_i_core_bar\[3\] vssd vssd vccd vccd net906 sky130_fd_sc_hd__clkinv_2
XFILLER_29_3846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_048_ la_data_in_mprj_bar\[65\] vssd vssd vccd vccd net680 sky130_fd_sc_hd__clkinv_2
XFILLER_4_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output545_A net1081 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1176_A net1177 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output712_A net712 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__478__B net2117 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1343_A net458 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2090 mprj_logic1\[194\] vssd vssd vccd vccd net2090 sky130_fd_sc_hd__buf_6
XFILLER_26_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] la_data_in_enable\[57\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[57\] sky130_fd_sc_hd__nand2_2
XFILLER_36_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1510_A net1511 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_39_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1977_A net1978 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__388__B net1646 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2193_A mprj_logic1\[141\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input276_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__383__A_N net293 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input443_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__579__A net1535 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput320 la_oenb_mprj[39] vssd vssd vccd vccd net320 sky130_fd_sc_hd__clkbuf_4
Xinput331 la_oenb_mprj[49] vssd vssd vccd vccd net331 sky130_fd_sc_hd__buf_4
XFILLER_0_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput342 la_oenb_mprj[59] vssd vssd vccd vccd net342 sky130_fd_sc_hd__buf_4
XANTENNA__298__B net1394 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput353 la_oenb_mprj[69] vssd vssd vccd vccd net353 sky130_fd_sc_hd__buf_6
XFILLER_48_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput364 la_oenb_mprj[79] vssd vssd vccd vccd net364 sky130_fd_sc_hd__buf_6
Xinput375 la_oenb_mprj[89] vssd vssd vccd vccd net375 sky130_fd_sc_hd__clkbuf_4
XFILLER_29_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput386 la_oenb_mprj[99] vssd vssd vccd vccd net386 sky130_fd_sc_hd__buf_6
Xinput397 mprj_adr_o_core[18] vssd vssd vccd vccd net397 sky130_fd_sc_hd__buf_6
XFILLER_48_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_597_ net1607 net1953 vssd vssd vccd vccd net720 sky130_fd_sc_hd__and2_4
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output495_A net1131 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output662_A net662 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__480__C net17 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2 la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput805 net805 vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__buf_8
XFILLER_47_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput816 net816 vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__buf_8
Xoutput827 net827 vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__buf_8
Xoutput838 net838 vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__buf_8
XFILLER_42_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output927_A net1182 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput849 net1271 vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__buf_8
XFILLER_6_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1460_A net1461 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1558_A net334 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1725_A net951 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_520_ net303 net2030 vssd vssd vccd vccd net762 sky130_fd_sc_hd__and2_4
XTAP_2702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2039_A mprj_logic1\[217\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_451_ net1535 net2165 net1622 vssd vssd vccd vccd net571 sky130_fd_sc_hd__and3b_4
XTAP_2757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_382_ net292 net1659 net36 vssd vssd vccd vccd net495 sky130_fd_sc_hd__and3b_4
XFILLER_15_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2206_A net2207 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input393_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__581__B net1986 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input87_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__102__A la_data_in_mprj_bar\[119\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput150 la_iena_mprj[116] vssd vssd vccd vccd net150 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput161 la_iena_mprj[126] vssd vssd vccd vccd net161 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput172 la_iena_mprj[20] vssd vssd vccd vccd net172 sky130_fd_sc_hd__clkbuf_4
XTAP_4660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput183 la_iena_mprj[30] vssd vssd vccd vccd net183 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output508_A net1119 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput194 la_iena_mprj[40] vssd vssd vccd vccd net194 sky130_fd_sc_hd__clkbuf_4
XTAP_4671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1041_A net741 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1139_A net557 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output877_A net1277 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__491__B net2082 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1675_A mprj_logic1\[80\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput602 net602 vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_8
XFILLER_9_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput613 net613 vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_8
Xoutput624 net624 vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_8
XFILLER_29_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput635 net635 vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_8
Xoutput646 net646 vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_8
Xoutput657 net657 vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_8
XANTENNA_wire1842_A mprj_logic1\[34\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput668 net668 vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_8
XFILLER_47_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput679 net679 vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_8
XFILLER_29_2794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1900 net1901 vssd vssd vccd vccd net1900 sky130_fd_sc_hd__buf_6
XFILLER_28_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input141_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1911 net1912 vssd vssd vccd vccd net1911 sky130_fd_sc_hd__buf_6
XFILLER_3_4390 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1922 net1923 vssd vssd vccd vccd net1922 sky130_fd_sc_hd__buf_6
XANTENNA_wire2156_A net2157 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input239_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1933 mprj_logic1\[311\] vssd vssd vccd vccd net1933 sky130_fd_sc_hd__buf_6
XANTENNA__421__A_N net335 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1944 mprj_logic1\[306\] vssd vssd vccd vccd net1944 sky130_fd_sc_hd__buf_6
XTAP_3200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1955 net1956 vssd vssd vccd vccd net1955 sky130_fd_sc_hd__buf_6
XTAP_3211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1966 mprj_logic1\[298\] vssd vssd vccd vccd net1966 sky130_fd_sc_hd__buf_6
XFILLER_19_4321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1977 net1978 vssd vssd vccd vccd net1977 sky130_fd_sc_hd__buf_6
XTAP_3233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1988 net1989 vssd vssd vccd vccd net1988 sky130_fd_sc_hd__buf_6
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1999 net2000 vssd vssd vccd vccd net1999 sky130_fd_sc_hd__buf_6
XANTENNA__576__B net1996 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input406_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_200 net1837 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 net1988 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 net2137 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_503_ net354 net2053 vssd vssd vccd vccd net813 sky130_fd_sc_hd__and2_4
XTAP_2532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 net384 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 net1888 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 mprj_logic1\[78\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_434_ net1552 net2196 net1339 vssd vssd vccd vccd net552 sky130_fd_sc_hd__and3b_4
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__592__A net382 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ net1696 net1363 vssd vssd vccd vccd net933 sky130_fd_sc_hd__and2_2
XFILLER_9_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_296_ mprj_logic1\[1\] net1 vssd vssd vccd vccd net955 sky130_fd_sc_hd__and2_4
XFILLER_13_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1089_A net540 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[40\]_B la_data_in_enable\[40\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_29_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1256_A net860 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__486__B net2097 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1423_A net1424 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1792_A mprj_logic1\[429\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__007__A la_data_in_mprj_bar\[24\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] la_data_in_enable\[1\] vssd vssd vccd
+ vccd la_data_in_mprj_bar\[1\] sky130_fd_sc_hd__nand2_1
Xoutput465 net1065 vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__buf_8
XFILLER_5_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_B la_data_in_enable\[31\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xoutput476 net1055 vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__buf_8
XFILLER_44_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__444__A_N net1542 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput487 net487 vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__buf_8
XFILLER_9_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput498 net1128 vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__buf_8
XFILLER_25_3178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1207 net920 vssd vssd vccd vccd net1207 sky130_fd_sc_hd__buf_6
Xwire1218 net1219 vssd vssd vccd vccd net1218 sky130_fd_sc_hd__buf_6
XFILLER_47_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1229 net1230 vssd vssd vccd vccd net1229 sky130_fd_sc_hd__buf_6
XFILLER_9_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__396__B mprj_logic1\[101\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_B la_data_in_enable\[98\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_150_ la_data_in_mprj_bar\[3\] vssd vssd vccd vccd net652 sky130_fd_sc_hd__inv_2
XFILLER_36_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_081_ la_data_in_mprj_bar\[98\] vssd vssd vccd vccd net716 sky130_fd_sc_hd__clkinv_4
XFILLER_12_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input189_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input356_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_B la_data_in_enable\[22\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_43_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__587__A net377 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1730 net1731 vssd vssd vccd vccd net1730 sky130_fd_sc_hd__buf_6
Xwire1741 mprj_logic1\[455\] vssd vssd vccd vccd net1741 sky130_fd_sc_hd__buf_6
Xwire1752 mprj_logic1\[450\] vssd vssd vccd vccd net1752 sky130_fd_sc_hd__buf_6
Xwire1763 net1764 vssd vssd vccd vccd net1763 sky130_fd_sc_hd__buf_6
XFILLER_1_2936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1774 mprj_logic1\[439\] vssd vssd vccd vccd net1774 sky130_fd_sc_hd__buf_6
XTAP_3030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1785 net1786 vssd vssd vccd vccd net1785 sky130_fd_sc_hd__buf_6
XTAP_3041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1796 mprj_logic1\[427\] vssd vssd vccd vccd net1796 sky130_fd_sc_hd__buf_6
XTAP_3052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[89\]_B net1325 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_417_ net330 mprj_logic1\[122\] net74 vssd vssd vccd vccd net533 sky130_fd_sc_hd__and3b_4
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_348_ mprj_logic1\[53\] net1387 vssd vssd vccd vccd net915 sky130_fd_sc_hd__and2_4
XANTENNA_wire1004_A net797 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output575_A net575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_279_ net1759 net150 vssd vssd vccd vccd la_data_in_enable\[116\] sky130_fd_sc_hd__and2_4
XFILLER_13_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__467__A_N net1528 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A net742 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1373_A net1374 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] net1327 vssd vssd vccd vccd la_data_in_mprj_bar\[87\]
+ sky130_fd_sc_hd__nand2_8
XFILLER_22_3318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1540_A net362 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1638_A mprj_logic1\[98\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__497__A net260 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1004 net797 vssd vssd vccd vccd net1004 sky130_fd_sc_hd__buf_6
Xwire1015 net785 vssd vssd vccd vccd net1015 sky130_fd_sc_hd__buf_6
Xwire1026 net765 vssd vssd vccd vccd net1026 sky130_fd_sc_hd__buf_6
XFILLER_2_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1037 net753 vssd vssd vccd vccd net1037 sky130_fd_sc_hd__buf_6
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1048 net802 vssd vssd vccd vccd net1048 sky130_fd_sc_hd__buf_6
XANTENNA__200__A mprj_logic1\[367\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1059 net471 vssd vssd vccd vccd net1059 sky130_fd_sc_hd__buf_6
XFILLER_21_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input104_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2119_A net2120 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_202_ mprj_logic1\[369\] net192 vssd vssd vccd vccd la_data_in_enable\[39\] sky130_fd_sc_hd__and2_4
XFILLER_51_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_133_ mprj_dat_i_core_bar\[19\] vssd vssd vccd vccd net891 sky130_fd_sc_hd__inv_2
XFILLER_10_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_064_ net975 vssd vssd vccd vccd net698 sky130_fd_sc_hd__clkinv_2
XFILLER_10_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__110__A net979 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1560 net33 vssd vssd vccd vccd net1560 sky130_fd_sc_hd__buf_6
Xwire1571 net312 vssd vssd vccd vccd net1571 sky130_fd_sc_hd__buf_6
Xwire1582 net287 vssd vssd vccd vccd net1582 sky130_fd_sc_hd__buf_6
XFILLER_19_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1593 net275 vssd vssd vccd vccd net1593 sky130_fd_sc_hd__buf_8
XFILLER_1_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1121_A net506 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output692_A net692 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1219_A net916 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__C net20 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] net1311 vssd vssd vccd vccd mprj_dat_i_core_bar\[15\]
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1490_A net1491 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1755_A net1756 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1922_A net1923 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__020__A la_data_in_mprj_bar\[37\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] la_data_in_enable\[113\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[113\] sky130_fd_sc_hd__nand2_2
XFILLER_6_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__393__C net48 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2069_A net2070 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input221_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input319_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__584__B net1979 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_116_ mprj_dat_i_core_bar\[2\] vssd vssd vccd vccd net903 sky130_fd_sc_hd__clkinv_2
XFILLER_51_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__105__A net982 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_047_ la_data_in_mprj_bar\[64\] vssd vssd vccd vccd net679 sky130_fd_sc_hd__clkinv_2
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output538_A net1091 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1071_A net585 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2080 net2081 vssd vssd vccd vccd net2080 sky130_fd_sc_hd__buf_6
XFILLER_43_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2091 net2092 vssd vssd vccd vccd net2091 sky130_fd_sc_hd__buf_6
XFILLER_21_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1336_A net96 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1390 net422 vssd vssd vccd vccd net1390 sky130_fd_sc_hd__buf_6
XFILLER_36_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__494__B net2073 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_B la_data_in_enable\[119\] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1503_A net1504 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1872_A net1873 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__388__C net42 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmax_length1310 wb_in_enable vssd vssd vccd vccd net1310 sky130_fd_sc_hd__buf_8
XFILLER_29_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input171_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input269_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2186_A net2187 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__579__B net1990 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input436_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[19\]_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput310 la_oenb_mprj[2] vssd vssd vccd vccd net310 sky130_fd_sc_hd__buf_4
XFILLER_22_4180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput321 la_oenb_mprj[3] vssd vssd vccd vccd net321 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input32_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput332 la_oenb_mprj[4] vssd vssd vccd vccd net332 sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput343 la_oenb_mprj[5] vssd vssd vccd vccd net343 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput354 la_oenb_mprj[6] vssd vssd vccd vccd net354 sky130_fd_sc_hd__clkbuf_4
Xinput365 la_oenb_mprj[7] vssd vssd vccd vccd net365 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput376 la_oenb_mprj[8] vssd vssd vccd vccd net376 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput387 la_oenb_mprj[9] vssd vssd vccd vccd net387 sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput398 mprj_adr_o_core[19] vssd vssd vccd vccd net398 sky130_fd_sc_hd__buf_6
XANTENNA__595__A net1528 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_596_ net1527 net1955 vssd vssd vccd vccd net845 sky130_fd_sc_hd__and2_4
XFILLER_32_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output488_A net488 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output655_A net655 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_3 la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput806 net806 vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__buf_8
Xoutput817 net817 vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__buf_8
XFILLER_6_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput828 net828 vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__buf_8
XFILLER_29_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1286_A net1287 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput839 net839 vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__buf_8
XFILLER_42_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output822_A net822 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__B net2088 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1453_A net1454 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1620_A net114 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__399__B mprj_logic1\[104\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ net1536 net2167 net1623 vssd vssd vccd vccd net570 sky130_fd_sc_hd__and3b_4
XTAP_2747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_381_ net291 net1661 net35 vssd vssd vccd vccd net494 sky130_fd_sc_hd__and3b_4
XFILLER_40_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2101_A mprj_logic1\[190\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input386_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput140 la_iena_mprj[107] vssd vssd vccd vccd net140 sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput151 la_iena_mprj[117] vssd vssd vccd vccd net151 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput162 la_iena_mprj[127] vssd vssd vccd vccd net162 sky130_fd_sc_hd__clkbuf_4
Xinput173 la_iena_mprj[21] vssd vssd vccd vccd net173 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput184 la_iena_mprj[31] vssd vssd vccd vccd net184 sky130_fd_sc_hd__clkbuf_4
XTAP_4661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 la_iena_mprj[41] vssd vssd vccd vccd net195 sky130_fd_sc_hd__clkbuf_4
XTAP_4672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_579_ net1535 net1990 vssd vssd vccd vccd net827 sky130_fd_sc_hd__and2_4
XFILLER_53_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output772_A net772 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__491__C net29 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput603 net603 vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_8
Xoutput614 net614 vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_8
XANTENNA_wire1668_A net1669 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput625 net625 vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_8
XFILLER_25_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput636 net636 vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_8
XFILLER_29_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput647 net647 vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_8
XFILLER_42_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput658 net658 vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_8
XFILLER_45_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput669 net669 vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_8
XFILLER_28_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1835_A net1836 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__373__A_N net332 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__203__A mprj_logic1\[370\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1901 mprj_logic1\[321\] vssd vssd vccd vccd net1901 sky130_fd_sc_hd__buf_6
XFILLER_41_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1912 net1913 vssd vssd vccd vccd net1912 sky130_fd_sc_hd__buf_6
Xwire1923 net1924 vssd vssd vccd vccd net1923 sky130_fd_sc_hd__buf_6
Xwire1934 net1935 vssd vssd vccd vccd net1934 sky130_fd_sc_hd__buf_6
Xwire1945 net1946 vssd vssd vccd vccd net1945 sky130_fd_sc_hd__buf_6
XFILLER_19_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input134_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1956 mprj_logic1\[301\] vssd vssd vccd vccd net1956 sky130_fd_sc_hd__buf_6
XANTENNA_wire2051_A mprj_logic1\[210\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1967 net1968 vssd vssd vccd vccd net1967 sky130_fd_sc_hd__buf_6
XANTENNA_wire2149_A net2150 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1978 mprj_logic1\[290\] vssd vssd vccd vccd net1978 sky130_fd_sc_hd__buf_6
XTAP_3234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1989 mprj_logic1\[285\] vssd vssd vccd vccd net1989 sky130_fd_sc_hd__buf_6
XFILLER_18_438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 net1865 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ net343 net2055 vssd vssd vccd vccd net802 sky130_fd_sc_hd__and2_4
XANTENNA_212 net2009 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input301_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_223 mprj_logic1\[142\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 net1354 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_245 net1984 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 net1575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_433_ net1553 net2197 net92 vssd vssd vccd vccd net551 sky130_fd_sc_hd__and3b_4
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__592__B net1967 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_364_ net1700 net1364 vssd vssd vccd vccd net932 sky130_fd_sc_hd__and2_2
XFILLER_35_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_295_ net1576 net2203 vssd vssd vccd vccd net960 sky130_fd_sc_hd__and2b_2
XFILLER_9_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output520_A net1108 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output618_A net618 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1151_A net1152 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1249_A net1250 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__486__C net23 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__396__A_N net1575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1416_A net415 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] la_data_in_enable\[32\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[32\] sky130_fd_sc_hd__nand2_4
XFILLER_18_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1785_A net1786 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__023__A la_data_in_mprj_bar\[40\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput466 net1064 vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__buf_8
XFILLER_25_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput477 net1054 vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__buf_8
XFILLER_47_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput488 net488 vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__buf_8
Xoutput499 net1127 vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__buf_8
XFILLER_47_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1208 net1209 vssd vssd vccd vccd net1208 sky130_fd_sc_hd__buf_6
XFILLER_5_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1219 net916 vssd vssd vccd vccd net1219 sky130_fd_sc_hd__buf_6
XFILLER_45_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__396__C net51 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3426 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_080_ la_data_in_mprj_bar\[97\] vssd vssd vccd vccd net715 sky130_fd_sc_hd__clkinv_4
XFILLER_17_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2099_A net2100 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input251_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input349_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1720 net1721 vssd vssd vccd vccd net1720 sky130_fd_sc_hd__buf_6
XANTENNA__587__B net1975 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1731 mprj_logic1\[459\] vssd vssd vccd vccd net1731 sky130_fd_sc_hd__buf_6
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1742 net1743 vssd vssd vccd vccd net1742 sky130_fd_sc_hd__buf_6
Xwire1753 net1754 vssd vssd vccd vccd net1753 sky130_fd_sc_hd__buf_6
Xwire1764 mprj_logic1\[444\] vssd vssd vccd vccd net1764 sky130_fd_sc_hd__buf_6
XFILLER_46_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1775 net1776 vssd vssd vccd vccd net1775 sky130_fd_sc_hd__buf_6
XTAP_3031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1786 mprj_logic1\[432\] vssd vssd vccd vccd net1786 sky130_fd_sc_hd__buf_6
XFILLER_37_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1797 mprj_logic1\[426\] vssd vssd vccd vccd net1797 sky130_fd_sc_hd__buf_6
XTAP_3053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_416_ net329 mprj_logic1\[121\] net73 vssd vssd vccd vccd net532 sky130_fd_sc_hd__and3b_4
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__108__A la_data_in_mprj_bar\[125\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_347_ mprj_logic1\[52\] net1389 vssd vssd vccd vccd net914 sky130_fd_sc_hd__and2_4
X_278_ net1761 net149 vssd vssd vccd vccd la_data_in_enable\[115\] sky130_fd_sc_hd__and2_4
XANTENNA_output470_A net1060 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output568_A net1138 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1199_A net1200 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output735_A net735 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1366_A net438 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__497__B net2064 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1533_A net370 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1700_A net1701 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire986_A la_data_in_mprj_bar\[113\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__411__A_N net324 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1005 net1006 vssd vssd vccd vccd net1005 sky130_fd_sc_hd__buf_6
XFILLER_40_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1016 net1017 vssd vssd vccd vccd net1016 sky130_fd_sc_hd__buf_6
XFILLER_25_2286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1027 net764 vssd vssd vccd vccd net1027 sky130_fd_sc_hd__buf_6
Xwire1038 net752 vssd vssd vccd vccd net1038 sky130_fd_sc_hd__buf_6
Xwire1049 net791 vssd vssd vccd vccd net1049 sky130_fd_sc_hd__buf_6
XFILLER_0_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2014_A mprj_logic1\[272\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_201_ mprj_logic1\[368\] net191 vssd vssd vccd vccd la_data_in_enable\[38\] sky130_fd_sc_hd__and2_4
XFILLER_11_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input299_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_132_ mprj_dat_i_core_bar\[18\] vssd vssd vccd vccd net890 sky130_fd_sc_hd__inv_2
XFILLER_8_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_063_ net976 vssd vssd vccd vccd net697 sky130_fd_sc_hd__clkinv_2
XFILLER_10_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input62_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__598__A net1606 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1550 net351 vssd vssd vccd vccd net1550 sky130_fd_sc_hd__buf_6
XFILLER_19_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1561 net1562 vssd vssd vccd vccd net1561 sky130_fd_sc_hd__buf_6
XFILLER_21_2662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1572 net311 vssd vssd vccd vccd net1572 sky130_fd_sc_hd__buf_8
Xwire1583 net286 vssd vssd vccd vccd net1583 sky130_fd_sc_hd__buf_6
XFILLER_19_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1594 net274 vssd vssd vccd vccd net1594 sky130_fd_sc_hd__buf_6
XFILLER_1_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__434__A_N net1552 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output852_A net1264 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1483_A net1484 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1650_A net1651 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__301__A net1698 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1915_A net1916 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] la_data_in_enable\[106\] vssd
+ vssd vccd vccd la_data_in_mprj_bar\[106\] sky130_fd_sc_hd__nand2_8
XFILLER_0_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__211__A mprj_logic1\[378\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input214_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__457__A_N net1529 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_115_ mprj_dat_i_core_bar\[1\] vssd vssd vccd vccd net892 sky130_fd_sc_hd__clkinv_2
XFILLER_45_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_046_ la_data_in_mprj_bar\[63\] vssd vssd vccd vccd net678 sky130_fd_sc_hd__clkinv_2
XFILLER_45_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__121__A mprj_dat_i_core_bar\[7\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1064_A net466 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2070 net2071 vssd vssd vccd vccd net2070 sky130_fd_sc_hd__buf_6
Xwire2081 mprj_logic1\[197\] vssd vssd vccd vccd net2081 sky130_fd_sc_hd__buf_6
XFILLER_36_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output600_A net600 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2092 net2093 vssd vssd vccd vccd net2092 sky130_fd_sc_hd__buf_6
XFILLER_43_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1380 net427 vssd vssd vccd vccd net1380 sky130_fd_sc_hd__buf_6
XFILLER_19_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1391 net1392 vssd vssd vccd vccd net1391 sky130_fd_sc_hd__buf_6
XANTENNA_wire1231_A net943 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1329_A la_data_in_enable\[85\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__494__C net1566 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1698_A net1699 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3896 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1865_A net1866 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_B net1310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__A net1820 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xmax_length1311 wb_in_enable vssd vssd vccd vccd net1311 sky130_fd_sc_hd__buf_8
XFILLER_11_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2081_A mprj_logic1\[197\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input164_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2179_A mprj_logic1\[14\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput300 la_oenb_mprj[20] vssd vssd vccd vccd net300 sky130_fd_sc_hd__buf_4
XFILLER_1_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[19\]_B net1311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput311 la_oenb_mprj[30] vssd vssd vccd vccd net311 sky130_fd_sc_hd__buf_6
Xinput322 la_oenb_mprj[40] vssd vssd vccd vccd net322 sky130_fd_sc_hd__buf_6
XFILLER_22_4192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput333 la_oenb_mprj[50] vssd vssd vccd vccd net333 sky130_fd_sc_hd__buf_4
XANTENNA_input331_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput344 la_oenb_mprj[60] vssd vssd vccd vccd net344 sky130_fd_sc_hd__buf_4
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input429_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput355 la_oenb_mprj[70] vssd vssd vccd vccd net355 sky130_fd_sc_hd__buf_6
XFILLER_2_4297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput366 la_oenb_mprj[80] vssd vssd vccd vccd net366 sky130_fd_sc_hd__buf_6
XANTENNA_input25_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput377 la_oenb_mprj[90] vssd vssd vccd vccd net377 sky130_fd_sc_hd__buf_4
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput388 mprj_adr_o_core[0] vssd vssd vccd vccd net388 sky130_fd_sc_hd__buf_6
Xinput399 mprj_adr_o_core[1] vssd vssd vccd vccd net399 sky130_fd_sc_hd__buf_6
XFILLER_18_4217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__595__B net1957 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_595_ net1528 net1957 vssd vssd vccd vccd net844 sky130_fd_sc_hd__and2_4
XFILLER_31_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_4 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput807 net807 vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__buf_8
Xoutput818 net818 vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__buf_8
XFILLER_49_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output550_A net550 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput829 net829 vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__buf_8
XFILLER_6_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_029_ la_data_in_mprj_bar\[46\] vssd vssd vccd vccd net659 sky130_fd_sc_hd__inv_2
XFILLER_42_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1279_A net876 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__C net1598 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output815_A net815 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1446_A net409 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] la_data_in_enable\[62\] vssd vssd
+ vccd vccd la_data_in_mprj_bar\[62\] sky130_fd_sc_hd__nand2_4
XFILLER_39_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1982_A net1983 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__026__A la_data_in_mprj_bar\[43\] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__399__C net55 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_380_ net282 net1663 net26 vssd vssd vccd vccd net485 sky130_fd_sc_hd__and3b_1
XFILLER_13_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input281_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input379_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput130 la_data_out_mprj[99] vssd vssd vccd vccd net130 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput141 la_iena_mprj[108] vssd vssd vccd vccd net141 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput152 la_iena_mprj[118] vssd vssd vccd vccd net152 sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput163 la_iena_mprj[12] vssd vssd vccd vccd net163 sky130_fd_sc_hd__clkbuf_4
XTAP_4640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 la_iena_mprj[22] vssd vssd vccd vccd net174 sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput185 la_iena_mprj[32] vssd vssd vccd vccd net185 sky130_fd_sc_hd__clkbuf_4
XTAP_4662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput196 la_iena_mprj[42] vssd vssd vccd vccd net196 sky130_fd_sc_hd__buf_4
XTAP_4673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_578_ net1536 net1992 vssd vssd vccd vccd net826 sky130_fd_sc_hd__and2_4
XFILLER_16_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output598_A net598 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output765_A net1026 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1396_A net1397 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output932_A net1162 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput604 net604 vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput615 net615 vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_8
XFILLER_44_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput626 net626 vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_8
Xoutput637 net637 vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_8
XANTENNA_wire1563_A net328 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput648 net648 vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_8
XFILLER_28_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput659 net659 vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_8
XFILLER_42_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1730_A net1731 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
.ends

