* NGSPICE file created from constant_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_4 abstract view
.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_16 abstract view
.subckt sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_8 abstract view
.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

.subckt constant_block one vccd vssd zero
XFILLER_0_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_0 vssd vssd vccd vccd sky130_fd_sc_hd__fill_4
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xconst_zero_buf const_source/LO vssd vssd vccd vccd zero sky130_fd_sc_hd__buf_16
XFILLER_1_4 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xconst_source vssd vssd vccd vccd const_source/HI const_source/LO sky130_fd_sc_hd__conb_1
XFILLER_1_8 vssd vssd vccd vccd sky130_fd_sc_hd__fill_8
XFILLER_1_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_4
XFILLER_1_16 vssd vssd vccd vccd sky130_fd_sc_hd__fill_8
Xconst_one_buf const_source/HI vssd vssd vccd vccd one sky130_fd_sc_hd__buf_16
XTAP_0 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_0 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_0 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
.ends

