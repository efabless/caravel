module caravel_power_routing ();
endmodule
