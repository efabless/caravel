* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_8 abstract view
.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt digital_pll VGND VPWR clockp[0] clockp[1] dco div[0] div[1] div[2] div[3]
+ div[4] enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__338__A1 ext_trim[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_294_ _297_/C _302_/C _301_/A VGND VGND VPWR VPWR _294_/X sky130_fd_sc_hd__or3_2
X_363_ _328_/A _363_/D _318_/X VGND VGND VPWR VPWR _363_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_346_ _288_/B ext_trim[3] dco VGND VGND VPWR VPWR _346_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_277_ _362_/Q _272_/B _363_/Q _267_/B _226_/B VGND VGND VPWR VPWR _359_/D sky130_fd_sc_hd__a311o_2
X_200_ _196_/A _199_/Y _196_/A _199_/Y VGND VGND VPWR VPWR _200_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _331_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_329_ _292_/B _232_/B _370_/Q VGND VGND VPWR VPWR _329_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _332_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _334_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_362_ _328_/A _362_/D _319_/X VGND VGND VPWR VPWR _362_/Q sky130_fd_sc_hd__dfrtp_2
X_293_ _367_/Q _221_/B _302_/B _370_/Q _232_/B VGND VGND VPWR VPWR _293_/X sky130_fd_sc_hd__o311a_2
X_276_ _276_/A _276_/B VGND VGND VPWR VPWR _360_/D sky130_fd_sc_hd__or2_2
X_345_ _300_/X ext_trim[17] dco VGND VGND VPWR VPWR _345_/X sky130_fd_sc_hd__mux2_1
X_328_ _328_/A VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__buf_2
X_259_ _366_/Q _220_/Y _262_/A VGND VGND VPWR VPWR _259_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _333_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _335_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_361_ _328_/A _361_/D _320_/X VGND VGND VPWR VPWR _361_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_292_ _301_/A _292_/B VGND VGND VPWR VPWR _299_/B sky130_fd_sc_hd__nand2_2
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_344_ _286_/X ext_trim[4] dco VGND VGND VPWR VPWR _344_/X sky130_fd_sc_hd__mux2_1
X_275_ _267_/A _267_/B _360_/Q _359_/Q _272_/D VGND VGND VPWR VPWR _276_/B sky130_fd_sc_hd__o221a_2
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _344_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_327_ _327_/A VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__buf_1
X_258_ _262_/A _262_/B VGND VGND VPWR VPWR _258_/X sky130_fd_sc_hd__or2_2
X_189_ _371_/Q _226_/B VGND VGND VPWR VPWR _371_/D sky130_fd_sc_hd__or2_2
XANTENNA__210__B1 div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _342_/X VGND
+ VGND VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvn_8
XANTENNA__201__B1 div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_360_ _328_/A _360_/D _321_/X VGND VGND VPWR VPWR _360_/Q sky130_fd_sc_hd__dfrtp_2
X_291_ _369_/Q _368_/Q _367_/Q _370_/Q VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__a31o_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_274_ _272_/D _268_/A _273_/Y _276_/A VGND VGND VPWR VPWR _361_/D sky130_fd_sc_hd__a31o_2
X_343_ _301_/Y ext_trim[18] dco VGND VGND VPWR VPWR _343_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _345_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_326_ _370_/Q VGND VGND VPWR VPWR _326_/X sky130_fd_sc_hd__buf_1
X_257_ _236_/A _251_/X _256_/Y _368_/Q _236_/Y VGND VGND VPWR VPWR _368_/D sky130_fd_sc_hd__a32o_2
X_188_ _372_/Q _272_/D _371_/Q _226_/B VGND VGND VPWR VPWR _372_/D sky130_fd_sc_hd__a22o_2
X_309_ _327_/A VGND VGND VPWR VPWR _309_/X sky130_fd_sc_hd__buf_1
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__210__A1 div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _343_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XANTENNA__201__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_290_ _369_/Q _368_/Q _297_/C _370_/Q VGND VGND VPWR VPWR _290_/X sky130_fd_sc_hd__a31o_2
X_342_ _283_/X ext_trim[5] dco VGND VGND VPWR VPWR _342_/X sky130_fd_sc_hd__mux2_1
X_273_ _267_/A _267_/B _267_/C VGND VGND VPWR VPWR _273_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ _327_/A VGND VGND VPWR VPWR _325_/X sky130_fd_sc_hd__buf_1
X_256_ _256_/A _256_/B VGND VGND VPWR VPWR _256_/Y sky130_fd_sc_hd__nand2_2
X_187_ _372_/Q _226_/B _373_/Q _272_/D VGND VGND VPWR VPWR _373_/D sky130_fd_sc_hd__a22o_2
X_308_ _327_/A VGND VGND VPWR VPWR _308_/X sky130_fd_sc_hd__buf_1
X_239_ _288_/A _239_/B VGND VGND VPWR VPWR _239_/Y sky130_fd_sc_hd__nor2_2
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_272_ _362_/Q _272_/B _363_/Q _272_/D VGND VGND VPWR VPWR _276_/A sky130_fd_sc_hd__and4_2
X_341_ _299_/B ext_trim[19] dco VGND VGND VPWR VPWR _341_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _350_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XANTENNA__340__A1 ext_trim[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XANTENNA__181__A enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__331__A1 ext_trim[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_186_ _374_/Q _272_/D _359_/Q _226_/B VGND VGND VPWR VPWR _374_/D sky130_fd_sc_hd__a22o_2
X_324_ _327_/A VGND VGND VPWR VPWR _324_/X sky130_fd_sc_hd__buf_1
X_255_ _297_/A _236_/A _254_/X VGND VGND VPWR VPWR _369_/D sky130_fd_sc_hd__o21ai_2
X_169_ _374_/Q VGND VGND VPWR VPWR _193_/B sky130_fd_sc_hd__inv_2
X_307_ _327_/A VGND VGND VPWR VPWR _307_/X sky130_fd_sc_hd__buf_1
X_238_ _224_/A _220_/A _224_/B _237_/X VGND VGND VPWR VPWR _262_/A sky130_fd_sc_hd__o22a_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _351_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_340_ _279_/X ext_trim[6] dco VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__mux2_1
X_271_ _362_/Q _272_/B _363_/Q _269_/Y _272_/D VGND VGND VPWR VPWR _362_/D sky130_fd_sc_hd__o221a_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__181__B resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _350_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_185_ _375_/Q _272_/D _360_/Q _226_/B VGND VGND VPWR VPWR _375_/D sky130_fd_sc_hd__a22o_2
X_323_ _327_/A VGND VGND VPWR VPWR _323_/X sky130_fd_sc_hd__buf_1
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_254_ _244_/Y _253_/A _244_/A _253_/Y _236_/Y VGND VGND VPWR VPWR _254_/X sky130_fd_sc_hd__a221o_2
X_306_ _327_/A VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__buf_1
X_168_ _359_/Q VGND VGND VPWR VPWR _267_/B sky130_fd_sc_hd__inv_2
X_237_ _365_/Q _220_/Y _224_/A _220_/A VGND VGND VPWR VPWR _237_/X sky130_fd_sc_hd__a22o_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__204__A1 div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_270_ _164_/Y _269_/Y _226_/B VGND VGND VPWR VPWR _363_/D sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _351_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_322_ _327_/A VGND VGND VPWR VPWR _322_/X sky130_fd_sc_hd__buf_1
XFILLER_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_184_ _376_/Q _272_/D _361_/Q _226_/B VGND VGND VPWR VPWR _376_/D sky130_fd_sc_hd__a22o_2
X_253_ _253_/A VGND VGND VPWR VPWR _253_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ _327_/A VGND VGND VPWR VPWR _305_/X sky130_fd_sc_hd__buf_1
X_167_ _360_/Q VGND VGND VPWR VPWR _267_/A sky130_fd_sc_hd__inv_2
X_236_ _236_/A VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _219_/A _219_/B VGND VGND VPWR VPWR _220_/A sky130_fd_sc_hd__or2_2
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _334_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__330__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__343__A1 ext_trim[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__352__A1 ext_trim[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__334__A1 ext_trim[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__356__D osc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_321_ _327_/A VGND VGND VPWR VPWR _321_/X sky130_fd_sc_hd__buf_1
X_183_ _377_/Q _272_/D _362_/Q _226_/B VGND VGND VPWR VPWR _377_/D sky130_fd_sc_hd__a22o_2
X_252_ _280_/B _220_/A _251_/X VGND VGND VPWR VPWR _253_/A sky130_fd_sc_hd__o21ai_2
X_304_ _288_/A _239_/B _302_/B _370_/Q _232_/B VGND VGND VPWR VPWR _304_/X sky130_fd_sc_hd__o311a_2
X_235_ _301_/A _220_/Y _224_/X _234_/X VGND VGND VPWR VPWR _236_/A sky130_fd_sc_hd__o31a_2
X_166_ _361_/Q VGND VGND VPWR VPWR _267_/C sky130_fd_sc_hd__inv_2
XANTENNA__333__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_218_ _164_/Y _165_/Y div[4] _216_/B _214_/X VGND VGND VPWR VPWR _219_/B sky130_fd_sc_hd__o221ai_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _335_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__341__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_320_ _327_/A VGND VGND VPWR VPWR _320_/X sky130_fd_sc_hd__buf_1
X_182_ dco _182_/B VGND VGND VPWR VPWR _327_/A sky130_fd_sc_hd__nor2_2
X_251_ _256_/A _256_/B VGND VGND VPWR VPWR _251_/X sky130_fd_sc_hd__or2_2
XANTENNA__336__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_165_ _378_/Q VGND VGND VPWR VPWR _165_/Y sky130_fd_sc_hd__inv_2
X_303_ _297_/A _368_/Q _367_/Q _302_/X VGND VGND VPWR VPWR _303_/X sky130_fd_sc_hd__o31a_2
X_234_ _219_/B _225_/Y _220_/A _233_/X _226_/X VGND VGND VPWR VPWR _234_/X sky130_fd_sc_hd__o221a_2
Xringosc.iss.reseten0 ringosc.iss.const1/HI _182_/B VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_1
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_217_ _201_/Y _203_/Y _205_/Y _211_/Y _216_/Y VGND VGND VPWR VPWR _219_/A sky130_fd_sc_hd__o221a_2
XANTENNA__344__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__339__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _336_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_181_ enable resetb VGND VGND VPWR VPWR _182_/B sky130_fd_sc_hd__nand2_2
X_250_ _301_/A _236_/A _249_/X VGND VGND VPWR VPWR _370_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__352__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_164_ _363_/Q VGND VGND VPWR VPWR _164_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_302_ _370_/Q _302_/B _302_/C VGND VGND VPWR VPWR _302_/X sky130_fd_sc_hd__and3_2
X_233_ _365_/Q _364_/Q _233_/C VGND VGND VPWR VPWR _233_/X sky130_fd_sc_hd__or3_2
XANTENNA__347__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_216_ div[4] _216_/B VGND VGND VPWR VPWR _216_/Y sky130_fd_sc_hd__nand2_2
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XANTENNA__355__A1 ext_trim[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__346__A1 ext_trim[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__337__A1 ext_trim[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__355__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _337_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_180_ _378_/Q _272_/D _363_/Q _226_/B VGND VGND VPWR VPWR _378_/D sky130_fd_sc_hd__a22o_2
X_378_ _328_/A _378_/D _327_/X VGND VGND VPWR VPWR _378_/Q sky130_fd_sc_hd__dfrtp_2
X_232_ _370_/Q _232_/B VGND VGND VPWR VPWR _233_/C sky130_fd_sc_hd__or2_2
X_301_ _301_/A _301_/B VGND VGND VPWR VPWR _301_/Y sky130_fd_sc_hd__nor2_2
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _340_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_215_ _214_/A _214_/B _214_/X VGND VGND VPWR VPWR _216_/B sky130_fd_sc_hd__a21bo_2
XANTENNA__207__A div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_377_ _328_/A _377_/D _327_/A VGND VGND VPWR VPWR _377_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _344_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_300_ _221_/A _366_/Q _301_/A _302_/C _296_/X VGND VGND VPWR VPWR _300_/X sky130_fd_sc_hd__o41a_2
X_231_ _297_/C _302_/B VGND VGND VPWR VPWR _232_/B sky130_fd_sc_hd__or2_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _332_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _341_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_214_ _214_/A _214_/B VGND VGND VPWR VPWR _214_/X sky130_fd_sc_hd__or2_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_376_ _328_/A _376_/D _305_/X VGND VGND VPWR VPWR _376_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _345_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_230_ _302_/B VGND VGND VPWR VPWR _301_/B sky130_fd_sc_hd__inv_2
X_359_ _328_/A _359_/D _322_/X VGND VGND VPWR VPWR _359_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _333_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_213_ _362_/Q _377_/Q _190_/Y _197_/X VGND VGND VPWR VPWR _214_/B sky130_fd_sc_hd__o2bb2a_2
XANTENNA__349__A1 ext_trim[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_375_ _328_/A _375_/D _306_/X VGND VGND VPWR VPWR _375_/Q sky130_fd_sc_hd__dfrtp_2
X_358_ _328_/A _358_/D _323_/X VGND VGND VPWR VPWR _358_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ _297_/A _368_/Q _370_/Q _284_/X VGND VGND VPWR VPWR _289_/X sky130_fd_sc_hd__o31a_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_212_ _363_/Q _378_/Q _164_/Y _165_/Y VGND VGND VPWR VPWR _214_/A sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _352_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_374_ _328_/A _374_/D _307_/X VGND VGND VPWR VPWR _374_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _346_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _328_/A _357_/D _324_/X VGND VGND VPWR VPWR _358_/D sky130_fd_sc_hd__dfrtp_2
X_288_ _288_/A _288_/B VGND VGND VPWR VPWR _288_/X sky130_fd_sc_hd__or2_2
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_211_ div[1] _207_/B _210_/X VGND VGND VPWR VPWR _211_/Y sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _353_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VGND VPWR
+ VPWR ringosc.ibufp00/A sky130_fd_sc_hd__einvn_8
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__330__A1 ext_trim[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_373_ _328_/A _373_/D _308_/X VGND VGND VPWR VPWR _373_/Q sky130_fd_sc_hd__dfrtp_2
X_356_ _328_/A osc _325_/X VGND VGND VPWR VPWR _357_/D sky130_fd_sc_hd__dfrtp_2
X_287_ _297_/A _368_/Q _370_/Q _288_/A _284_/X VGND VGND VPWR VPWR _287_/X sky130_fd_sc_hd__o41a_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _347_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ div[1] _207_/B div[0] _209_/Y _207_/Y VGND VGND VPWR VPWR _210_/X sky130_fd_sc_hd__o221a_2
X_339_ _303_/X ext_trim[20] dco VGND VGND VPWR VPWR _339_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _355_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_372_ _328_/A _372_/D _309_/X VGND VGND VPWR VPWR _372_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__182__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_355_ _304_/X ext_trim[25] dco VGND VGND VPWR VPWR _355_/X sky130_fd_sc_hd__mux2_1
X_286_ _297_/A _368_/Q _370_/Q _367_/Q _284_/X VGND VGND VPWR VPWR _286_/X sky130_fd_sc_hd__o41a_2
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__177__A div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ _362_/Q _272_/B VGND VGND VPWR VPWR _269_/Y sky130_fd_sc_hd__nand2_2
X_338_ _290_/X ext_trim[7] dco VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_371_ _328_/A _371_/D _310_/X VGND VGND VPWR VPWR _371_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_354_ _282_/X ext_trim[12] dco VGND VGND VPWR VPWR _354_/X sky130_fd_sc_hd__mux2_1
X_285_ _297_/A _368_/Q _370_/Q _297_/C _284_/X VGND VGND VPWR VPWR _285_/X sky130_fd_sc_hd__o41a_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_199_ _361_/Q _376_/Q _192_/Y VGND VGND VPWR VPWR _199_/Y sky130_fd_sc_hd__a21oi_2
X_268_ _268_/A VGND VGND VPWR VPWR _272_/B sky130_fd_sc_hd__inv_2
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_337_ _293_/X ext_trim[21] dco VGND VGND VPWR VPWR _337_/X sky130_fd_sc_hd__mux2_1
XANTENNA__351__A1 ext_trim[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__342__A1 ext_trim[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__333__A1 ext_trim[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_370_ _328_/A _370_/D _311_/X VGND VGND VPWR VPWR _370_/Q sky130_fd_sc_hd__dfrtp_2
X_353_ _291_/X ext_trim[13] dco VGND VGND VPWR VPWR _353_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _352_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_284_ _370_/Q _302_/C _288_/B VGND VGND VPWR VPWR _284_/X sky130_fd_sc_hd__o21a_2
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_267_ _267_/A _267_/B _267_/C VGND VGND VPWR VPWR _268_/A sky130_fd_sc_hd__or3_2
X_198_ _191_/X _197_/X _191_/X _197_/X VGND VGND VPWR VPWR _202_/B sky130_fd_sc_hd__a2bb2o_2
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _338_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_336_ _281_/X ext_trim[8] dco VGND VGND VPWR VPWR _336_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_319_ _327_/A VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__buf_1
XANTENNA__331__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _353_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _370_/Q _302_/C _288_/A _288_/B VGND VGND VPWR VPWR _283_/X sky130_fd_sc_hd__o31a_2
X_352_ _233_/C ext_trim[0] dco VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__mux2_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_197_ _361_/Q _376_/Q _192_/Y _196_/Y VGND VGND VPWR VPWR _197_/X sky130_fd_sc_hd__o2bb2a_2
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _339_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_266_ _364_/Q _236_/A _224_/B _236_/Y VGND VGND VPWR VPWR _364_/D sky130_fd_sc_hd__o22a_2
X_335_ _296_/X ext_trim[22] dco VGND VGND VPWR VPWR _335_/X sky130_fd_sc_hd__mux2_1
XANTENNA__334__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_249_ _246_/Y _248_/A _246_/A _248_/Y _236_/Y VGND VGND VPWR VPWR _249_/X sky130_fd_sc_hd__a221o_2
X_318_ _327_/A VGND VGND VPWR VPWR _318_/X sky130_fd_sc_hd__buf_1
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _336_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__342__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ _370_/Q _302_/C _367_/Q _288_/B VGND VGND VPWR VPWR _282_/X sky130_fd_sc_hd__o31a_2
XANTENNA__337__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_351_ _298_/X ext_trim[14] dco VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__mux2_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ _285_/X ext_trim[9] dco VGND VGND VPWR VPWR _334_/X sky130_fd_sc_hd__mux2_1
X_196_ _196_/A VGND VGND VPWR VPWR _196_/Y sky130_fd_sc_hd__inv_2
X_265_ _224_/A _236_/A _236_/Y _264_/X VGND VGND VPWR VPWR _365_/D sky130_fd_sc_hd__o22ai_2
XANTENNA__354__A1 ext_trim[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__350__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_248_ _248_/A VGND VGND VPWR VPWR _248_/Y sky130_fd_sc_hd__inv_2
X_317_ _327_/A VGND VGND VPWR VPWR _317_/X sky130_fd_sc_hd__buf_1
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__345__A1 ext_trim[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_179_ _272_/D VGND VGND VPWR VPWR _226_/B sky130_fd_sc_hd__inv_2
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _346_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__336__A1 ext_trim[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XANTENNA__345__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _337_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XANTENNA__218__B1 div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_350_ _289_/X ext_trim[1] dco VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__mux2_1
XANTENNA__353__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_281_ _297_/C _302_/C _370_/Q _288_/B VGND VGND VPWR VPWR _281_/X sky130_fd_sc_hd__o31a_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__202__A div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__348__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ _360_/Q _375_/Q _193_/Y _194_/X VGND VGND VPWR VPWR _196_/A sky130_fd_sc_hd__a22o_2
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_333_ _326_/X ext_trim[23] dco VGND VGND VPWR VPWR _333_/X sky130_fd_sc_hd__mux2_1
X_264_ _224_/B _237_/X _224_/B _237_/X VGND VGND VPWR VPWR _264_/X sky130_fd_sc_hd__a2bb2o_2
X_247_ _370_/Q _220_/Y _301_/A _220_/A VGND VGND VPWR VPWR _248_/A sky130_fd_sc_hd__o22a_2
X_316_ _327_/A VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _347_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_178_ _358_/D _358_/Q _358_/D _358_/Q VGND VGND VPWR VPWR _272_/D sky130_fd_sc_hd__a2bb2o_2
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_280_ _369_/Q _280_/B VGND VGND VPWR VPWR _302_/C sky130_fd_sc_hd__or2_2
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ _360_/Q _375_/Q _360_/Q _375_/Q VGND VGND VPWR VPWR _194_/X sky130_fd_sc_hd__o2bb2a_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _288_/X ext_trim[10] dco VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__mux2_1
X_263_ _236_/A _258_/X _262_/Y _366_/Q _236_/Y VGND VGND VPWR VPWR _366_/D sky130_fd_sc_hd__a32o_2
XFILLER_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_177_ div[0] VGND VGND VPWR VPWR _177_/Y sky130_fd_sc_hd__inv_2
X_315_ _327_/A VGND VGND VPWR VPWR _315_/X sky130_fd_sc_hd__buf_1
X_246_ _246_/A VGND VGND VPWR VPWR _246_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ _369_/Q _368_/Q VGND VGND VPWR VPWR _302_/B sky130_fd_sc_hd__or2_2
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__clkinv_2
XANTENNA__216__A div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ _267_/B _193_/B VGND VGND VPWR VPWR _193_/Y sky130_fd_sc_hd__nor2_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _302_/X ext_trim[24] dco VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__mux2_1
X_262_ _262_/A _262_/B VGND VGND VPWR VPWR _262_/Y sky130_fd_sc_hd__nand2_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__348__A1 ext_trim[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__339__A1 ext_trim[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ _327_/A VGND VGND VPWR VPWR _314_/X sky130_fd_sc_hd__buf_1
X_245_ _256_/B _244_/A _256_/A _220_/A _301_/B VGND VGND VPWR VPWR _246_/A sky130_fd_sc_hd__o32a_2
X_176_ _364_/Q VGND VGND VPWR VPWR _224_/B sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _342_/X VGND VGND
+ VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvp_2
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_228_ _297_/C VGND VGND VPWR VPWR _239_/B sky130_fd_sc_hd__inv_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.ibufp11 ringosc.ibufp11/A VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkinv_8
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_192_ _361_/Q _376_/Q VGND VGND VPWR VPWR _192_/Y sky130_fd_sc_hd__nor2_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _287_/X ext_trim[11] dco VGND VGND VPWR VPWR _330_/X sky130_fd_sc_hd__mux2_1
X_261_ _367_/Q _260_/X _367_/Q _260_/X VGND VGND VPWR VPWR _367_/D sky130_fd_sc_hd__o2bb2a_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_313_ _327_/A VGND VGND VPWR VPWR _313_/X sky130_fd_sc_hd__buf_1
X_175_ _365_/Q VGND VGND VPWR VPWR _224_/A sky130_fd_sc_hd__inv_2
X_244_ _244_/A VGND VGND VPWR VPWR _244_/Y sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _343_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_227_ _367_/Q _366_/Q VGND VGND VPWR VPWR _297_/C sky130_fd_sc_hd__or2_2
XFILLER_8_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _328_/A sky130_fd_sc_hd__clkinv_8
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _221_/B _220_/A _236_/A _259_/X VGND VGND VPWR VPWR _260_/X sky130_fd_sc_hd__o211a_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ _362_/Q _377_/Q _190_/Y VGND VGND VPWR VPWR _191_/X sky130_fd_sc_hd__a21o_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_174_ _366_/Q VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__inv_2
X_243_ _297_/A _220_/Y _369_/Q _220_/A VGND VGND VPWR VPWR _244_/A sky130_fd_sc_hd__o22a_2
X_312_ _327_/A VGND VGND VPWR VPWR _312_/X sky130_fd_sc_hd__buf_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _330_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvn_8
X_226_ _372_/Q _226_/B _373_/Q _371_/Q VGND VGND VPWR VPWR _226_/X sky130_fd_sc_hd__and4_2
X_209_ _209_/A VGND VGND VPWR VPWR _209_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ _362_/Q _377_/Q VGND VGND VPWR VPWR _190_/Y sky130_fd_sc_hd__nor2_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_311_ _327_/A VGND VGND VPWR VPWR _311_/X sky130_fd_sc_hd__buf_1
X_173_ _367_/Q VGND VGND VPWR VPWR _221_/A sky130_fd_sc_hd__inv_2
X_242_ _368_/Q _220_/Y _280_/B _220_/A VGND VGND VPWR VPWR _256_/B sky130_fd_sc_hd__a22o_2
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_225_ _177_/Y _209_/A _210_/X _205_/A _216_/Y VGND VGND VPWR VPWR _225_/Y sky130_fd_sc_hd__o2111ai_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _331_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ _267_/B _193_/B _193_/Y VGND VGND VPWR VPWR _209_/A sky130_fd_sc_hd__a21oi_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__211__A1 div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ _327_/A VGND VGND VPWR VPWR _310_/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _348_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_241_ _239_/Y _262_/B _262_/A _220_/A _239_/B VGND VGND VPWR VPWR _256_/A sky130_fd_sc_hd__o32a_2
X_172_ _368_/Q VGND VGND VPWR VPWR _280_/B sky130_fd_sc_hd__inv_2
X_224_ _224_/A _224_/B _292_/B VGND VGND VPWR VPWR _224_/X sky130_fd_sc_hd__or3_2
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _340_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_207_ div[1] _207_/B VGND VGND VPWR VPWR _207_/Y sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _349_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_240_ _366_/Q _220_/Y _221_/B _220_/A VGND VGND VPWR VPWR _262_/B sky130_fd_sc_hd__a22o_2
X_171_ _369_/Q VGND VGND VPWR VPWR _297_/A sky130_fd_sc_hd__inv_2
X_369_ _328_/A _369_/D _312_/X VGND VGND VPWR VPWR _369_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__350__A1 ext_trim[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_223_ _297_/A _280_/B _223_/C VGND VGND VPWR VPWR _292_/B sky130_fd_sc_hd__or3_2
XANTENNA__341__A1 ext_trim[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__332__A1 ext_trim[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _341_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_206_ _193_/Y _194_/X _193_/Y _194_/X VGND VGND VPWR VPWR _207_/B sky130_fd_sc_hd__o2bb2ai_2
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _354_/X VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_2
X_170_ _370_/Q VGND VGND VPWR VPWR _301_/A sky130_fd_sc_hd__inv_2
X_368_ _328_/A _368_/D _313_/X VGND VGND VPWR VPWR _368_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_299_ _329_/X _299_/B VGND VGND VPWR VPWR _299_/X sky130_fd_sc_hd__and2_2
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_222_ _223_/C VGND VGND VPWR VPWR _288_/A sky130_fd_sc_hd__inv_2
X_205_ _205_/A VGND VGND VPWR VPWR _205_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _348_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _355_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_2
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_367_ _328_/A _367_/D _314_/X VGND VGND VPWR VPWR _367_/Q sky130_fd_sc_hd__dfrtp_2
X_298_ _301_/A _302_/C _221_/A _297_/X _296_/X VGND VGND VPWR VPWR _298_/X sky130_fd_sc_hd__o311a_2
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_221_ _221_/A _221_/B VGND VGND VPWR VPWR _223_/C sky130_fd_sc_hd__or2_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_204_ div[2] _200_/X _203_/A _201_/Y VGND VGND VPWR VPWR _205_/A sky130_fd_sc_hd__o211a_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__332__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _349_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__353__A1 ext_trim[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__344__A1 ext_trim[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__340__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_366_ _328_/A _366_/D _315_/X VGND VGND VPWR VPWR _366_/Q sky130_fd_sc_hd__dfrtp_2
X_297_ _297_/A _368_/Q _297_/C _301_/A VGND VGND VPWR VPWR _297_/X sky130_fd_sc_hd__or4_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__335__A1 ext_trim[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__335__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_220_ _220_/A VGND VGND VPWR VPWR _220_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_349_ _295_/X ext_trim[15] dco VGND VGND VPWR VPWR _349_/X sky130_fd_sc_hd__mux2_1
X_203_ _203_/A VGND VGND VPWR VPWR _203_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.iss.ctrlen0 _182_/B _354_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__343__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XANTENNA__338__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_296_ _367_/Q _221_/B _302_/C _301_/A _295_/X VGND VGND VPWR VPWR _296_/X sky130_fd_sc_hd__o41a_2
X_365_ _328_/A _365_/D _316_/X VGND VGND VPWR VPWR _365_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__351__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ _367_/Q _288_/B VGND VGND VPWR VPWR _279_/X sky130_fd_sc_hd__or2_2
X_348_ _284_/X ext_trim[2] dco VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__mux2_1
X_202_ div[3] _202_/B VGND VGND VPWR VPWR _203_/A sky130_fd_sc_hd__or2_2
XANTENNA__346__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _338_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__354__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__349__S dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_364_ _328_/A _364_/D _317_/X VGND VGND VPWR VPWR _364_/Q sky130_fd_sc_hd__dfrtp_2
X_295_ _301_/A _302_/B _221_/A _294_/X _293_/X VGND VGND VPWR VPWR _295_/X sky130_fd_sc_hd__o311a_2
X_278_ _370_/Q _302_/B VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__or2_2
X_347_ _299_/X ext_trim[16] dco VGND VGND VPWR VPWR _347_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_201_ div[3] _202_/B div[2] _200_/X VGND VGND VPWR VPWR _201_/Y sky130_fd_sc_hd__a22oi_2
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _330_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvp_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _339_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__347__A1 ext_trim[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

