magic
tech sky130A
magscale 1 2
timestamp 1636973520
<< obsli1 >>
rect 1288 1071 68816 3281
<< obsm1 >>
rect 14 552 68816 3460
<< metal2 >>
rect 18 3800 74 4400
rect 294 3800 350 4400
rect 570 3800 626 4400
rect 846 3800 902 4400
rect 1122 3800 1178 4400
rect 1398 3800 1454 4400
rect 1674 3800 1730 4400
rect 1950 3800 2006 4400
rect 2226 3800 2282 4400
rect 2502 3800 2558 4400
rect 2778 3800 2834 4400
rect 3054 3800 3110 4400
rect 3330 3800 3386 4400
rect 3606 3800 3662 4400
rect 3882 3800 3938 4400
rect 4158 3800 4214 4400
rect 4434 3800 4490 4400
rect 4710 3800 4766 4400
rect 4986 3800 5042 4400
rect 5262 3800 5318 4400
rect 5538 3800 5594 4400
rect 5814 3800 5870 4400
rect 6090 3800 6146 4400
rect 6366 3800 6422 4400
rect 6642 3800 6698 4400
rect 6918 3800 6974 4400
rect 7194 3800 7250 4400
rect 7470 3800 7526 4400
rect 7746 3800 7802 4400
rect 8022 3800 8078 4400
rect 8298 3800 8354 4400
rect 8574 3800 8630 4400
rect 8850 3800 8906 4400
rect 9126 3800 9182 4400
rect 9402 3800 9458 4400
rect 9678 3800 9734 4400
rect 9954 3800 10010 4400
rect 10230 3800 10286 4400
rect 10506 3800 10562 4400
rect 10782 3800 10838 4400
rect 11058 3800 11114 4400
rect 11334 3800 11390 4400
rect 11610 3800 11666 4400
rect 11886 3800 11942 4400
rect 12162 3800 12218 4400
rect 12438 3800 12494 4400
rect 12714 3800 12770 4400
rect 12990 3800 13046 4400
rect 13266 3800 13322 4400
rect 13542 3800 13598 4400
rect 13818 3800 13874 4400
rect 14094 3800 14150 4400
rect 14370 3800 14426 4400
rect 14646 3800 14702 4400
rect 14922 3800 14978 4400
rect 15198 3800 15254 4400
rect 15474 3800 15530 4400
rect 15750 3800 15806 4400
rect 16026 3800 16082 4400
rect 16302 3800 16358 4400
rect 16578 3800 16634 4400
rect 16854 3800 16910 4400
rect 17130 3800 17186 4400
rect 17406 3800 17462 4400
rect 17682 3800 17738 4400
rect 17958 3800 18014 4400
rect 18234 3800 18290 4400
rect 18510 3800 18566 4400
rect 18786 3800 18842 4400
rect 19062 3800 19118 4400
rect 19338 3800 19394 4400
rect 19614 3800 19670 4400
rect 19890 3800 19946 4400
rect 20166 3800 20222 4400
rect 20442 3800 20498 4400
rect 20718 3800 20774 4400
rect 20994 3800 21050 4400
rect 21270 3800 21326 4400
rect 21546 3800 21602 4400
rect 21822 3800 21878 4400
rect 22098 3800 22154 4400
rect 22374 3800 22430 4400
rect 22650 3800 22706 4400
rect 22926 3800 22982 4400
rect 23202 3800 23258 4400
rect 23478 3800 23534 4400
rect 23754 3800 23810 4400
rect 24030 3800 24086 4400
rect 24306 3800 24362 4400
rect 24582 3800 24638 4400
rect 24858 3800 24914 4400
rect 25134 3800 25190 4400
rect 25410 3800 25466 4400
rect 25686 3800 25742 4400
rect 25962 3800 26018 4400
rect 26238 3800 26294 4400
rect 26514 3800 26570 4400
rect 26790 3800 26846 4400
rect 27066 3800 27122 4400
rect 27342 3800 27398 4400
rect 27618 3800 27674 4400
rect 27894 3800 27950 4400
rect 28170 3800 28226 4400
rect 28446 3800 28502 4400
rect 28722 3800 28778 4400
rect 28998 3800 29054 4400
rect 29274 3800 29330 4400
rect 29550 3800 29606 4400
rect 29826 3800 29882 4400
rect 30102 3800 30158 4400
rect 30378 3800 30434 4400
rect 30654 3800 30710 4400
rect 30930 3800 30986 4400
rect 31206 3800 31262 4400
rect 31482 3800 31538 4400
rect 31758 3800 31814 4400
rect 32034 3800 32090 4400
rect 32310 3800 32366 4400
rect 32586 3800 32642 4400
rect 32862 3800 32918 4400
rect 33138 3800 33194 4400
rect 33414 3800 33470 4400
rect 33690 3800 33746 4400
rect 33966 3800 34022 4400
rect 34242 3800 34298 4400
rect 34518 3800 34574 4400
rect 34794 3800 34850 4400
rect 35070 3800 35126 4400
rect 35346 3800 35402 4400
rect 35622 3800 35678 4400
rect 35898 3800 35954 4400
rect 36174 3800 36230 4400
rect 36450 3800 36506 4400
rect 36726 3800 36782 4400
rect 37002 3800 37058 4400
rect 37278 3800 37334 4400
rect 37554 3800 37610 4400
rect 37830 3800 37886 4400
rect 38106 3800 38162 4400
rect 38382 3800 38438 4400
rect 38658 3800 38714 4400
rect 38934 3800 38990 4400
rect 39210 3800 39266 4400
rect 39486 3800 39542 4400
rect 39762 3800 39818 4400
rect 40038 3800 40094 4400
rect 40314 3800 40370 4400
rect 40590 3800 40646 4400
rect 40866 3800 40922 4400
rect 41142 3800 41198 4400
rect 41418 3800 41474 4400
rect 41694 3800 41750 4400
rect 41970 3800 42026 4400
rect 42246 3800 42302 4400
rect 42522 3800 42578 4400
rect 42798 3800 42854 4400
rect 43074 3800 43130 4400
rect 43350 3800 43406 4400
rect 43626 3800 43682 4400
rect 43902 3800 43958 4400
rect 44178 3800 44234 4400
rect 44454 3800 44510 4400
rect 44730 3800 44786 4400
rect 45006 3800 45062 4400
rect 45282 3800 45338 4400
rect 45558 3800 45614 4400
rect 45834 3800 45890 4400
rect 46110 3800 46166 4400
rect 46386 3800 46442 4400
rect 46662 3800 46718 4400
rect 46938 3800 46994 4400
rect 47214 3800 47270 4400
rect 47490 3800 47546 4400
rect 47766 3800 47822 4400
rect 48042 3800 48098 4400
rect 48318 3800 48374 4400
rect 48594 3800 48650 4400
rect 48870 3800 48926 4400
rect 49146 3800 49202 4400
rect 49422 3800 49478 4400
rect 49698 3800 49754 4400
rect 49974 3800 50030 4400
rect 50250 3800 50306 4400
rect 50526 3800 50582 4400
rect 50802 3800 50858 4400
rect 51078 3800 51134 4400
rect 51354 3800 51410 4400
rect 51630 3800 51686 4400
rect 51906 3800 51962 4400
rect 52182 3800 52238 4400
rect 52458 3800 52514 4400
rect 52734 3800 52790 4400
rect 53010 3800 53066 4400
rect 53286 3800 53342 4400
rect 53562 3800 53618 4400
rect 53838 3800 53894 4400
rect 54114 3800 54170 4400
rect 54390 3800 54446 4400
rect 54666 3800 54722 4400
rect 54942 3800 54998 4400
rect 55218 3800 55274 4400
rect 55494 3800 55550 4400
rect 55770 3800 55826 4400
rect 56046 3800 56102 4400
rect 56322 3800 56378 4400
rect 56598 3800 56654 4400
rect 56874 3800 56930 4400
rect 57150 3800 57206 4400
rect 57426 3800 57482 4400
rect 57702 3800 57758 4400
rect 57978 3800 58034 4400
rect 58254 3800 58310 4400
rect 58530 3800 58586 4400
rect 58806 3800 58862 4400
rect 59082 3800 59138 4400
rect 59358 3800 59414 4400
rect 59634 3800 59690 4400
rect 59910 3800 59966 4400
rect 60186 3800 60242 4400
rect 60462 3800 60518 4400
rect 60738 3800 60794 4400
rect 61014 3800 61070 4400
rect 61290 3800 61346 4400
rect 61566 3800 61622 4400
rect 61842 3800 61898 4400
rect 62118 3800 62174 4400
rect 62394 3800 62450 4400
rect 62670 3800 62726 4400
rect 62946 3800 63002 4400
rect 63222 3800 63278 4400
rect 63498 3800 63554 4400
rect 63774 3800 63830 4400
rect 64050 3800 64106 4400
rect 64326 3800 64382 4400
rect 64602 3800 64658 4400
rect 64878 3800 64934 4400
rect 65154 3800 65210 4400
rect 65430 3800 65486 4400
rect 65706 3800 65762 4400
rect 65982 3800 66038 4400
rect 66258 3800 66314 4400
rect 66534 3800 66590 4400
rect 66810 3800 66866 4400
rect 67086 3800 67142 4400
rect 67362 3800 67418 4400
rect 67638 3800 67694 4400
rect 67914 3800 67970 4400
rect 7238 1040 7338 3312
rect 13238 1040 13338 3312
rect 19238 1040 19338 3312
rect 25238 1040 25338 3312
rect 31238 1040 31338 3312
rect 37238 1040 37338 3312
rect 43238 1040 43338 3312
rect 49238 1040 49338 3312
rect 55238 1040 55338 3312
rect 61238 1040 61338 3312
rect 67238 1040 67338 3312
rect 18 0 74 600
rect 294 0 350 600
rect 570 0 626 600
rect 846 0 902 600
rect 1122 0 1178 600
rect 1398 0 1454 600
rect 1674 0 1730 600
rect 1950 0 2006 600
rect 2226 0 2282 600
rect 2502 0 2558 600
rect 2778 0 2834 600
rect 3054 0 3110 600
rect 3330 0 3386 600
rect 3606 0 3662 600
rect 3882 0 3938 600
rect 4158 0 4214 600
rect 4434 0 4490 600
rect 4710 0 4766 600
rect 4986 0 5042 600
rect 5262 0 5318 600
rect 5538 0 5594 600
rect 5814 0 5870 600
rect 6090 0 6146 600
rect 6366 0 6422 600
rect 6642 0 6698 600
rect 6918 0 6974 600
rect 7194 0 7250 600
rect 7470 0 7526 600
rect 7746 0 7802 600
rect 8022 0 8078 600
rect 8298 0 8354 600
rect 8574 0 8630 600
rect 8850 0 8906 600
rect 9126 0 9182 600
rect 9402 0 9458 600
rect 9678 0 9734 600
rect 9954 0 10010 600
rect 10230 0 10286 600
rect 10506 0 10562 600
rect 10782 0 10838 600
rect 11058 0 11114 600
rect 11334 0 11390 600
rect 11610 0 11666 600
rect 11886 0 11942 600
rect 12162 0 12218 600
rect 12438 0 12494 600
rect 12714 0 12770 600
rect 12990 0 13046 600
rect 13266 0 13322 600
rect 13542 0 13598 600
rect 13818 0 13874 600
rect 14094 0 14150 600
rect 14370 0 14426 600
rect 14646 0 14702 600
rect 14922 0 14978 600
rect 15198 0 15254 600
rect 15474 0 15530 600
rect 15750 0 15806 600
rect 16026 0 16082 600
rect 16302 0 16358 600
rect 16578 0 16634 600
rect 16854 0 16910 600
rect 17130 0 17186 600
rect 17406 0 17462 600
rect 17682 0 17738 600
rect 17958 0 18014 600
rect 18234 0 18290 600
rect 18510 0 18566 600
rect 18786 0 18842 600
rect 19062 0 19118 600
rect 19338 0 19394 600
rect 19614 0 19670 600
rect 19890 0 19946 600
rect 20166 0 20222 600
rect 20442 0 20498 600
rect 20718 0 20774 600
rect 20994 0 21050 600
rect 21270 0 21326 600
rect 21546 0 21602 600
rect 21822 0 21878 600
rect 22098 0 22154 600
rect 22374 0 22430 600
rect 22650 0 22706 600
rect 22926 0 22982 600
rect 23202 0 23258 600
rect 23478 0 23534 600
rect 23754 0 23810 600
rect 24030 0 24086 600
rect 24306 0 24362 600
rect 24582 0 24638 600
rect 24858 0 24914 600
rect 25134 0 25190 600
rect 25410 0 25466 600
rect 25686 0 25742 600
rect 25962 0 26018 600
rect 26238 0 26294 600
rect 26514 0 26570 600
rect 26790 0 26846 600
rect 27066 0 27122 600
rect 27342 0 27398 600
rect 27618 0 27674 600
rect 27894 0 27950 600
rect 28170 0 28226 600
rect 28446 0 28502 600
rect 28722 0 28778 600
rect 28998 0 29054 600
rect 29274 0 29330 600
rect 29550 0 29606 600
rect 29826 0 29882 600
rect 30102 0 30158 600
rect 30378 0 30434 600
rect 30654 0 30710 600
rect 30930 0 30986 600
rect 31206 0 31262 600
rect 31482 0 31538 600
rect 31758 0 31814 600
rect 32034 0 32090 600
rect 32310 0 32366 600
rect 32586 0 32642 600
rect 32862 0 32918 600
rect 33138 0 33194 600
rect 33414 0 33470 600
rect 33690 0 33746 600
rect 33966 0 34022 600
rect 34242 0 34298 600
rect 34518 0 34574 600
rect 34794 0 34850 600
rect 35070 0 35126 600
rect 35346 0 35402 600
rect 35622 0 35678 600
rect 35898 0 35954 600
rect 36174 0 36230 600
rect 36450 0 36506 600
rect 36726 0 36782 600
rect 37002 0 37058 600
rect 37278 0 37334 600
rect 37554 0 37610 600
rect 37830 0 37886 600
rect 38106 0 38162 600
rect 38382 0 38438 600
rect 38658 0 38714 600
rect 38934 0 38990 600
rect 39210 0 39266 600
rect 39486 0 39542 600
rect 39762 0 39818 600
rect 40038 0 40094 600
rect 40314 0 40370 600
rect 40590 0 40646 600
rect 40866 0 40922 600
rect 41142 0 41198 600
rect 41418 0 41474 600
rect 41694 0 41750 600
rect 41970 0 42026 600
rect 42246 0 42302 600
rect 42522 0 42578 600
rect 42798 0 42854 600
rect 43074 0 43130 600
rect 43350 0 43406 600
rect 43626 0 43682 600
rect 43902 0 43958 600
rect 44178 0 44234 600
rect 44454 0 44510 600
rect 44730 0 44786 600
rect 45006 0 45062 600
rect 45282 0 45338 600
rect 45558 0 45614 600
rect 45834 0 45890 600
rect 46110 0 46166 600
rect 46386 0 46442 600
rect 46662 0 46718 600
rect 46938 0 46994 600
rect 47214 0 47270 600
rect 47490 0 47546 600
rect 47766 0 47822 600
rect 48042 0 48098 600
rect 48318 0 48374 600
rect 48594 0 48650 600
rect 48870 0 48926 600
rect 49146 0 49202 600
rect 49422 0 49478 600
rect 49698 0 49754 600
rect 49974 0 50030 600
rect 50250 0 50306 600
rect 50526 0 50582 600
rect 50802 0 50858 600
rect 51078 0 51134 600
rect 51354 0 51410 600
rect 51630 0 51686 600
rect 51906 0 51962 600
rect 52182 0 52238 600
rect 52458 0 52514 600
rect 52734 0 52790 600
rect 53010 0 53066 600
rect 53286 0 53342 600
rect 53562 0 53618 600
rect 53838 0 53894 600
rect 54114 0 54170 600
rect 54390 0 54446 600
rect 54666 0 54722 600
rect 54942 0 54998 600
<< obsm2 >>
rect 130 3744 238 3800
rect 406 3744 514 3800
rect 682 3744 790 3800
rect 958 3744 1066 3800
rect 1234 3744 1342 3800
rect 1510 3744 1618 3800
rect 1786 3744 1894 3800
rect 2062 3744 2170 3800
rect 2338 3744 2446 3800
rect 2614 3744 2722 3800
rect 2890 3744 2998 3800
rect 3166 3744 3274 3800
rect 3442 3744 3550 3800
rect 3718 3744 3826 3800
rect 3994 3744 4102 3800
rect 4270 3744 4378 3800
rect 4546 3744 4654 3800
rect 4822 3744 4930 3800
rect 5098 3744 5206 3800
rect 5374 3744 5482 3800
rect 5650 3744 5758 3800
rect 5926 3744 6034 3800
rect 6202 3744 6310 3800
rect 6478 3744 6586 3800
rect 6754 3744 6862 3800
rect 7030 3744 7138 3800
rect 7306 3744 7414 3800
rect 7582 3744 7690 3800
rect 7858 3744 7966 3800
rect 8134 3744 8242 3800
rect 8410 3744 8518 3800
rect 8686 3744 8794 3800
rect 8962 3744 9070 3800
rect 9238 3744 9346 3800
rect 9514 3744 9622 3800
rect 9790 3744 9898 3800
rect 10066 3744 10174 3800
rect 10342 3744 10450 3800
rect 10618 3744 10726 3800
rect 10894 3744 11002 3800
rect 11170 3744 11278 3800
rect 11446 3744 11554 3800
rect 11722 3744 11830 3800
rect 11998 3744 12106 3800
rect 12274 3744 12382 3800
rect 12550 3744 12658 3800
rect 12826 3744 12934 3800
rect 13102 3744 13210 3800
rect 13378 3744 13486 3800
rect 13654 3744 13762 3800
rect 13930 3744 14038 3800
rect 14206 3744 14314 3800
rect 14482 3744 14590 3800
rect 14758 3744 14866 3800
rect 15034 3744 15142 3800
rect 15310 3744 15418 3800
rect 15586 3744 15694 3800
rect 15862 3744 15970 3800
rect 16138 3744 16246 3800
rect 16414 3744 16522 3800
rect 16690 3744 16798 3800
rect 16966 3744 17074 3800
rect 17242 3744 17350 3800
rect 17518 3744 17626 3800
rect 17794 3744 17902 3800
rect 18070 3744 18178 3800
rect 18346 3744 18454 3800
rect 18622 3744 18730 3800
rect 18898 3744 19006 3800
rect 19174 3744 19282 3800
rect 19450 3744 19558 3800
rect 19726 3744 19834 3800
rect 20002 3744 20110 3800
rect 20278 3744 20386 3800
rect 20554 3744 20662 3800
rect 20830 3744 20938 3800
rect 21106 3744 21214 3800
rect 21382 3744 21490 3800
rect 21658 3744 21766 3800
rect 21934 3744 22042 3800
rect 22210 3744 22318 3800
rect 22486 3744 22594 3800
rect 22762 3744 22870 3800
rect 23038 3744 23146 3800
rect 23314 3744 23422 3800
rect 23590 3744 23698 3800
rect 23866 3744 23974 3800
rect 24142 3744 24250 3800
rect 24418 3744 24526 3800
rect 24694 3744 24802 3800
rect 24970 3744 25078 3800
rect 25246 3744 25354 3800
rect 25522 3744 25630 3800
rect 25798 3744 25906 3800
rect 26074 3744 26182 3800
rect 26350 3744 26458 3800
rect 26626 3744 26734 3800
rect 26902 3744 27010 3800
rect 27178 3744 27286 3800
rect 27454 3744 27562 3800
rect 27730 3744 27838 3800
rect 28006 3744 28114 3800
rect 28282 3744 28390 3800
rect 28558 3744 28666 3800
rect 28834 3744 28942 3800
rect 29110 3744 29218 3800
rect 29386 3744 29494 3800
rect 29662 3744 29770 3800
rect 29938 3744 30046 3800
rect 30214 3744 30322 3800
rect 30490 3744 30598 3800
rect 30766 3744 30874 3800
rect 31042 3744 31150 3800
rect 31318 3744 31426 3800
rect 31594 3744 31702 3800
rect 31870 3744 31978 3800
rect 32146 3744 32254 3800
rect 32422 3744 32530 3800
rect 32698 3744 32806 3800
rect 32974 3744 33082 3800
rect 33250 3744 33358 3800
rect 33526 3744 33634 3800
rect 33802 3744 33910 3800
rect 34078 3744 34186 3800
rect 34354 3744 34462 3800
rect 34630 3744 34738 3800
rect 34906 3744 35014 3800
rect 35182 3744 35290 3800
rect 35458 3744 35566 3800
rect 35734 3744 35842 3800
rect 36010 3744 36118 3800
rect 36286 3744 36394 3800
rect 36562 3744 36670 3800
rect 36838 3744 36946 3800
rect 37114 3744 37222 3800
rect 37390 3744 37498 3800
rect 37666 3744 37774 3800
rect 37942 3744 38050 3800
rect 38218 3744 38326 3800
rect 38494 3744 38602 3800
rect 38770 3744 38878 3800
rect 39046 3744 39154 3800
rect 39322 3744 39430 3800
rect 39598 3744 39706 3800
rect 39874 3744 39982 3800
rect 40150 3744 40258 3800
rect 40426 3744 40534 3800
rect 40702 3744 40810 3800
rect 40978 3744 41086 3800
rect 41254 3744 41362 3800
rect 41530 3744 41638 3800
rect 41806 3744 41914 3800
rect 42082 3744 42190 3800
rect 42358 3744 42466 3800
rect 42634 3744 42742 3800
rect 42910 3744 43018 3800
rect 43186 3744 43294 3800
rect 43462 3744 43570 3800
rect 43738 3744 43846 3800
rect 44014 3744 44122 3800
rect 44290 3744 44398 3800
rect 44566 3744 44674 3800
rect 44842 3744 44950 3800
rect 45118 3744 45226 3800
rect 45394 3744 45502 3800
rect 45670 3744 45778 3800
rect 45946 3744 46054 3800
rect 46222 3744 46330 3800
rect 46498 3744 46606 3800
rect 46774 3744 46882 3800
rect 47050 3744 47158 3800
rect 47326 3744 47434 3800
rect 47602 3744 47710 3800
rect 47878 3744 47986 3800
rect 48154 3744 48262 3800
rect 48430 3744 48538 3800
rect 48706 3744 48814 3800
rect 48982 3744 49090 3800
rect 49258 3744 49366 3800
rect 49534 3744 49642 3800
rect 49810 3744 49918 3800
rect 50086 3744 50194 3800
rect 50362 3744 50470 3800
rect 50638 3744 50746 3800
rect 50914 3744 51022 3800
rect 51190 3744 51298 3800
rect 51466 3744 51574 3800
rect 51742 3744 51850 3800
rect 52018 3744 52126 3800
rect 52294 3744 52402 3800
rect 52570 3744 52678 3800
rect 52846 3744 52954 3800
rect 53122 3744 53230 3800
rect 53398 3744 53506 3800
rect 53674 3744 53782 3800
rect 53950 3744 54058 3800
rect 54226 3744 54334 3800
rect 54502 3744 54610 3800
rect 54778 3744 54886 3800
rect 55054 3744 55162 3800
rect 55330 3744 55438 3800
rect 55606 3744 55714 3800
rect 55882 3744 55990 3800
rect 56158 3744 56266 3800
rect 56434 3744 56542 3800
rect 56710 3744 56818 3800
rect 56986 3744 57094 3800
rect 57262 3744 57370 3800
rect 57538 3744 57646 3800
rect 57814 3744 57922 3800
rect 58090 3744 58198 3800
rect 58366 3744 58474 3800
rect 58642 3744 58750 3800
rect 58918 3744 59026 3800
rect 59194 3744 59302 3800
rect 59470 3744 59578 3800
rect 59746 3744 59854 3800
rect 60022 3744 60130 3800
rect 60298 3744 60406 3800
rect 60574 3744 60682 3800
rect 60850 3744 60958 3800
rect 61126 3744 61234 3800
rect 61402 3744 61510 3800
rect 61678 3744 61786 3800
rect 61954 3744 62062 3800
rect 62230 3744 62338 3800
rect 62506 3744 62614 3800
rect 62782 3744 62890 3800
rect 63058 3744 63166 3800
rect 63334 3744 63442 3800
rect 63610 3744 63718 3800
rect 63886 3744 63994 3800
rect 64162 3744 64270 3800
rect 64438 3744 64546 3800
rect 64714 3744 64822 3800
rect 64990 3744 65098 3800
rect 65266 3744 65374 3800
rect 65542 3744 65650 3800
rect 65818 3744 65926 3800
rect 66094 3744 66202 3800
rect 66370 3744 66478 3800
rect 66646 3744 66754 3800
rect 66922 3744 67030 3800
rect 67198 3744 67306 3800
rect 67474 3744 67582 3800
rect 67750 3744 67858 3800
rect 20 3368 67968 3744
rect 20 984 7182 3368
rect 7394 984 13182 3368
rect 13394 984 19182 3368
rect 19394 984 25182 3368
rect 25394 984 31182 3368
rect 31394 984 37182 3368
rect 37394 984 43182 3368
rect 43394 984 49182 3368
rect 49394 984 55182 3368
rect 55394 984 61182 3368
rect 61394 984 67182 3368
rect 67394 984 67968 3368
rect 20 656 67968 984
rect 130 546 238 656
rect 406 546 514 656
rect 682 546 790 656
rect 958 546 1066 656
rect 1234 546 1342 656
rect 1510 546 1618 656
rect 1786 546 1894 656
rect 2062 546 2170 656
rect 2338 546 2446 656
rect 2614 546 2722 656
rect 2890 546 2998 656
rect 3166 546 3274 656
rect 3442 546 3550 656
rect 3718 546 3826 656
rect 3994 546 4102 656
rect 4270 546 4378 656
rect 4546 546 4654 656
rect 4822 546 4930 656
rect 5098 546 5206 656
rect 5374 546 5482 656
rect 5650 546 5758 656
rect 5926 546 6034 656
rect 6202 546 6310 656
rect 6478 546 6586 656
rect 6754 546 6862 656
rect 7030 546 7138 656
rect 7306 546 7414 656
rect 7582 546 7690 656
rect 7858 546 7966 656
rect 8134 546 8242 656
rect 8410 546 8518 656
rect 8686 546 8794 656
rect 8962 546 9070 656
rect 9238 546 9346 656
rect 9514 546 9622 656
rect 9790 546 9898 656
rect 10066 546 10174 656
rect 10342 546 10450 656
rect 10618 546 10726 656
rect 10894 546 11002 656
rect 11170 546 11278 656
rect 11446 546 11554 656
rect 11722 546 11830 656
rect 11998 546 12106 656
rect 12274 546 12382 656
rect 12550 546 12658 656
rect 12826 546 12934 656
rect 13102 546 13210 656
rect 13378 546 13486 656
rect 13654 546 13762 656
rect 13930 546 14038 656
rect 14206 546 14314 656
rect 14482 546 14590 656
rect 14758 546 14866 656
rect 15034 546 15142 656
rect 15310 546 15418 656
rect 15586 546 15694 656
rect 15862 546 15970 656
rect 16138 546 16246 656
rect 16414 546 16522 656
rect 16690 546 16798 656
rect 16966 546 17074 656
rect 17242 546 17350 656
rect 17518 546 17626 656
rect 17794 546 17902 656
rect 18070 546 18178 656
rect 18346 546 18454 656
rect 18622 546 18730 656
rect 18898 546 19006 656
rect 19174 546 19282 656
rect 19450 546 19558 656
rect 19726 546 19834 656
rect 20002 546 20110 656
rect 20278 546 20386 656
rect 20554 546 20662 656
rect 20830 546 20938 656
rect 21106 546 21214 656
rect 21382 546 21490 656
rect 21658 546 21766 656
rect 21934 546 22042 656
rect 22210 546 22318 656
rect 22486 546 22594 656
rect 22762 546 22870 656
rect 23038 546 23146 656
rect 23314 546 23422 656
rect 23590 546 23698 656
rect 23866 546 23974 656
rect 24142 546 24250 656
rect 24418 546 24526 656
rect 24694 546 24802 656
rect 24970 546 25078 656
rect 25246 546 25354 656
rect 25522 546 25630 656
rect 25798 546 25906 656
rect 26074 546 26182 656
rect 26350 546 26458 656
rect 26626 546 26734 656
rect 26902 546 27010 656
rect 27178 546 27286 656
rect 27454 546 27562 656
rect 27730 546 27838 656
rect 28006 546 28114 656
rect 28282 546 28390 656
rect 28558 546 28666 656
rect 28834 546 28942 656
rect 29110 546 29218 656
rect 29386 546 29494 656
rect 29662 546 29770 656
rect 29938 546 30046 656
rect 30214 546 30322 656
rect 30490 546 30598 656
rect 30766 546 30874 656
rect 31042 546 31150 656
rect 31318 546 31426 656
rect 31594 546 31702 656
rect 31870 546 31978 656
rect 32146 546 32254 656
rect 32422 546 32530 656
rect 32698 546 32806 656
rect 32974 546 33082 656
rect 33250 546 33358 656
rect 33526 546 33634 656
rect 33802 546 33910 656
rect 34078 546 34186 656
rect 34354 546 34462 656
rect 34630 546 34738 656
rect 34906 546 35014 656
rect 35182 546 35290 656
rect 35458 546 35566 656
rect 35734 546 35842 656
rect 36010 546 36118 656
rect 36286 546 36394 656
rect 36562 546 36670 656
rect 36838 546 36946 656
rect 37114 546 37222 656
rect 37390 546 37498 656
rect 37666 546 37774 656
rect 37942 546 38050 656
rect 38218 546 38326 656
rect 38494 546 38602 656
rect 38770 546 38878 656
rect 39046 546 39154 656
rect 39322 546 39430 656
rect 39598 546 39706 656
rect 39874 546 39982 656
rect 40150 546 40258 656
rect 40426 546 40534 656
rect 40702 546 40810 656
rect 40978 546 41086 656
rect 41254 546 41362 656
rect 41530 546 41638 656
rect 41806 546 41914 656
rect 42082 546 42190 656
rect 42358 546 42466 656
rect 42634 546 42742 656
rect 42910 546 43018 656
rect 43186 546 43294 656
rect 43462 546 43570 656
rect 43738 546 43846 656
rect 44014 546 44122 656
rect 44290 546 44398 656
rect 44566 546 44674 656
rect 44842 546 44950 656
rect 45118 546 45226 656
rect 45394 546 45502 656
rect 45670 546 45778 656
rect 45946 546 46054 656
rect 46222 546 46330 656
rect 46498 546 46606 656
rect 46774 546 46882 656
rect 47050 546 47158 656
rect 47326 546 47434 656
rect 47602 546 47710 656
rect 47878 546 47986 656
rect 48154 546 48262 656
rect 48430 546 48538 656
rect 48706 546 48814 656
rect 48982 546 49090 656
rect 49258 546 49366 656
rect 49534 546 49642 656
rect 49810 546 49918 656
rect 50086 546 50194 656
rect 50362 546 50470 656
rect 50638 546 50746 656
rect 50914 546 51022 656
rect 51190 546 51298 656
rect 51466 546 51574 656
rect 51742 546 51850 656
rect 52018 546 52126 656
rect 52294 546 52402 656
rect 52570 546 52678 656
rect 52846 546 52954 656
rect 53122 546 53230 656
rect 53398 546 53506 656
rect 53674 546 53782 656
rect 53950 546 54058 656
rect 54226 546 54334 656
rect 54502 546 54610 656
rect 54778 546 54886 656
rect 55054 546 67968 656
<< metal3 >>
rect 0 4088 600 4208
rect 0 3816 600 3936
rect 0 3544 600 3664
rect 0 3272 600 3392
rect 0 3000 600 3120
rect 0 2728 600 2848
rect 0 2456 600 2576
rect 0 2184 600 2304
rect 1288 2270 68816 2370
rect 0 1912 600 2032
rect 0 1640 600 1760
rect 0 1368 600 1488
rect 0 1096 600 1216
rect 1288 1190 68816 1290
rect 0 824 600 944
rect 0 552 600 672
rect 0 280 600 400
rect 0 8 600 128
<< obsm3 >>
rect 680 2450 4311 4178
rect 680 2190 1208 2450
rect 680 1370 4311 2190
rect 680 1110 1208 1370
rect 680 38 4311 1110
<< labels >>
rlabel metal3 s 0 3816 600 3936 6 HI[0]
port 1 nsew signal output
rlabel metal3 s 0 3544 600 3664 6 HI[100]
port 2 nsew signal output
rlabel metal3 s 0 3272 600 3392 6 HI[101]
port 3 nsew signal output
rlabel metal3 s 0 3000 600 3120 6 HI[102]
port 4 nsew signal output
rlabel metal3 s 0 2728 600 2848 6 HI[103]
port 5 nsew signal output
rlabel metal3 s 0 2456 600 2576 6 HI[104]
port 6 nsew signal output
rlabel metal3 s 0 2184 600 2304 6 HI[105]
port 7 nsew signal output
rlabel metal3 s 0 1912 600 2032 6 HI[106]
port 8 nsew signal output
rlabel metal3 s 0 1640 600 1760 6 HI[107]
port 9 nsew signal output
rlabel metal3 s 0 1368 600 1488 6 HI[108]
port 10 nsew signal output
rlabel metal3 s 0 1096 600 1216 6 HI[109]
port 11 nsew signal output
rlabel metal3 s 0 4088 600 4208 6 HI[10]
port 12 nsew signal output
rlabel metal3 s 0 824 600 944 6 HI[110]
port 13 nsew signal output
rlabel metal3 s 0 280 600 400 6 HI[111]
port 14 nsew signal output
rlabel metal3 s 0 8 600 128 6 HI[112]
port 15 nsew signal output
rlabel metal3 s 0 552 600 672 6 HI[113]
port 16 nsew signal output
rlabel metal2 s 14094 3800 14150 4400 6 HI[114]
port 17 nsew signal output
rlabel metal2 s 12990 3800 13046 4400 6 HI[115]
port 18 nsew signal output
rlabel metal2 s 13818 3800 13874 4400 6 HI[116]
port 19 nsew signal output
rlabel metal2 s 13542 3800 13598 4400 6 HI[117]
port 20 nsew signal output
rlabel metal2 s 9402 3800 9458 4400 6 HI[118]
port 21 nsew signal output
rlabel metal2 s 13266 3800 13322 4400 6 HI[119]
port 22 nsew signal output
rlabel metal2 s 12438 3800 12494 4400 6 HI[11]
port 23 nsew signal output
rlabel metal2 s 11334 3800 11390 4400 6 HI[120]
port 24 nsew signal output
rlabel metal2 s 12714 3800 12770 4400 6 HI[121]
port 25 nsew signal output
rlabel metal2 s 6366 3800 6422 4400 6 HI[122]
port 26 nsew signal output
rlabel metal2 s 12162 3800 12218 4400 6 HI[123]
port 27 nsew signal output
rlabel metal2 s 11886 3800 11942 4400 6 HI[124]
port 28 nsew signal output
rlabel metal2 s 11610 3800 11666 4400 6 HI[125]
port 29 nsew signal output
rlabel metal2 s 9678 3800 9734 4400 6 HI[126]
port 30 nsew signal output
rlabel metal2 s 11058 3800 11114 4400 6 HI[127]
port 31 nsew signal output
rlabel metal2 s 10782 3800 10838 4400 6 HI[128]
port 32 nsew signal output
rlabel metal2 s 10506 3800 10562 4400 6 HI[129]
port 33 nsew signal output
rlabel metal2 s 570 3800 626 4400 6 HI[12]
port 34 nsew signal output
rlabel metal2 s 10230 3800 10286 4400 6 HI[130]
port 35 nsew signal output
rlabel metal2 s 9954 3800 10010 4400 6 HI[131]
port 36 nsew signal output
rlabel metal2 s 7746 3800 7802 4400 6 HI[132]
port 37 nsew signal output
rlabel metal2 s 4986 3800 5042 4400 6 HI[133]
port 38 nsew signal output
rlabel metal2 s 9126 3800 9182 4400 6 HI[134]
port 39 nsew signal output
rlabel metal2 s 8850 3800 8906 4400 6 HI[135]
port 40 nsew signal output
rlabel metal2 s 8574 3800 8630 4400 6 HI[136]
port 41 nsew signal output
rlabel metal2 s 8298 3800 8354 4400 6 HI[137]
port 42 nsew signal output
rlabel metal2 s 8022 3800 8078 4400 6 HI[138]
port 43 nsew signal output
rlabel metal2 s 5814 3800 5870 4400 6 HI[139]
port 44 nsew signal output
rlabel metal2 s 14370 3800 14426 4400 6 HI[13]
port 45 nsew signal output
rlabel metal2 s 7470 3800 7526 4400 6 HI[140]
port 46 nsew signal output
rlabel metal2 s 7194 3800 7250 4400 6 HI[141]
port 47 nsew signal output
rlabel metal2 s 6918 3800 6974 4400 6 HI[142]
port 48 nsew signal output
rlabel metal2 s 6642 3800 6698 4400 6 HI[143]
port 49 nsew signal output
rlabel metal2 s 18 3800 74 4400 6 HI[144]
port 50 nsew signal output
rlabel metal2 s 6090 3800 6146 4400 6 HI[145]
port 51 nsew signal output
rlabel metal2 s 3606 3800 3662 4400 6 HI[146]
port 52 nsew signal output
rlabel metal2 s 5538 3800 5594 4400 6 HI[147]
port 53 nsew signal output
rlabel metal2 s 5262 3800 5318 4400 6 HI[148]
port 54 nsew signal output
rlabel metal2 s 294 3800 350 4400 6 HI[149]
port 55 nsew signal output
rlabel metal2 s 4434 3800 4490 4400 6 HI[14]
port 56 nsew signal output
rlabel metal2 s 4710 3800 4766 4400 6 HI[150]
port 57 nsew signal output
rlabel metal2 s 3882 3800 3938 4400 6 HI[151]
port 58 nsew signal output
rlabel metal2 s 4158 3800 4214 4400 6 HI[152]
port 59 nsew signal output
rlabel metal2 s 3330 3800 3386 4400 6 HI[153]
port 60 nsew signal output
rlabel metal2 s 1122 3800 1178 4400 6 HI[154]
port 61 nsew signal output
rlabel metal2 s 3054 3800 3110 4400 6 HI[155]
port 62 nsew signal output
rlabel metal2 s 2778 3800 2834 4400 6 HI[156]
port 63 nsew signal output
rlabel metal2 s 2502 3800 2558 4400 6 HI[157]
port 64 nsew signal output
rlabel metal2 s 2226 3800 2282 4400 6 HI[158]
port 65 nsew signal output
rlabel metal2 s 1950 3800 2006 4400 6 HI[159]
port 66 nsew signal output
rlabel metal2 s 14646 3800 14702 4400 6 HI[15]
port 67 nsew signal output
rlabel metal2 s 1398 3800 1454 4400 6 HI[160]
port 68 nsew signal output
rlabel metal2 s 1674 3800 1730 4400 6 HI[161]
port 69 nsew signal output
rlabel metal2 s 846 3800 902 4400 6 HI[162]
port 70 nsew signal output
rlabel metal2 s 11886 0 11942 600 6 HI[163]
port 71 nsew signal output
rlabel metal2 s 28998 0 29054 600 6 HI[164]
port 72 nsew signal output
rlabel metal2 s 17958 0 18014 600 6 HI[165]
port 73 nsew signal output
rlabel metal2 s 11058 0 11114 600 6 HI[166]
port 74 nsew signal output
rlabel metal2 s 45282 0 45338 600 6 HI[167]
port 75 nsew signal output
rlabel metal2 s 7746 0 7802 600 6 HI[168]
port 76 nsew signal output
rlabel metal2 s 8574 0 8630 600 6 HI[169]
port 77 nsew signal output
rlabel metal2 s 29550 0 29606 600 6 HI[16]
port 78 nsew signal output
rlabel metal2 s 45558 0 45614 600 6 HI[170]
port 79 nsew signal output
rlabel metal2 s 10782 0 10838 600 6 HI[171]
port 80 nsew signal output
rlabel metal2 s 29826 0 29882 600 6 HI[172]
port 81 nsew signal output
rlabel metal2 s 51354 0 51410 600 6 HI[173]
port 82 nsew signal output
rlabel metal2 s 10230 0 10286 600 6 HI[174]
port 83 nsew signal output
rlabel metal2 s 54666 0 54722 600 6 HI[175]
port 84 nsew signal output
rlabel metal2 s 19062 0 19118 600 6 HI[176]
port 85 nsew signal output
rlabel metal2 s 6366 0 6422 600 6 HI[177]
port 86 nsew signal output
rlabel metal2 s 30378 0 30434 600 6 HI[178]
port 87 nsew signal output
rlabel metal2 s 8298 0 8354 600 6 HI[179]
port 88 nsew signal output
rlabel metal2 s 294 0 350 600 6 HI[17]
port 89 nsew signal output
rlabel metal2 s 46110 0 46166 600 6 HI[180]
port 90 nsew signal output
rlabel metal2 s 23754 0 23810 600 6 HI[181]
port 91 nsew signal output
rlabel metal2 s 14094 0 14150 600 6 HI[182]
port 92 nsew signal output
rlabel metal2 s 30930 0 30986 600 6 HI[183]
port 93 nsew signal output
rlabel metal2 s 51630 0 51686 600 6 HI[184]
port 94 nsew signal output
rlabel metal2 s 6090 0 6146 600 6 HI[185]
port 95 nsew signal output
rlabel metal2 s 31206 0 31262 600 6 HI[186]
port 96 nsew signal output
rlabel metal2 s 46386 0 46442 600 6 HI[187]
port 97 nsew signal output
rlabel metal2 s 13818 0 13874 600 6 HI[188]
port 98 nsew signal output
rlabel metal2 s 31482 0 31538 600 6 HI[189]
port 99 nsew signal output
rlabel metal2 s 2778 0 2834 600 6 HI[18]
port 100 nsew signal output
rlabel metal2 s 16854 0 16910 600 6 HI[190]
port 101 nsew signal output
rlabel metal2 s 46662 0 46718 600 6 HI[191]
port 102 nsew signal output
rlabel metal2 s 20718 0 20774 600 6 HI[192]
port 103 nsew signal output
rlabel metal2 s 11334 0 11390 600 6 HI[193]
port 104 nsew signal output
rlabel metal2 s 51906 0 51962 600 6 HI[194]
port 105 nsew signal output
rlabel metal2 s 8850 0 8906 600 6 HI[195]
port 106 nsew signal output
rlabel metal2 s 9126 0 9182 600 6 HI[196]
port 107 nsew signal output
rlabel metal2 s 32310 0 32366 600 6 HI[197]
port 108 nsew signal output
rlabel metal2 s 21270 0 21326 600 6 HI[198]
port 109 nsew signal output
rlabel metal2 s 46938 0 46994 600 6 HI[199]
port 110 nsew signal output
rlabel metal2 s 32586 0 32642 600 6 HI[19]
port 111 nsew signal output
rlabel metal2 s 52182 0 52238 600 6 HI[1]
port 112 nsew signal output
rlabel metal2 s 12990 0 13046 600 6 HI[200]
port 113 nsew signal output
rlabel metal2 s 32862 0 32918 600 6 HI[201]
port 114 nsew signal output
rlabel metal2 s 21822 0 21878 600 6 HI[202]
port 115 nsew signal output
rlabel metal2 s 47214 0 47270 600 6 HI[203]
port 116 nsew signal output
rlabel metal2 s 33138 0 33194 600 6 HI[204]
port 117 nsew signal output
rlabel metal2 s 24858 0 24914 600 6 HI[205]
port 118 nsew signal output
rlabel metal2 s 4986 0 5042 600 6 HI[206]
port 119 nsew signal output
rlabel metal2 s 47490 0 47546 600 6 HI[207]
port 120 nsew signal output
rlabel metal2 s 22374 0 22430 600 6 HI[208]
port 121 nsew signal output
rlabel metal2 s 846 0 902 600 6 HI[209]
port 122 nsew signal output
rlabel metal2 s 54114 0 54170 600 6 HI[20]
port 123 nsew signal output
rlabel metal2 s 2226 0 2282 600 6 HI[210]
port 124 nsew signal output
rlabel metal2 s 47766 0 47822 600 6 HI[211]
port 125 nsew signal output
rlabel metal2 s 33966 0 34022 600 6 HI[212]
port 126 nsew signal output
rlabel metal2 s 22926 0 22982 600 6 HI[213]
port 127 nsew signal output
rlabel metal2 s 4434 0 4490 600 6 HI[214]
port 128 nsew signal output
rlabel metal2 s 34242 0 34298 600 6 HI[215]
port 129 nsew signal output
rlabel metal2 s 48042 0 48098 600 6 HI[216]
port 130 nsew signal output
rlabel metal2 s 18510 0 18566 600 6 HI[217]
port 131 nsew signal output
rlabel metal2 s 34518 0 34574 600 6 HI[218]
port 132 nsew signal output
rlabel metal2 s 23478 0 23534 600 6 HI[219]
port 133 nsew signal output
rlabel metal2 s 48318 0 48374 600 6 HI[21]
port 134 nsew signal output
rlabel metal2 s 34794 0 34850 600 6 HI[220]
port 135 nsew signal output
rlabel metal2 s 7470 0 7526 600 6 HI[221]
port 136 nsew signal output
rlabel metal2 s 5538 0 5594 600 6 HI[222]
port 137 nsew signal output
rlabel metal2 s 35070 0 35126 600 6 HI[223]
port 138 nsew signal output
rlabel metal2 s 24030 0 24086 600 6 HI[224]
port 139 nsew signal output
rlabel metal2 s 52458 0 52514 600 6 HI[225]
port 140 nsew signal output
rlabel metal2 s 35346 0 35402 600 6 HI[226]
port 141 nsew signal output
rlabel metal2 s 28722 0 28778 600 6 HI[227]
port 142 nsew signal output
rlabel metal2 s 18 0 74 600 6 HI[228]
port 143 nsew signal output
rlabel metal2 s 35622 0 35678 600 6 HI[229]
port 144 nsew signal output
rlabel metal2 s 24582 0 24638 600 6 HI[22]
port 145 nsew signal output
rlabel metal2 s 12714 0 12770 600 6 HI[230]
port 146 nsew signal output
rlabel metal2 s 35898 0 35954 600 6 HI[231]
port 147 nsew signal output
rlabel metal2 s 39210 0 39266 600 6 HI[232]
port 148 nsew signal output
rlabel metal2 s 48594 0 48650 600 6 HI[233]
port 149 nsew signal output
rlabel metal2 s 36174 0 36230 600 6 HI[234]
port 150 nsew signal output
rlabel metal2 s 25134 0 25190 600 6 HI[235]
port 151 nsew signal output
rlabel metal2 s 20166 0 20222 600 6 HI[236]
port 152 nsew signal output
rlabel metal2 s 36450 0 36506 600 6 HI[237]
port 153 nsew signal output
rlabel metal2 s 52734 0 52790 600 6 HI[238]
port 154 nsew signal output
rlabel metal2 s 54942 0 54998 600 6 HI[239]
port 155 nsew signal output
rlabel metal2 s 36726 0 36782 600 6 HI[23]
port 156 nsew signal output
rlabel metal2 s 25686 0 25742 600 6 HI[240]
port 157 nsew signal output
rlabel metal2 s 12162 0 12218 600 6 HI[241]
port 158 nsew signal output
rlabel metal2 s 37002 0 37058 600 6 HI[242]
port 159 nsew signal output
rlabel metal2 s 13266 0 13322 600 6 HI[243]
port 160 nsew signal output
rlabel metal2 s 20994 0 21050 600 6 HI[244]
port 161 nsew signal output
rlabel metal2 s 37278 0 37334 600 6 HI[245]
port 162 nsew signal output
rlabel metal2 s 26238 0 26294 600 6 HI[246]
port 163 nsew signal output
rlabel metal2 s 14646 0 14702 600 6 HI[247]
port 164 nsew signal output
rlabel metal2 s 37554 0 37610 600 6 HI[248]
port 165 nsew signal output
rlabel metal2 s 53010 0 53066 600 6 HI[249]
port 166 nsew signal output
rlabel metal2 s 33414 0 33470 600 6 HI[24]
port 167 nsew signal output
rlabel metal2 s 37830 0 37886 600 6 HI[250]
port 168 nsew signal output
rlabel metal2 s 26790 0 26846 600 6 HI[251]
port 169 nsew signal output
rlabel metal2 s 22098 0 22154 600 6 HI[252]
port 170 nsew signal output
rlabel metal2 s 38106 0 38162 600 6 HI[253]
port 171 nsew signal output
rlabel metal2 s 15750 0 15806 600 6 HI[254]
port 172 nsew signal output
rlabel metal2 s 14922 0 14978 600 6 HI[255]
port 173 nsew signal output
rlabel metal2 s 38382 0 38438 600 6 HI[256]
port 174 nsew signal output
rlabel metal2 s 27342 0 27398 600 6 HI[257]
port 175 nsew signal output
rlabel metal2 s 16302 0 16358 600 6 HI[258]
port 176 nsew signal output
rlabel metal2 s 38658 0 38714 600 6 HI[259]
port 177 nsew signal output
rlabel metal2 s 16578 0 16634 600 6 HI[25]
port 178 nsew signal output
rlabel metal2 s 1950 0 2006 600 6 HI[260]
port 179 nsew signal output
rlabel metal2 s 38934 0 38990 600 6 HI[261]
port 180 nsew signal output
rlabel metal2 s 1674 0 1730 600 6 HI[262]
port 181 nsew signal output
rlabel metal2 s 17130 0 17186 600 6 HI[263]
port 182 nsew signal output
rlabel metal2 s 14370 0 14426 600 6 HI[264]
port 183 nsew signal output
rlabel metal2 s 48870 0 48926 600 6 HI[265]
port 184 nsew signal output
rlabel metal2 s 28170 0 28226 600 6 HI[266]
port 185 nsew signal output
rlabel metal2 s 17682 0 17738 600 6 HI[267]
port 186 nsew signal output
rlabel metal2 s 42522 0 42578 600 6 HI[268]
port 187 nsew signal output
rlabel metal2 s 39486 0 39542 600 6 HI[269]
port 188 nsew signal output
rlabel metal2 s 6642 0 6698 600 6 HI[26]
port 189 nsew signal output
rlabel metal2 s 18234 0 18290 600 6 HI[270]
port 190 nsew signal output
rlabel metal2 s 7194 0 7250 600 6 HI[271]
port 191 nsew signal output
rlabel metal2 s 39762 0 39818 600 6 HI[272]
port 192 nsew signal output
rlabel metal2 s 10506 0 10562 600 6 HI[273]
port 193 nsew signal output
rlabel metal2 s 24306 0 24362 600 6 HI[274]
port 194 nsew signal output
rlabel metal2 s 49146 0 49202 600 6 HI[275]
port 195 nsew signal output
rlabel metal2 s 40038 0 40094 600 6 HI[276]
port 196 nsew signal output
rlabel metal2 s 5262 0 5318 600 6 HI[277]
port 197 nsew signal output
rlabel metal2 s 19338 0 19394 600 6 HI[278]
port 198 nsew signal output
rlabel metal2 s 29274 0 29330 600 6 HI[279]
port 199 nsew signal output
rlabel metal2 s 40314 0 40370 600 6 HI[27]
port 200 nsew signal output
rlabel metal2 s 3054 0 3110 600 6 HI[280]
port 201 nsew signal output
rlabel metal2 s 49422 0 49478 600 6 HI[281]
port 202 nsew signal output
rlabel metal2 s 6918 0 6974 600 6 HI[282]
port 203 nsew signal output
rlabel metal2 s 40590 0 40646 600 6 HI[283]
port 204 nsew signal output
rlabel metal2 s 1398 0 1454 600 6 HI[284]
port 205 nsew signal output
rlabel metal2 s 20442 0 20498 600 6 HI[285]
port 206 nsew signal output
rlabel metal2 s 32034 0 32090 600 6 HI[286]
port 207 nsew signal output
rlabel metal2 s 40866 0 40922 600 6 HI[287]
port 208 nsew signal output
rlabel metal2 s 3330 0 3386 600 6 HI[288]
port 209 nsew signal output
rlabel metal2 s 30102 0 30158 600 6 HI[289]
port 210 nsew signal output
rlabel metal2 s 3882 0 3938 600 6 HI[28]
port 211 nsew signal output
rlabel metal2 s 41142 0 41198 600 6 HI[290]
port 212 nsew signal output
rlabel metal2 s 4710 0 4766 600 6 HI[291]
port 213 nsew signal output
rlabel metal2 s 21546 0 21602 600 6 HI[292]
port 214 nsew signal output
rlabel metal2 s 9678 0 9734 600 6 HI[293]
port 215 nsew signal output
rlabel metal2 s 41418 0 41474 600 6 HI[294]
port 216 nsew signal output
rlabel metal2 s 49698 0 49754 600 6 HI[295]
port 217 nsew signal output
rlabel metal2 s 30654 0 30710 600 6 HI[296]
port 218 nsew signal output
rlabel metal2 s 2502 0 2558 600 6 HI[297]
port 219 nsew signal output
rlabel metal2 s 41694 0 41750 600 6 HI[298]
port 220 nsew signal output
rlabel metal2 s 33690 0 33746 600 6 HI[299]
port 221 nsew signal output
rlabel metal2 s 22650 0 22706 600 6 HI[29]
port 222 nsew signal output
rlabel metal2 s 4158 0 4214 600 6 HI[2]
port 223 nsew signal output
rlabel metal2 s 41970 0 42026 600 6 HI[300]
port 224 nsew signal output
rlabel metal2 s 49974 0 50030 600 6 HI[301]
port 225 nsew signal output
rlabel metal2 s 23202 0 23258 600 6 HI[302]
port 226 nsew signal output
rlabel metal2 s 13542 0 13598 600 6 HI[303]
port 227 nsew signal output
rlabel metal2 s 42246 0 42302 600 6 HI[304]
port 228 nsew signal output
rlabel metal2 s 27618 0 27674 600 6 HI[305]
port 229 nsew signal output
rlabel metal2 s 50250 0 50306 600 6 HI[306]
port 230 nsew signal output
rlabel metal2 s 53286 0 53342 600 6 HI[307]
port 231 nsew signal output
rlabel metal2 s 54390 0 54446 600 6 HI[308]
port 232 nsew signal output
rlabel metal2 s 43074 0 43130 600 6 HI[309]
port 233 nsew signal output
rlabel metal2 s 31758 0 31814 600 6 HI[30]
port 234 nsew signal output
rlabel metal2 s 12438 0 12494 600 6 HI[310]
port 235 nsew signal output
rlabel metal2 s 42798 0 42854 600 6 HI[311]
port 236 nsew signal output
rlabel metal2 s 15198 0 15254 600 6 HI[312]
port 237 nsew signal output
rlabel metal2 s 43626 0 43682 600 6 HI[313]
port 238 nsew signal output
rlabel metal2 s 50526 0 50582 600 6 HI[314]
port 239 nsew signal output
rlabel metal2 s 44730 0 44786 600 6 HI[315]
port 240 nsew signal output
rlabel metal2 s 15474 0 15530 600 6 HI[316]
port 241 nsew signal output
rlabel metal2 s 25410 0 25466 600 6 HI[317]
port 242 nsew signal output
rlabel metal2 s 19890 0 19946 600 6 HI[318]
port 243 nsew signal output
rlabel metal2 s 43350 0 43406 600 6 HI[319]
port 244 nsew signal output
rlabel metal2 s 570 0 626 600 6 HI[31]
port 245 nsew signal output
rlabel metal2 s 25962 0 26018 600 6 HI[320]
port 246 nsew signal output
rlabel metal2 s 1122 0 1178 600 6 HI[321]
port 247 nsew signal output
rlabel metal2 s 45834 0 45890 600 6 HI[322]
port 248 nsew signal output
rlabel metal2 s 50802 0 50858 600 6 HI[323]
port 249 nsew signal output
rlabel metal2 s 26514 0 26570 600 6 HI[324]
port 250 nsew signal output
rlabel metal2 s 16026 0 16082 600 6 HI[325]
port 251 nsew signal output
rlabel metal2 s 43902 0 43958 600 6 HI[326]
port 252 nsew signal output
rlabel metal2 s 3606 0 3662 600 6 HI[327]
port 253 nsew signal output
rlabel metal2 s 27066 0 27122 600 6 HI[328]
port 254 nsew signal output
rlabel metal2 s 8022 0 8078 600 6 HI[329]
port 255 nsew signal output
rlabel metal2 s 44178 0 44234 600 6 HI[32]
port 256 nsew signal output
rlabel metal2 s 5814 0 5870 600 6 HI[330]
port 257 nsew signal output
rlabel metal2 s 53562 0 53618 600 6 HI[331]
port 258 nsew signal output
rlabel metal2 s 18786 0 18842 600 6 HI[332]
port 259 nsew signal output
rlabel metal2 s 44454 0 44510 600 6 HI[333]
port 260 nsew signal output
rlabel metal2 s 27894 0 27950 600 6 HI[334]
port 261 nsew signal output
rlabel metal2 s 9954 0 10010 600 6 HI[335]
port 262 nsew signal output
rlabel metal2 s 9402 0 9458 600 6 HI[336]
port 263 nsew signal output
rlabel metal2 s 51078 0 51134 600 6 HI[337]
port 264 nsew signal output
rlabel metal2 s 19614 0 19670 600 6 HI[338]
port 265 nsew signal output
rlabel metal2 s 17406 0 17462 600 6 HI[339]
port 266 nsew signal output
rlabel metal2 s 28446 0 28502 600 6 HI[33]
port 267 nsew signal output
rlabel metal2 s 11610 0 11666 600 6 HI[340]
port 268 nsew signal output
rlabel metal2 s 53838 0 53894 600 6 HI[341]
port 269 nsew signal output
rlabel metal2 s 45006 0 45062 600 6 HI[342]
port 270 nsew signal output
rlabel metal2 s 67914 3800 67970 4400 6 HI[343]
port 271 nsew signal output
rlabel metal2 s 14922 3800 14978 4400 6 HI[344]
port 272 nsew signal output
rlabel metal2 s 15198 3800 15254 4400 6 HI[345]
port 273 nsew signal output
rlabel metal2 s 15474 3800 15530 4400 6 HI[346]
port 274 nsew signal output
rlabel metal2 s 15750 3800 15806 4400 6 HI[347]
port 275 nsew signal output
rlabel metal2 s 16026 3800 16082 4400 6 HI[348]
port 276 nsew signal output
rlabel metal2 s 16302 3800 16358 4400 6 HI[349]
port 277 nsew signal output
rlabel metal2 s 16578 3800 16634 4400 6 HI[34]
port 278 nsew signal output
rlabel metal2 s 16854 3800 16910 4400 6 HI[350]
port 279 nsew signal output
rlabel metal2 s 17130 3800 17186 4400 6 HI[351]
port 280 nsew signal output
rlabel metal2 s 17406 3800 17462 4400 6 HI[352]
port 281 nsew signal output
rlabel metal2 s 17682 3800 17738 4400 6 HI[353]
port 282 nsew signal output
rlabel metal2 s 17958 3800 18014 4400 6 HI[354]
port 283 nsew signal output
rlabel metal2 s 18234 3800 18290 4400 6 HI[355]
port 284 nsew signal output
rlabel metal2 s 18510 3800 18566 4400 6 HI[356]
port 285 nsew signal output
rlabel metal2 s 18786 3800 18842 4400 6 HI[357]
port 286 nsew signal output
rlabel metal2 s 19062 3800 19118 4400 6 HI[358]
port 287 nsew signal output
rlabel metal2 s 19338 3800 19394 4400 6 HI[359]
port 288 nsew signal output
rlabel metal2 s 19614 3800 19670 4400 6 HI[35]
port 289 nsew signal output
rlabel metal2 s 19890 3800 19946 4400 6 HI[360]
port 290 nsew signal output
rlabel metal2 s 20166 3800 20222 4400 6 HI[361]
port 291 nsew signal output
rlabel metal2 s 20442 3800 20498 4400 6 HI[362]
port 292 nsew signal output
rlabel metal2 s 20718 3800 20774 4400 6 HI[363]
port 293 nsew signal output
rlabel metal2 s 20994 3800 21050 4400 6 HI[364]
port 294 nsew signal output
rlabel metal2 s 21270 3800 21326 4400 6 HI[365]
port 295 nsew signal output
rlabel metal2 s 21546 3800 21602 4400 6 HI[366]
port 296 nsew signal output
rlabel metal2 s 21822 3800 21878 4400 6 HI[367]
port 297 nsew signal output
rlabel metal2 s 22098 3800 22154 4400 6 HI[368]
port 298 nsew signal output
rlabel metal2 s 22374 3800 22430 4400 6 HI[369]
port 299 nsew signal output
rlabel metal2 s 22650 3800 22706 4400 6 HI[36]
port 300 nsew signal output
rlabel metal2 s 22926 3800 22982 4400 6 HI[370]
port 301 nsew signal output
rlabel metal2 s 23202 3800 23258 4400 6 HI[371]
port 302 nsew signal output
rlabel metal2 s 23478 3800 23534 4400 6 HI[372]
port 303 nsew signal output
rlabel metal2 s 23754 3800 23810 4400 6 HI[373]
port 304 nsew signal output
rlabel metal2 s 24030 3800 24086 4400 6 HI[374]
port 305 nsew signal output
rlabel metal2 s 24306 3800 24362 4400 6 HI[375]
port 306 nsew signal output
rlabel metal2 s 24582 3800 24638 4400 6 HI[376]
port 307 nsew signal output
rlabel metal2 s 24858 3800 24914 4400 6 HI[377]
port 308 nsew signal output
rlabel metal2 s 25134 3800 25190 4400 6 HI[378]
port 309 nsew signal output
rlabel metal2 s 25410 3800 25466 4400 6 HI[379]
port 310 nsew signal output
rlabel metal2 s 25686 3800 25742 4400 6 HI[37]
port 311 nsew signal output
rlabel metal2 s 25962 3800 26018 4400 6 HI[380]
port 312 nsew signal output
rlabel metal2 s 26238 3800 26294 4400 6 HI[381]
port 313 nsew signal output
rlabel metal2 s 26514 3800 26570 4400 6 HI[382]
port 314 nsew signal output
rlabel metal2 s 26790 3800 26846 4400 6 HI[383]
port 315 nsew signal output
rlabel metal2 s 27066 3800 27122 4400 6 HI[384]
port 316 nsew signal output
rlabel metal2 s 27342 3800 27398 4400 6 HI[385]
port 317 nsew signal output
rlabel metal2 s 27618 3800 27674 4400 6 HI[386]
port 318 nsew signal output
rlabel metal2 s 27894 3800 27950 4400 6 HI[387]
port 319 nsew signal output
rlabel metal2 s 28170 3800 28226 4400 6 HI[388]
port 320 nsew signal output
rlabel metal2 s 28446 3800 28502 4400 6 HI[389]
port 321 nsew signal output
rlabel metal2 s 28722 3800 28778 4400 6 HI[38]
port 322 nsew signal output
rlabel metal2 s 28998 3800 29054 4400 6 HI[390]
port 323 nsew signal output
rlabel metal2 s 29274 3800 29330 4400 6 HI[391]
port 324 nsew signal output
rlabel metal2 s 29550 3800 29606 4400 6 HI[392]
port 325 nsew signal output
rlabel metal2 s 29826 3800 29882 4400 6 HI[393]
port 326 nsew signal output
rlabel metal2 s 30102 3800 30158 4400 6 HI[394]
port 327 nsew signal output
rlabel metal2 s 30378 3800 30434 4400 6 HI[395]
port 328 nsew signal output
rlabel metal2 s 30654 3800 30710 4400 6 HI[396]
port 329 nsew signal output
rlabel metal2 s 30930 3800 30986 4400 6 HI[397]
port 330 nsew signal output
rlabel metal2 s 31206 3800 31262 4400 6 HI[398]
port 331 nsew signal output
rlabel metal2 s 31482 3800 31538 4400 6 HI[399]
port 332 nsew signal output
rlabel metal2 s 31758 3800 31814 4400 6 HI[39]
port 333 nsew signal output
rlabel metal2 s 32034 3800 32090 4400 6 HI[3]
port 334 nsew signal output
rlabel metal2 s 32310 3800 32366 4400 6 HI[400]
port 335 nsew signal output
rlabel metal2 s 32586 3800 32642 4400 6 HI[401]
port 336 nsew signal output
rlabel metal2 s 32862 3800 32918 4400 6 HI[402]
port 337 nsew signal output
rlabel metal2 s 33138 3800 33194 4400 6 HI[403]
port 338 nsew signal output
rlabel metal2 s 33414 3800 33470 4400 6 HI[404]
port 339 nsew signal output
rlabel metal2 s 33690 3800 33746 4400 6 HI[405]
port 340 nsew signal output
rlabel metal2 s 33966 3800 34022 4400 6 HI[406]
port 341 nsew signal output
rlabel metal2 s 34242 3800 34298 4400 6 HI[407]
port 342 nsew signal output
rlabel metal2 s 34518 3800 34574 4400 6 HI[408]
port 343 nsew signal output
rlabel metal2 s 34794 3800 34850 4400 6 HI[409]
port 344 nsew signal output
rlabel metal2 s 35070 3800 35126 4400 6 HI[40]
port 345 nsew signal output
rlabel metal2 s 35346 3800 35402 4400 6 HI[410]
port 346 nsew signal output
rlabel metal2 s 35622 3800 35678 4400 6 HI[411]
port 347 nsew signal output
rlabel metal2 s 35898 3800 35954 4400 6 HI[412]
port 348 nsew signal output
rlabel metal2 s 36174 3800 36230 4400 6 HI[413]
port 349 nsew signal output
rlabel metal2 s 36450 3800 36506 4400 6 HI[414]
port 350 nsew signal output
rlabel metal2 s 36726 3800 36782 4400 6 HI[415]
port 351 nsew signal output
rlabel metal2 s 37002 3800 37058 4400 6 HI[416]
port 352 nsew signal output
rlabel metal2 s 37278 3800 37334 4400 6 HI[417]
port 353 nsew signal output
rlabel metal2 s 37554 3800 37610 4400 6 HI[418]
port 354 nsew signal output
rlabel metal2 s 37830 3800 37886 4400 6 HI[419]
port 355 nsew signal output
rlabel metal2 s 38106 3800 38162 4400 6 HI[41]
port 356 nsew signal output
rlabel metal2 s 38382 3800 38438 4400 6 HI[420]
port 357 nsew signal output
rlabel metal2 s 38658 3800 38714 4400 6 HI[421]
port 358 nsew signal output
rlabel metal2 s 38934 3800 38990 4400 6 HI[422]
port 359 nsew signal output
rlabel metal2 s 39210 3800 39266 4400 6 HI[423]
port 360 nsew signal output
rlabel metal2 s 39486 3800 39542 4400 6 HI[424]
port 361 nsew signal output
rlabel metal2 s 39762 3800 39818 4400 6 HI[425]
port 362 nsew signal output
rlabel metal2 s 40038 3800 40094 4400 6 HI[426]
port 363 nsew signal output
rlabel metal2 s 40314 3800 40370 4400 6 HI[427]
port 364 nsew signal output
rlabel metal2 s 40590 3800 40646 4400 6 HI[428]
port 365 nsew signal output
rlabel metal2 s 40866 3800 40922 4400 6 HI[429]
port 366 nsew signal output
rlabel metal2 s 41142 3800 41198 4400 6 HI[42]
port 367 nsew signal output
rlabel metal2 s 41418 3800 41474 4400 6 HI[430]
port 368 nsew signal output
rlabel metal2 s 41694 3800 41750 4400 6 HI[431]
port 369 nsew signal output
rlabel metal2 s 41970 3800 42026 4400 6 HI[432]
port 370 nsew signal output
rlabel metal2 s 42246 3800 42302 4400 6 HI[433]
port 371 nsew signal output
rlabel metal2 s 42522 3800 42578 4400 6 HI[434]
port 372 nsew signal output
rlabel metal2 s 42798 3800 42854 4400 6 HI[435]
port 373 nsew signal output
rlabel metal2 s 43074 3800 43130 4400 6 HI[436]
port 374 nsew signal output
rlabel metal2 s 43350 3800 43406 4400 6 HI[437]
port 375 nsew signal output
rlabel metal2 s 43626 3800 43682 4400 6 HI[438]
port 376 nsew signal output
rlabel metal2 s 43902 3800 43958 4400 6 HI[439]
port 377 nsew signal output
rlabel metal2 s 44178 3800 44234 4400 6 HI[43]
port 378 nsew signal output
rlabel metal2 s 44454 3800 44510 4400 6 HI[440]
port 379 nsew signal output
rlabel metal2 s 44730 3800 44786 4400 6 HI[441]
port 380 nsew signal output
rlabel metal2 s 45006 3800 45062 4400 6 HI[442]
port 381 nsew signal output
rlabel metal2 s 45282 3800 45338 4400 6 HI[443]
port 382 nsew signal output
rlabel metal2 s 45558 3800 45614 4400 6 HI[444]
port 383 nsew signal output
rlabel metal2 s 45834 3800 45890 4400 6 HI[445]
port 384 nsew signal output
rlabel metal2 s 46110 3800 46166 4400 6 HI[446]
port 385 nsew signal output
rlabel metal2 s 46386 3800 46442 4400 6 HI[447]
port 386 nsew signal output
rlabel metal2 s 46662 3800 46718 4400 6 HI[448]
port 387 nsew signal output
rlabel metal2 s 46938 3800 46994 4400 6 HI[449]
port 388 nsew signal output
rlabel metal2 s 47214 3800 47270 4400 6 HI[44]
port 389 nsew signal output
rlabel metal2 s 47490 3800 47546 4400 6 HI[450]
port 390 nsew signal output
rlabel metal2 s 47766 3800 47822 4400 6 HI[451]
port 391 nsew signal output
rlabel metal2 s 48042 3800 48098 4400 6 HI[452]
port 392 nsew signal output
rlabel metal2 s 48318 3800 48374 4400 6 HI[453]
port 393 nsew signal output
rlabel metal2 s 48594 3800 48650 4400 6 HI[454]
port 394 nsew signal output
rlabel metal2 s 48870 3800 48926 4400 6 HI[455]
port 395 nsew signal output
rlabel metal2 s 49146 3800 49202 4400 6 HI[456]
port 396 nsew signal output
rlabel metal2 s 49422 3800 49478 4400 6 HI[457]
port 397 nsew signal output
rlabel metal2 s 49698 3800 49754 4400 6 HI[458]
port 398 nsew signal output
rlabel metal2 s 49974 3800 50030 4400 6 HI[459]
port 399 nsew signal output
rlabel metal2 s 50250 3800 50306 4400 6 HI[45]
port 400 nsew signal output
rlabel metal2 s 50526 3800 50582 4400 6 HI[460]
port 401 nsew signal output
rlabel metal2 s 50802 3800 50858 4400 6 HI[461]
port 402 nsew signal output
rlabel metal2 s 51078 3800 51134 4400 6 HI[462]
port 403 nsew signal output
rlabel metal2 s 51354 3800 51410 4400 6 HI[46]
port 404 nsew signal output
rlabel metal2 s 51630 3800 51686 4400 6 HI[47]
port 405 nsew signal output
rlabel metal2 s 51906 3800 51962 4400 6 HI[48]
port 406 nsew signal output
rlabel metal2 s 52182 3800 52238 4400 6 HI[49]
port 407 nsew signal output
rlabel metal2 s 52458 3800 52514 4400 6 HI[4]
port 408 nsew signal output
rlabel metal2 s 52734 3800 52790 4400 6 HI[50]
port 409 nsew signal output
rlabel metal2 s 53010 3800 53066 4400 6 HI[51]
port 410 nsew signal output
rlabel metal2 s 53286 3800 53342 4400 6 HI[52]
port 411 nsew signal output
rlabel metal2 s 53562 3800 53618 4400 6 HI[53]
port 412 nsew signal output
rlabel metal2 s 53838 3800 53894 4400 6 HI[54]
port 413 nsew signal output
rlabel metal2 s 54114 3800 54170 4400 6 HI[55]
port 414 nsew signal output
rlabel metal2 s 54390 3800 54446 4400 6 HI[56]
port 415 nsew signal output
rlabel metal2 s 54666 3800 54722 4400 6 HI[57]
port 416 nsew signal output
rlabel metal2 s 54942 3800 54998 4400 6 HI[58]
port 417 nsew signal output
rlabel metal2 s 55218 3800 55274 4400 6 HI[59]
port 418 nsew signal output
rlabel metal2 s 55494 3800 55550 4400 6 HI[5]
port 419 nsew signal output
rlabel metal2 s 55770 3800 55826 4400 6 HI[60]
port 420 nsew signal output
rlabel metal2 s 56046 3800 56102 4400 6 HI[61]
port 421 nsew signal output
rlabel metal2 s 56322 3800 56378 4400 6 HI[62]
port 422 nsew signal output
rlabel metal2 s 56598 3800 56654 4400 6 HI[63]
port 423 nsew signal output
rlabel metal2 s 56874 3800 56930 4400 6 HI[64]
port 424 nsew signal output
rlabel metal2 s 57150 3800 57206 4400 6 HI[65]
port 425 nsew signal output
rlabel metal2 s 57426 3800 57482 4400 6 HI[66]
port 426 nsew signal output
rlabel metal2 s 57702 3800 57758 4400 6 HI[67]
port 427 nsew signal output
rlabel metal2 s 57978 3800 58034 4400 6 HI[68]
port 428 nsew signal output
rlabel metal2 s 58254 3800 58310 4400 6 HI[69]
port 429 nsew signal output
rlabel metal2 s 58530 3800 58586 4400 6 HI[6]
port 430 nsew signal output
rlabel metal2 s 58806 3800 58862 4400 6 HI[70]
port 431 nsew signal output
rlabel metal2 s 59082 3800 59138 4400 6 HI[71]
port 432 nsew signal output
rlabel metal2 s 59358 3800 59414 4400 6 HI[72]
port 433 nsew signal output
rlabel metal2 s 59634 3800 59690 4400 6 HI[73]
port 434 nsew signal output
rlabel metal2 s 59910 3800 59966 4400 6 HI[74]
port 435 nsew signal output
rlabel metal2 s 60186 3800 60242 4400 6 HI[75]
port 436 nsew signal output
rlabel metal2 s 60462 3800 60518 4400 6 HI[76]
port 437 nsew signal output
rlabel metal2 s 60738 3800 60794 4400 6 HI[77]
port 438 nsew signal output
rlabel metal2 s 61014 3800 61070 4400 6 HI[78]
port 439 nsew signal output
rlabel metal2 s 61290 3800 61346 4400 6 HI[79]
port 440 nsew signal output
rlabel metal2 s 61566 3800 61622 4400 6 HI[7]
port 441 nsew signal output
rlabel metal2 s 61842 3800 61898 4400 6 HI[80]
port 442 nsew signal output
rlabel metal2 s 62118 3800 62174 4400 6 HI[81]
port 443 nsew signal output
rlabel metal2 s 62394 3800 62450 4400 6 HI[82]
port 444 nsew signal output
rlabel metal2 s 62670 3800 62726 4400 6 HI[83]
port 445 nsew signal output
rlabel metal2 s 62946 3800 63002 4400 6 HI[84]
port 446 nsew signal output
rlabel metal2 s 63222 3800 63278 4400 6 HI[85]
port 447 nsew signal output
rlabel metal2 s 63498 3800 63554 4400 6 HI[86]
port 448 nsew signal output
rlabel metal2 s 63774 3800 63830 4400 6 HI[87]
port 449 nsew signal output
rlabel metal2 s 64050 3800 64106 4400 6 HI[88]
port 450 nsew signal output
rlabel metal2 s 64326 3800 64382 4400 6 HI[89]
port 451 nsew signal output
rlabel metal2 s 64602 3800 64658 4400 6 HI[8]
port 452 nsew signal output
rlabel metal2 s 64878 3800 64934 4400 6 HI[90]
port 453 nsew signal output
rlabel metal2 s 65154 3800 65210 4400 6 HI[91]
port 454 nsew signal output
rlabel metal2 s 65430 3800 65486 4400 6 HI[92]
port 455 nsew signal output
rlabel metal2 s 65706 3800 65762 4400 6 HI[93]
port 456 nsew signal output
rlabel metal2 s 65982 3800 66038 4400 6 HI[94]
port 457 nsew signal output
rlabel metal2 s 66258 3800 66314 4400 6 HI[95]
port 458 nsew signal output
rlabel metal2 s 66534 3800 66590 4400 6 HI[96]
port 459 nsew signal output
rlabel metal2 s 66810 3800 66866 4400 6 HI[97]
port 460 nsew signal output
rlabel metal2 s 67086 3800 67142 4400 6 HI[98]
port 461 nsew signal output
rlabel metal2 s 67362 3800 67418 4400 6 HI[99]
port 462 nsew signal output
rlabel metal2 s 67638 3800 67694 4400 6 HI[9]
port 463 nsew signal output
rlabel metal3 s 1288 1190 68816 1290 6 vccd1
port 464 nsew power input
rlabel metal2 s 7238 1040 7338 3312 6 vccd1
port 464 nsew power input
rlabel metal2 s 19238 1040 19338 3312 6 vccd1
port 464 nsew power input
rlabel metal2 s 31238 1040 31338 3312 6 vccd1
port 464 nsew power input
rlabel metal2 s 43238 1040 43338 3312 6 vccd1
port 464 nsew power input
rlabel metal2 s 55238 1040 55338 3312 6 vccd1
port 464 nsew power input
rlabel metal2 s 67238 1040 67338 3312 6 vccd1
port 464 nsew power input
rlabel metal3 s 1288 2270 68816 2370 6 vssd1
port 465 nsew ground input
rlabel metal2 s 13238 1040 13338 3312 6 vssd1
port 465 nsew ground input
rlabel metal2 s 25238 1040 25338 3312 6 vssd1
port 465 nsew ground input
rlabel metal2 s 37238 1040 37338 3312 6 vssd1
port 465 nsew ground input
rlabel metal2 s 49238 1040 49338 3312 6 vssd1
port 465 nsew ground input
rlabel metal2 s 61238 1040 61338 3312 6 vssd1
port 465 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 70000 4400
string LEFview TRUE
string GDS_FILE /project/openlane/mprj_logic_high/runs/mprj_logic_high/results/magic/mprj_logic_high.gds
string GDS_END 514418
string GDS_START 24116
<< end >>

