* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_2 abstract view
.subckt sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_4 abstract view
.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_67_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6914_ _6967_/CLK _6914_/D fanout586/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6845_ _6889_/CLK _6845_/D fanout582/X VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6776_ _6780_/CLK _6776_/D fanout575/X VGND VGND VPWR VPWR _6776_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3988_ _6549_/A0 hold955/X _3992_/S VGND VGND VPWR VPWR _3988_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5727_ _5726_/Y _5759_/B _5712_/Y VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5658_ _5667_/A0 _5658_/A1 _5665_/S VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4609_ _4620_/A _4595_/A _4786_/B _4923_/B _4333_/A VGND VGND VPWR VPWR _5216_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ _3924_/B hold266/X hold44/X VGND VGND VPWR VPWR _5589_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold340 _7066_/Q VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold351 _3908_/X VGND VGND VPWR VPWR _6587_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 hold362/A VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _7034_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _6547_/X VGND VGND VPWR VPWR _7274_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _5436_/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7259_ _7259_/CLK _7259_/D fanout613/X VGND VGND VPWR VPWR _7259_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1040 _6533_/X VGND VGND VPWR VPWR _7262_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1051 _5538_/X VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _3980_/X VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1073 _6687_/Q VGND VGND VPWR VPWR _4034_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _4097_/X VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1095 _6725_/Q VGND VGND VPWR VPWR _4095_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_202 _6465_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _6543_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_224 _3922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _3340_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 hold67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 _3508_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 _3918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4960_ _4629_/Y _4951_/X _4958_/X _4959_/X VGND VGND VPWR VPWR _4960_/X sky130_fd_sc_hd__o211a_1
X_3911_ hold24/X hold200/X _3912_/S VGND VGND VPWR VPWR _3911_/X sky130_fd_sc_hd__mux2_1
X_4891_ _5089_/C _4308_/D _4480_/B _4890_/Y VGND VGND VPWR VPWR _4891_/X sky130_fd_sc_hd__a31o_1
X_6630_ _7218_/CLK _6630_/D VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfxtp_1
X_3842_ _6956_/Q _3424_/X _3571_/X hold94/A _3841_/X VGND VGND VPWR VPWR _3843_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6561_ _6761_/CLK _6561_/D _3291_/A VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfstp_2
X_3773_ _7035_/Q _3547_/X _3558_/X _6611_/Q _3772_/X VGND VGND VPWR VPWR _3773_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5512_ _6548_/B _5512_/B _5675_/D _5657_/D VGND VGND VPWR VPWR _5520_/S sky130_fd_sc_hd__nand4_4
X_6492_ _7257_/Q _6492_/A2 _6492_/B1 _4164_/Y _6491_/X VGND VGND VPWR VPWR _6492_/X
+ sky130_fd_sc_hd__a221o_1
X_5443_ hold307/X _3919_/C _5448_/S VGND VGND VPWR VPWR _5443_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5374_ hold170/X hold83/X _5376_/S VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__mux2_1
X_7113_ _7245_/CLK _7113_/D fanout599/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_2
X_4325_ _4691_/B _4254_/Y _4304_/Y _4870_/B _4320_/Y VGND VGND VPWR VPWR _4325_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7044_ _7120_/CLK _7044_/D fanout606/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_1
X_4256_ _4870_/B _4247_/Y _4429_/D VGND VGND VPWR VPWR _4256_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4187_ hold174/X _4053_/X _4187_/S VGND VGND VPWR VPWR _4187_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6828_ _6828_/CLK _6828_/D fanout583/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6759_ _7260_/CLK _6759_/D fanout572/X VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold170 _6892_/Q VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _5401_/X VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _7148_/Q VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4110_ hold21/X hold206/X _4111_/S VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__mux2_1
X_5090_ _5090_/A _5090_/B _5263_/B VGND VGND VPWR VPWR _5090_/X sky130_fd_sc_hd__and3_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4041_ _4055_/A1 _6898_/Q _3346_/D hold64/X _5494_/A VGND VGND VPWR VPWR _5341_/C
+ sky130_fd_sc_hd__o311a_4
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5992_ _6768_/Q _5776_/X _5991_/X _6025_/B _5990_/X VGND VGND VPWR VPWR _5992_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_92_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4943_ _4939_/A _4682_/B _4678_/A _4942_/X VGND VGND VPWR VPWR _4954_/D sky130_fd_sc_hd__a211o_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4874_ _4859_/C _5255_/A _5255_/C _4687_/B _4718_/D VGND VGND VPWR VPWR _4874_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_33_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6613_ _7251_/CLK _6613_/D VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfxtp_1
X_3825_ _3825_/A _3825_/B _3825_/C _3825_/D VGND VGND VPWR VPWR _3825_/Y sky130_fd_sc_hd__nor4_1
XFILLER_165_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6544_ _6550_/A0 hold820/X _6547_/S VGND VGND VPWR VPWR _6544_/X sky130_fd_sc_hd__mux2_1
X_3756_ _6815_/Q _5341_/A _5485_/B _3496_/X _6995_/Q VGND VGND VPWR VPWR _3756_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_192_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6475_ _3693_/Y _6475_/A1 _6480_/S VGND VGND VPWR VPWR _7223_/D sky130_fd_sc_hd__mux2_1
X_3687_ _6599_/Q _6530_/C _3466_/X _5593_/B _7089_/Q VGND VGND VPWR VPWR _3687_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5426_ _5430_/S hold846/X _3433_/X _3922_/X VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__a22o_1
Xoutput220 _7293_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput231 _7303_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput242 _7283_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
Xoutput253 _7311_/X VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput264 _6820_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5357_ hold21/X hold242/X _5358_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
Xoutput275 hold94/A VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
XFILLER_102_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput286 _6836_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xoutput297 _6838_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
XFILLER_87_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4308_ _4647_/C _4310_/B _4310_/C _4308_/D VGND VGND VPWR VPWR _4308_/Y sky130_fd_sc_hd__nand4_2
X_5288_ _6524_/A _6536_/B _5327_/D _6536_/D VGND VGND VPWR VPWR _5294_/S sky130_fd_sc_hd__and4_2
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7027_ _7167_/CLK _7027_/D fanout604/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4239_ _4637_/A _4747_/A VGND VGND VPWR VPWR _4734_/B sky130_fd_sc_hd__and2b_1
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire347 _6158_/Y VGND VGND VPWR VPWR wire347/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire358 _5125_/C VGND VGND VPWR VPWR wire358/X sky130_fd_sc_hd__clkbuf_1
Xwire369 _5969_/Y VGND VGND VPWR VPWR _5974_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_183_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout480 hold72/X VGND VGND VPWR VPWR _6548_/C sky130_fd_sc_hd__buf_12
Xfanout491 hold17/X VGND VGND VPWR VPWR _6548_/A sky130_fd_sc_hd__buf_12
XFILLER_65_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3610_ _6734_/Q _5341_/A _3721_/A3 _3607_/X _3609_/X VGND VGND VPWR VPWR _3610_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_174_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4590_ _4815_/A _4606_/B _4923_/A _4606_/D VGND VGND VPWR VPWR _4591_/B sky130_fd_sc_hd__and4_1
XFILLER_190_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3541_ _7039_/Q _3538_/X _3539_/X input52/X _3537_/X VGND VGND VPWR VPWR _3541_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold906 _5529_/X VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 _6919_/Q VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 _5547_/X VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 _4028_/X VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6260_ _7059_/Q _5732_/X _6108_/X _6454_/B1 _6955_/Q VGND VGND VPWR VPWR _6260_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_182_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3472_ _6855_/Q _5327_/D _3902_/A3 _3471_/X input20/X VGND VGND VPWR VPWR _3472_/X
+ sky130_fd_sc_hd__a32o_1
X_5211_ _5210_/X _4726_/Y _5064_/X _5085_/X VGND VGND VPWR VPWR _5211_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6191_ wire357/X _6190_/Y _6872_/Q _6466_/A1 VGND VGND VPWR VPWR _6191_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5142_ _5141_/X _5142_/B _5261_/C _5142_/D VGND VGND VPWR VPWR _5145_/B sky130_fd_sc_hd__nand4b_1
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5073_ _5070_/X _5073_/B _5270_/C VGND VGND VPWR VPWR _5073_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_111_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4024_ _4024_/A0 _4152_/B _4028_/S VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5975_ _6878_/Q _5726_/Y _5963_/X _5974_/Y _3246_/Y VGND VGND VPWR VPWR _5975_/X
+ sky130_fd_sc_hd__o221a_2
X_4926_ _5040_/C _4527_/X _4567_/Y _4707_/Y _4552_/Y VGND VGND VPWR VPWR _5100_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_100_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4857_ _4859_/C _5255_/A _4857_/C VGND VGND VPWR VPWR _4857_/X sky130_fd_sc_hd__and3_1
XFILLER_178_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3808_ input30/X _3466_/X _5311_/C _3807_/X _3805_/X VGND VGND VPWR VPWR _3808_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4788_ _4788_/A _5263_/B _4945_/C VGND VGND VPWR VPWR _4788_/X sky130_fd_sc_hd__and3_1
XFILLER_181_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6527_ _3919_/C hold404/X _6529_/S VGND VGND VPWR VPWR _6527_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ input23/X _3471_/X _5404_/B _6922_/Q _3695_/X VGND VGND VPWR VPWR _3739_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_109_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6458_ _6687_/Q _6101_/X _6448_/X _6450_/X _6457_/X VGND VGND VPWR VPWR _6458_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_133_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5409_ _5404_/B _3925_/X _5412_/S hold895/X VGND VGND VPWR VPWR _5409_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6389_ _6389_/A _6389_/B _6389_/C _6440_/D VGND VGND VPWR VPWR _6390_/D sky130_fd_sc_hd__nor4_1
XFILLER_102_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5760_ _6292_/S _3307_/B _5759_/X VGND VGND VPWR VPWR _6343_/S sky130_fd_sc_hd__a21oi_4
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ _4711_/A _4711_/B _4711_/C VGND VGND VPWR VPWR _4717_/C sky130_fd_sc_hd__nand3_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ hold153/X hold21/X _5692_/S VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4642_ _4698_/A _4656_/C _4647_/C _4657_/C VGND VGND VPWR VPWR _5173_/C sky130_fd_sc_hd__nor4b_2
XFILLER_163_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4573_ _4573_/A _4573_/B _4573_/C VGND VGND VPWR VPWR _4576_/C sky130_fd_sc_hd__nand3_1
Xmax_cap400 _5763_/X VGND VGND VPWR VPWR _6073_/B2 sky130_fd_sc_hd__buf_12
Xhold703 _5384_/X VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap411 hold38/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__buf_12
X_6312_ _7069_/Q _6103_/X _6119_/X _7053_/Q _6311_/X VGND VGND VPWR VPWR _6312_/X
+ sky130_fd_sc_hd__a221o_1
Xhold714 _7099_/Q VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlygate4sd3_1
X_3524_ _6524_/A _5476_/B _5273_/D VGND VGND VPWR VPWR _4121_/B sky130_fd_sc_hd__and3_4
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold725 hold725/A VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlygate4sd3_1
X_7292_ _7292_/A VGND VGND VPWR VPWR _7292_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold736 _5336_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap444 _4164_/Y VGND VGND VPWR VPWR _4166_/B sky130_fd_sc_hd__buf_2
Xhold747 _6550_/X VGND VGND VPWR VPWR _7276_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _6633_/Q VGND VGND VPWR VPWR hold758/X sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ _6242_/X _6243_/A1 _6443_/S VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__mux2_1
Xhold769 _7090_/Q VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ hold37/X hold42/X hold28/A _5324_/B VGND VGND VPWR VPWR _5684_/C sky130_fd_sc_hd__and4b_4
XFILLER_170_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6174_ _7120_/Q _5750_/X _6129_/D _6904_/Q _6173_/X VGND VGND VPWR VPWR _6181_/C
+ sky130_fd_sc_hd__a221o_1
X_3386_ _5324_/B hold37/X hold42/X _3987_/A VGND VGND VPWR VPWR _3386_/X sky130_fd_sc_hd__and4_2
XFILLER_85_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5125_ _5125_/A _5125_/B _5125_/C VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__and3_1
XFILLER_111_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1403 _6954_/Q VGND VGND VPWR VPWR hold666/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 _7088_/Q VGND VGND VPWR VPWR hold521/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__1184_ _3812_/X VGND VGND VPWR VPWR clkbuf_0__1184_/X sky130_fd_sc_hd__clkbuf_16
Xhold1425 _7135_/Q VGND VGND VPWR VPWR hold780/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 _3407_/X VGND VGND VPWR VPWR hold1436/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _7015_/Q VGND VGND VPWR VPWR hold1447/X sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _5060_/B _5143_/D _4815_/A _4475_/B _4476_/A VGND VGND VPWR VPWR _5056_/X
+ sky130_fd_sc_hd__a41o_1
Xhold1458 _7223_/Q VGND VGND VPWR VPWR _6475_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _7224_/Q VGND VGND VPWR VPWR _6476_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4007_ hold544/X _3916_/C _4010_/S VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__mux2_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5958_ _5795_/D _6072_/C _6894_/Q _5776_/X _6958_/Q VGND VGND VPWR VPWR _5958_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4909_ _4909_/A _4909_/B _4909_/C VGND VGND VPWR VPWR _4909_/X sky130_fd_sc_hd__and3_1
X_5889_ _6915_/Q _6028_/B _5934_/C VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__and3_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7256_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_188_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_5 _7236_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6930_ _7145_/CLK _6930_/D fanout600/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6861_ _7017_/CLK _6861_/D fanout606/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7264_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5812_ _5810_/X _6072_/B _5804_/X _5811_/X _5807_/X VGND VGND VPWR VPWR _5812_/X
+ sky130_fd_sc_hd__a2111o_1
X_6792_ _7156_/CLK _6792_/D fanout602/X VGND VGND VPWR VPWR _7291_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5743_ _5742_/X _5759_/B _5741_/Y _6143_/D _5712_/Y VGND VGND VPWR VPWR _7188_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5674_ _5692_/A1 _5674_/A1 _5674_/S VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4625_ _4670_/D _4625_/B _4859_/A VGND VGND VPWR VPWR _4675_/B sky130_fd_sc_hd__and3_1
XFILLER_175_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold500 _6915_/Q VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 _4074_/X VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _4556_/A _4556_/B _4556_/C VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__nor3_1
Xhold522 _7089_/Q VGND VGND VPWR VPWR hold522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _3990_/X VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3507_/A _3507_/B _3507_/C _3507_/D VGND VGND VPWR VPWR _3508_/D sky130_fd_sc_hd__nor4_1
Xhold544 _6664_/Q VGND VGND VPWR VPWR hold544/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold555 _6761_/Q VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7275_ _7275_/CLK _7275_/D fanout596/X VGND VGND VPWR VPWR _7275_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold566 _4065_/X VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4487_/A _4487_/B _4487_/C VGND VGND VPWR VPWR _4493_/C sky130_fd_sc_hd__nand3_1
Xhold577 hold577/A VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold588 _4015_/X VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6226_ _7042_/Q _6117_/C _6108_/X _6107_/X _7002_/Q VGND VGND VPWR VPWR _6226_/X
+ sky130_fd_sc_hd__a32o_1
X_3438_ _6530_/D _5548_/D _5494_/C VGND VGND VPWR VPWR _3438_/X sky130_fd_sc_hd__and3_4
Xhold599 _6707_/Q VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6935_/Q _6462_/B1 _6153_/X _6154_/X _6156_/X VGND VGND VPWR VPWR _6157_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _5620_/A _6548_/C VGND VGND VPWR VPWR _3369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1200 _4180_/X VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 _4083_/X VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1222 _7291_/A VGND VGND VPWR VPWR _4191_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5108_ _4716_/A _4738_/B _4689_/A VGND VGND VPWR VPWR _5109_/C sky130_fd_sc_hd__o21ai_1
Xhold1233 _4091_/X VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1244 hold1407/X VGND VGND VPWR VPWR _5558_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _6080_/X _6025_/B _6085_/X _6083_/X _6087_/X VGND VGND VPWR VPWR _6088_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold1255 _3946_/A1 VGND VGND VPWR VPWR hold581/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1266 _6476_/A1 VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1277 _3950_/A1 VGND VGND VPWR VPWR hold700/A sky130_fd_sc_hd__dlygate4sd3_1
X_5039_ _4815_/A _4333_/A _4843_/C _4843_/A VGND VGND VPWR VPWR _5234_/A sky130_fd_sc_hd__a211oi_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1288 _7169_/Q VGND VGND VPWR VPWR _5687_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_406 _6953_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1299 _7075_/Q VGND VGND VPWR VPWR _5580_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_417 _3922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_428 _6446_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _3312_/C sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _3313_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6498_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6503_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_6
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4410_ _4247_/Y _4248_/X _5128_/B _4256_/Y VGND VGND VPWR VPWR _4439_/D sky130_fd_sc_hd__o211a_1
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5390_ _3281_/Y _5394_/S _3922_/X _3559_/X VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_160_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4341_ _4815_/A _5089_/A VGND VGND VPWR VPWR _4487_/C sky130_fd_sc_hd__nand2_1
XFILLER_172_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7060_ _7174_/CLK _7060_/D fanout602/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_4
X_4272_ _4698_/A _4657_/C VGND VGND VPWR VPWR _4730_/A sky130_fd_sc_hd__nor2_8
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6011_ _6644_/Q _5783_/X _5791_/X _6560_/Q _6010_/X VGND VGND VPWR VPWR _6011_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6913_ _7067_/CLK _6913_/D fanout584/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6844_ _6855_/CLK hold48/X fanout583/X VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6775_ _6828_/CLK _6775_/D fanout573/X VGND VGND VPWR VPWR _6775_/Q sky130_fd_sc_hd__dfstp_2
X_3987_ _3987_/A _6548_/A _6548_/B _5657_/D VGND VGND VPWR VPWR _3992_/S sky130_fd_sc_hd__nand4_4
XFILLER_148_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5726_ _5782_/C _5795_/C _5795_/D VGND VGND VPWR VPWR _5726_/Y sky130_fd_sc_hd__nand3_4
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5657_ _6548_/B _5684_/B _5675_/D _5657_/D VGND VGND VPWR VPWR _5665_/S sky130_fd_sc_hd__nand4_4
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4608_ _5089_/A _4923_/B VGND VGND VPWR VPWR _4611_/B sky130_fd_sc_hd__nand2_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ hold24/X _5588_/A1 hold44/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__mux2_1
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold330 _7050_/Q VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold341 _5570_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _5040_/C _4529_/X _4535_/Y _4555_/B _4299_/Y VGND VGND VPWR VPWR _4556_/A
+ sky130_fd_sc_hd__o32ai_1
Xhold352 _6899_/Q VGND VGND VPWR VPWR hold352/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold363 _7170_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _5534_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _6744_/Q VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _7243_/Q VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__dlygate4sd3_1
X_7258_ _7259_/CLK _7258_/D _6472_/A VGND VGND VPWR VPWR _7258_/Q sky130_fd_sc_hd__dfrtp_4
X_6209_ _7129_/Q _6116_/X _6118_/X _7057_/Q _6208_/X VGND VGND VPWR VPWR _6214_/B
+ sky130_fd_sc_hd__a221o_1
X_7189_ _7254_/CLK _7189_/D fanout594/X VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_58_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1030 _3930_/X VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 _7248_/Q VGND VGND VPWR VPWR _6529_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 _7143_/Q VGND VGND VPWR VPWR _5658_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1063 _6958_/Q VGND VGND VPWR VPWR _5448_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 _4034_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 _7144_/Q VGND VGND VPWR VPWR _5659_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 _4095_/X VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_203 _6465_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _5476_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_225 _3922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _3340_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 hold83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 hold76/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _5323_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6967_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3910_ _6539_/A0 hold422/X _3912_/S VGND VGND VPWR VPWR _3910_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _4890_/A _5225_/A VGND VGND VPWR VPWR _4890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7248_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3841_ _7060_/Q _3563_/A _3902_/A3 _3488_/X _7076_/Q VGND VGND VPWR VPWR _3841_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6560_ _6689_/CLK _6560_/D fanout580/X VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfrtp_4
X_3772_ _6737_/Q _3386_/X wire447/X _3563_/X _7027_/Q VGND VGND VPWR VPWR _3772_/X
+ sky130_fd_sc_hd__a32o_1
X_5511_ _6511_/A1 hold426/X _5511_/S VGND VGND VPWR VPWR _5511_/X sky130_fd_sc_hd__mux2_1
X_6491_ _7259_/Q _6491_/A2 _6491_/B1 _7258_/Q VGND VGND VPWR VPWR _6491_/X sky130_fd_sc_hd__a22o_1
X_5442_ hold401/X _3916_/C _5448_/S VGND VGND VPWR VPWR _5442_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5373_ hold482/X _3925_/C _5376_/S VGND VGND VPWR VPWR _5373_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7097_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7112_ _7167_/CLK _7112_/D fanout604/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfstp_1
X_4324_ _4691_/B _4254_/Y _4304_/Y _4870_/B _4320_/Y VGND VGND VPWR VPWR _4509_/A
+ sky130_fd_sc_hd__o32a_2
XFILLER_59_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7043_ _7131_/CLK _7043_/D fanout606/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_4
X_4255_ _4255_/A _4970_/D _4722_/A _4777_/A VGND VGND VPWR VPWR _4429_/D sky130_fd_sc_hd__nand4_4
XFILLER_101_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4186_ _4186_/A0 _4185_/X _4188_/S VGND VGND VPWR VPWR _4186_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7171_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_3_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_82_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6827_ _6827_/CLK _6827_/D fanout573/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6758_ _6781_/CLK _6758_/D _3291_/A VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ _7177_/Q _7178_/Q _5710_/D _7179_/Q VGND VGND VPWR VPWR _5711_/B sky130_fd_sc_hd__a31o_1
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6689_ _6689_/CLK _6689_/D fanout578/X VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold160 hold160/A VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _5374_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _7133_/Q VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold193 _5663_/X VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4040_ _3925_/C hold430/X _4040_/S VGND VGND VPWR VPWR _4040_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5991_ _7244_/Q _5782_/C _6010_/D _6009_/C _6648_/Q VGND VGND VPWR VPWR _5991_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_91_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4942_ _4799_/A _4748_/B _4747_/Y _4719_/B _4945_/B VGND VGND VPWR VPWR _4942_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4873_ _4718_/D _4687_/B _5255_/C _4377_/X VGND VGND VPWR VPWR _4876_/B sky130_fd_sc_hd__a22oi_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6612_ _7256_/CLK _6612_/D VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3824_ _7164_/Q _3509_/X _3821_/X _3823_/X VGND VGND VPWR VPWR _3825_/D sky130_fd_sc_hd__a211o_1
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3755_ input7/X _4127_/C _5476_/C _5311_/C VGND VGND VPWR VPWR _3755_/X sky130_fd_sc_hd__and4_1
X_6543_ _6543_/A0 hold866/X _6547_/S VGND VGND VPWR VPWR _6543_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3686_ _6690_/Q _3481_/X _3682_/X _3683_/X _3685_/X VGND VGND VPWR VPWR _3686_/X
+ sky130_fd_sc_hd__a2111o_1
X_6474_ _3632_/Y _6474_/A1 _6480_/S VGND VGND VPWR VPWR _7222_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5425_ _3919_/C hold288/X _5430_/S VGND VGND VPWR VPWR _5425_/X sky130_fd_sc_hd__mux2_1
Xoutput210 _3278_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
Xoutput221 _7294_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput232 _7304_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput243 _7284_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput254 _7312_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_5356_ _6505_/A1 hold282/X _5358_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
Xoutput265 _6821_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
Xoutput276 _6731_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput287 _6741_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
Xoutput298 _6839_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
X_4307_ _4307_/A _4307_/B _4310_/D _4760_/B VGND VGND VPWR VPWR _4544_/D sky130_fd_sc_hd__nand4_4
X_5287_ hold969/X _6535_/A0 _5287_/S VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4238_ _5042_/A VGND VGND VPWR VPWR _4488_/B sky130_fd_sc_hd__inv_2
X_7026_ _7162_/CLK _7026_/D fanout605/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ _7249_/Q _5324_/B VGND VGND VPWR VPWR _4170_/D sky130_fd_sc_hd__nand2b_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire348 _3776_/Y VGND VGND VPWR VPWR _3811_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire359 _5124_/Y VGND VGND VPWR VPWR _5125_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_139_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout470 hold55/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__buf_8
Xfanout481 _3370_/B VGND VGND VPWR VPWR _4152_/B sky130_fd_sc_hd__buf_4
XFILLER_93_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout492 hold17/X VGND VGND VPWR VPWR _5630_/A sky130_fd_sc_hd__buf_8
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ hold56/A _3540_/B VGND VGND VPWR VPWR _3540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold907 _6654_/Q VGND VGND VPWR VPWR hold907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 _5405_/X VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3471_ _4127_/C _5575_/D _3528_/C VGND VGND VPWR VPWR _3471_/X sky130_fd_sc_hd__and3_2
Xhold929 _6673_/Q VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5210_ _5210_/A _5249_/B _5210_/C VGND VGND VPWR VPWR _5210_/X sky130_fd_sc_hd__and3_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6190_ _6190_/A _6190_/B _6190_/C _6440_/D VGND VGND VPWR VPWR _6190_/Y sky130_fd_sc_hd__nor4_1
X_5141_ _4428_/Y _4661_/X _5140_/X _5044_/A VGND VGND VPWR VPWR _5141_/X sky130_fd_sc_hd__o31a_1
XFILLER_97_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5072_ _4946_/X _4633_/Y _4613_/Y _4635_/Y _5248_/A3 VGND VGND VPWR VPWR _5270_/C
+ sky130_fd_sc_hd__a311o_1
X_4023_ _6524_/A _6536_/B _6536_/D _4158_/D VGND VGND VPWR VPWR _4028_/S sky130_fd_sc_hd__and4_2
XFILLER_37_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5974_ _5964_/X _5967_/X _5974_/C _5974_/D VGND VGND VPWR VPWR _5974_/Y sky130_fd_sc_hd__nand4bb_2
XFILLER_80_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4925_ _4897_/X _4923_/X _4925_/C _4925_/D VGND VGND VPWR VPWR _4928_/A sky130_fd_sc_hd__and4bb_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4856_ _4878_/A _4987_/A _4987_/B VGND VGND VPWR VPWR _4856_/X sky130_fd_sc_hd__and3_1
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3807_ _6662_/Q _3447_/X _5404_/B _6923_/Q _3806_/X VGND VGND VPWR VPWR _3807_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4787_ _4788_/A _4777_/C _4786_/X _4785_/Y VGND VGND VPWR VPWR _4790_/C sky130_fd_sc_hd__a211oi_1
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ _6550_/A0 hold662/X _6529_/S VGND VGND VPWR VPWR _6526_/X sky130_fd_sc_hd__mux2_1
X_3738_ _7162_/Q _3509_/X _3521_/X _7170_/Q VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6457_ _6624_/Q _6136_/A wire392/X _6454_/X _6456_/X VGND VGND VPWR VPWR _6457_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_173_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3669_ _6770_/Q _3482_/X _3665_/X _3667_/X _3668_/X VGND VGND VPWR VPWR _3669_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5408_ _3922_/C hold110/X _5412_/S VGND VGND VPWR VPWR _5408_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6388_ _7240_/Q _6115_/X _6385_/X _6387_/X VGND VGND VPWR VPWR _6389_/C sky130_fd_sc_hd__a211o_1
XFILLER_88_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5339_ hold5/X hold228/X _5340_/S VGND VGND VPWR VPWR _5339_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7065_/CLK _7009_/D fanout590/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7218_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3799_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4719_/B _4792_/C VGND VGND VPWR VPWR _4711_/C sky130_fd_sc_hd__nand2_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ hold864/X _6505_/A1 _5692_/S VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__mux2_1
X_4641_ _4718_/D _4641_/B VGND VGND VPWR VPWR _4685_/D sky130_fd_sc_hd__nand2_1
XFILLER_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4572_ _4751_/A _4923_/A _4606_/D _4589_/C VGND VGND VPWR VPWR _4573_/C sky130_fd_sc_hd__nand4_1
XFILLER_190_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap401 _6446_/B VGND VGND VPWR VPWR _6176_/B sky130_fd_sc_hd__buf_12
XFILLER_116_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6311_ _7005_/Q _6465_/A2 wire392/X _6325_/A2 _6885_/Q VGND VGND VPWR VPWR _6311_/X
+ sky130_fd_sc_hd__a32o_1
Xhold704 _7157_/Q VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3523_ _3523_/A _3523_/B _3523_/C _3523_/D VGND VGND VPWR VPWR _3523_/Y sky130_fd_sc_hd__nor4_1
XFILLER_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold715 _5607_/X VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 hold726/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
X_7291_ _7291_/A VGND VGND VPWR VPWR _7291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold737 _6875_/Q VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold748 _7146_/Q VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 _3970_/X VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3454_ _6959_/Q _3452_/X _4187_/S input71/X _3451_/X VGND VGND VPWR VPWR _3462_/C
+ sky130_fd_sc_hd__a221o_1
X_6242_ _6292_/S _6242_/A2 _6240_/Y _6241_/X VGND VGND VPWR VPWR _6242_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6173_ _6944_/Q _6347_/C _6425_/C _6116_/X _7128_/Q VGND VGND VPWR VPWR _6173_/X
+ sky130_fd_sc_hd__a32o_1
X_3385_ _5324_/B hold37/X hold42/X VGND VGND VPWR VPWR _3385_/X sky130_fd_sc_hd__and3_1
X_5124_ _4721_/C _4675_/B _5007_/C _4626_/X _5007_/A VGND VGND VPWR VPWR _5124_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1404 _5444_/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 _6692_/Q VGND VGND VPWR VPWR hold430/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1426 _7000_/Q VGND VGND VPWR VPWR hold458/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _5468_/X VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _5143_/A _5143_/C _5260_/B _5055_/D VGND VGND VPWR VPWR _5055_/Y sky130_fd_sc_hd__nand4_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1448 _6586_/Q VGND VGND VPWR VPWR _3906_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _7228_/Q VGND VGND VPWR VPWR _6480_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4006_ _4006_/A0 _4152_/B _4010_/S VGND VGND VPWR VPWR _4006_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _7094_/Q _5826_/B wire398/X _5795_/X _6902_/Q VGND VGND VPWR VPWR _5957_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_71_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4908_ _4522_/Y _4550_/Y _4648_/Y _4555_/B _5040_/C VGND VGND VPWR VPWR _4909_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5888_ hold91/A _5934_/C _5782_/C _5795_/C VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__o211a_1
XFILLER_166_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4839_ _5040_/A _4466_/X _4811_/X _4836_/X VGND VGND VPWR VPWR _4841_/A sky130_fd_sc_hd__o211a_1
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _7259_/Q _6509_/A2 _6509_/B1 _7258_/Q VGND VGND VPWR VPWR _6509_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold20 hold31/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__buf_8
XFILLER_152_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 _5959_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6860_ _7114_/CLK _6860_/D fanout604/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_2
X_5811_ _7103_/Q _6086_/B1 _5767_/X _7111_/Q _5792_/X VGND VGND VPWR VPWR _5811_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6791_ _6967_/CLK _6791_/D fanout585/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5742_ _7186_/Q _7185_/Q _6141_/B _6143_/D VGND VGND VPWR VPWR _5742_/X sky130_fd_sc_hd__a31o_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5673_ _5674_/S hold704/X _3550_/X _4073_/X VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4624_ _4984_/A _5128_/A _4704_/B VGND VGND VPWR VPWR _4723_/A sky130_fd_sc_hd__and3_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold501 _5400_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4555_ _5040_/C _4555_/B VGND VGND VPWR VPWR _4556_/B sky130_fd_sc_hd__nor2_1
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _5596_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold534/A VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _6653_/Q _3502_/X _3503_/X _7135_/Q _3505_/X VGND VGND VPWR VPWR _3507_/D
+ sky130_fd_sc_hd__a221o_1
Xhold545 _4007_/X VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _4137_/X VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7274_ _7274_/CLK _7274_/D fanout577/X VGND VGND VPWR VPWR _7274_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4486_ _4689_/B _4485_/X _4482_/Y VGND VGND VPWR VPWR _4487_/A sky130_fd_sc_hd__o21ai_1
XFILLER_89_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold567 _6930_/Q VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 hold578/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
Xhold589 hold589/A VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6954_/Q _6142_/X _6144_/X _7082_/Q _6224_/X VGND VGND VPWR VPWR _6230_/B
+ sky130_fd_sc_hd__a221o_1
X_3437_ _3437_/A _3437_/B _3437_/C _3437_/D VGND VGND VPWR VPWR _3508_/A sky130_fd_sc_hd__nor4_1
XFILLER_131_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _7103_/Q _6112_/X _6119_/X _7047_/Q _6155_/X VGND VGND VPWR VPWR _6156_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3368_ hold65/X hold26/X hold71/X _5620_/A VGND VGND VPWR VPWR _3368_/X sky130_fd_sc_hd__and4_4
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1201 _7295_/A VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 _7284_/A VGND VGND VPWR VPWR _4087_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1223 _4191_/X VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5107_ _5103_/X _5105_/X _5180_/A VGND VGND VPWR VPWR _5107_/X sky130_fd_sc_hd__o21ba_1
Xhold1234 hold1362/X VGND VGND VPWR VPWR _5369_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6087_ _6647_/Q _5783_/X _5784_/X _6624_/Q _6086_/X VGND VGND VPWR VPWR _6087_/X
+ sky130_fd_sc_hd__a221o_1
X_3299_ _7177_/Q _7176_/Q _7178_/Q _7179_/Q VGND VGND VPWR VPWR _3300_/B sky130_fd_sc_hd__nand4bb_2
Xhold1245 hold1412/X VGND VGND VPWR VPWR _5441_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _3906_/A1 VGND VGND VPWR VPWR hold579/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _3962_/A1 VGND VGND VPWR VPWR hold633/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _6477_/A1 VGND VGND VPWR VPWR hold754/A sky130_fd_sc_hd__dlygate4sd3_1
X_5038_ _4976_/C _5035_/X _5037_/X _4516_/A VGND VGND VPWR VPWR _5038_/X sky130_fd_sc_hd__o31a_1
Xhold1289 _6969_/Q VGND VGND VPWR VPWR _5461_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_407 _6609_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_418 _3922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_429 _5795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6989_ _7143_/CLK _6989_/D fanout588/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR input110/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4557_/A sky130_fd_sc_hd__buf_4
XFILLER_88_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6489_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6492_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6495_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6481_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4340_ _4620_/A _4606_/B _4597_/B VGND VGND VPWR VPWR _5089_/A sky130_fd_sc_hd__and3_2
XFILLER_99_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4271_ _4970_/D _4940_/C VGND VGND VPWR VPWR _4271_/Y sky130_fd_sc_hd__nand2_4
XFILLER_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6010_ _7245_/Q _6059_/S _6010_/C _6010_/D VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__and4_1
XFILLER_140_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ _7087_/CLK _6912_/D fanout589/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6843_ _6843_/CLK _6843_/D fanout584/X VGND VGND VPWR VPWR _7281_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6774_ _6835_/CLK _6774_/D fanout583/X VGND VGND VPWR VPWR _6774_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3986_ _3986_/A0 _6535_/A0 _3986_/S VGND VGND VPWR VPWR _3986_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5725_ _7183_/Q _5712_/Y _5724_/X _5759_/B VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__a22o_1
XFILLER_176_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5656_ _4053_/B hold216/X _5656_/S VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4607_ _4607_/A _4607_/B _4607_/C _4607_/D VGND VGND VPWR VPWR _4611_/A sky130_fd_sc_hd__nor4_1
XFILLER_191_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5587_ _3918_/B hold651/X hold44/X VGND VGND VPWR VPWR _5587_/X sky130_fd_sc_hd__mux2_1
Xhold320 _6698_/Q VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold331 _5552_/X VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4538_ _5090_/A _5090_/B _4597_/B _4561_/B VGND VGND VPWR VPWR _4555_/B sky130_fd_sc_hd__nand4_2
XFILLER_117_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold342 hold342/A VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _5382_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold364 _5688_/X VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold375/A VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7257_ _7259_/CLK _7257_/D _6472_/A VGND VGND VPWR VPWR _7257_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold386 _4117_/X VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _4469_/A _4469_/B _4469_/C VGND VGND VPWR VPWR _4476_/C sky130_fd_sc_hd__nand3_1
Xhold397 _6523_/X VGND VGND VPWR VPWR _7243_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _7169_/Q _6130_/A _6114_/X _6130_/X _6929_/Q VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a32o_1
X_7188_ _7259_/CLK _7188_/D fanout594/X VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _7186_/Q _6141_/B _6143_/D _7185_/Q VGND VGND VPWR VPWR _6139_/X sky130_fd_sc_hd__and4bb_4
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _4153_/X VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1031 _7264_/Q VGND VGND VPWR VPWR _6535_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1042 _6529_/X VGND VGND VPWR VPWR _7248_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1053 _6910_/Q VGND VGND VPWR VPWR _5394_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1064 _5448_/X VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1075 _7042_/Q VGND VGND VPWR VPWR _5543_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 _5659_/X VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _6602_/Q VGND VGND VPWR VPWR _3934_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 _6465_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _5795_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _3919_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 hold2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_248 hold89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 _3542_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6676_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3840_ _6828_/Q _3497_/X _3528_/X input17/X _3839_/X VGND VGND VPWR VPWR _3843_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3771_ _7043_/Q _5512_/B _5684_/C _3565_/X _6652_/Q VGND VGND VPWR VPWR _3771_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ hold21/X hold176/X _5511_/S VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6490_ _6489_/X hold211/A _6511_/S VGND VGND VPWR VPWR _7229_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5441_ _5441_/A0 _5649_/A0 _5448_/S VGND VGND VPWR VPWR _5441_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5372_ _3282_/Y _5376_/S _3922_/X _5372_/B2 VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__a2bb2o_1
X_7111_ _7111_/CLK _7111_/D fanout599/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_141_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4323_ _4320_/A _4523_/C _4322_/Y VGND VGND VPWR VPWR _4509_/D sky130_fd_sc_hd__o21ai_2
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7042_ _7130_/CLK _7042_/D fanout600/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_4
X_4254_ _4657_/C _4698_/A VGND VGND VPWR VPWR _4254_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_101_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4185_ hold136/X _4051_/X _4187_/S VGND VGND VPWR VPWR _4185_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6826_ _6827_/CLK _6826_/D fanout573/X VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6757_ _7239_/CLK _6757_/D fanout581/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_1
X_3969_ _5494_/A hold64/X _3969_/C VGND VGND VPWR VPWR _3974_/S sky130_fd_sc_hd__and3_4
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5708_ _5711_/A _5708_/B _5708_/C VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__and3_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6688_ _7268_/CLK _6688_/D fanout572/X VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5639_ hold8/X _5639_/B VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__nand2_8
XFILLER_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold150 _5437_/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7309_ _7309_/A VGND VGND VPWR VPWR _7309_/X sky130_fd_sc_hd__clkbuf_1
Xhold161 _6982_/Q VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _7062_/Q VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold183 _5646_/X VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _6902_/Q VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5990_ _6678_/Q _6072_/C _6028_/C VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__and3_1
X_4941_ _4635_/Y _4745_/Y _4939_/Y _4629_/Y VGND VGND VPWR VPWR _5270_/D sky130_fd_sc_hd__o22a_1
X_4872_ _4872_/A _4872_/B _4872_/C _4872_/D VGND VGND VPWR VPWR _4876_/A sky130_fd_sc_hd__nor4_1
X_6611_ _6689_/CLK _6611_/D fanout580/X VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3823_ _6900_/Q _5377_/C _3521_/X _7172_/Q _3822_/X VGND VGND VPWR VPWR _3823_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6542_ _6542_/A _6542_/B VGND VGND VPWR VPWR _6547_/S sky130_fd_sc_hd__nand2_4
XFILLER_158_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3754_ _3753_/X _3754_/A1 _3906_/S VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6473_ _3568_/Y _6473_/A1 _6480_/S VGND VGND VPWR VPWR _7221_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3685_ _6881_/Q _5359_/B _3547_/X _7033_/Q _3684_/X VGND VGND VPWR VPWR _3685_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_106_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5424_ _3916_/C hold348/X _5430_/S VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput200 _3253_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
XFILLER_160_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput211 _3277_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _3335_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput233 _7282_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput244 _7285_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
X_5355_ _3924_/B hold737/X _5358_/S VGND VGND VPWR VPWR _5355_/X sky130_fd_sc_hd__mux2_1
Xoutput255 _3293_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
Xoutput266 _6822_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput277 _6732_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
XFILLER_87_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput288 _6742_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
X_4306_ _4284_/C _4310_/B _4282_/C _4308_/D _4760_/B VGND VGND VPWR VPWR _4312_/A
+ sky130_fd_sc_hd__a41o_1
Xoutput299 _6840_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
X_5286_ hold437/X _6546_/A0 _5287_/S VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7025_ _7099_/CLK _7025_/D fanout598/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4237_ _4243_/A _4243_/B VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__nand2_4
XFILLER_114_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4168_ _7257_/D _4168_/B _7258_/D _4167_/Y VGND VGND VPWR VPWR _4170_/C sky130_fd_sc_hd__nor4b_2
XFILLER_110_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7237_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4099_ _5494_/A _3571_/X _3924_/X _4102_/S _4099_/B2 VGND VGND VPWR VPWR _4099_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6809_ _7254_/CLK _6809_/D _6472_/A VGND VGND VPWR VPWR _6809_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire349 _3717_/Y VGND VGND VPWR VPWR _3752_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_139_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7151_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_85_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6812_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout460 _5331_/C VGND VGND VPWR VPWR _5327_/D sky130_fd_sc_hd__buf_12
XFILLER_120_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout471 _5449_/B VGND VGND VPWR VPWR _4127_/C sky130_fd_sc_hd__buf_12
Xfanout482 _6543_/A0 VGND VGND VPWR VPWR _3370_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout493 _5620_/A VGND VGND VPWR VPWR _5476_/B sky130_fd_sc_hd__buf_12
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk _7277_/CLK VGND VGND VPWR VPWR _7111_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7132_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold908 _3995_/X VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold919 _7161_/Q VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3470_ _6524_/A _6530_/C _6530_/D VGND VGND VPWR VPWR _3470_/X sky130_fd_sc_hd__and3_2
XFILLER_127_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5140_ _5260_/A _5140_/B _5140_/C VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__and3_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5071_ _4946_/X _4633_/Y _4613_/Y _5248_/A3 _4643_/Y VGND VGND VPWR VPWR _5073_/B
+ sky130_fd_sc_hd__a311o_1
X_4022_ _4017_/B _3925_/X _4021_/S hold976/X VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5973_ _7110_/Q _5764_/X _5784_/X _7030_/Q _5972_/X VGND VGND VPWR VPWR _5974_/D
+ sky130_fd_sc_hd__a221oi_2
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4924_ _4211_/X _4581_/B _4589_/C _4923_/X VGND VGND VPWR VPWR _5177_/A sky130_fd_sc_hd__a31o_1
XFILLER_178_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4855_ _5255_/A _4718_/D _4755_/B _4982_/D _4377_/X VGND VGND VPWR VPWR _4983_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3806_ _6915_/Q _4158_/D _5281_/A2 _3492_/X _6667_/Q VGND VGND VPWR VPWR _3806_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_178_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4786_ _4788_/A _4786_/B _4939_/B VGND VGND VPWR VPWR _4786_/X sky130_fd_sc_hd__and3_1
X_6525_ _6543_/A0 hold872/X _6529_/S VGND VGND VPWR VPWR _6525_/X sky130_fd_sc_hd__mux2_1
X_3737_ _7098_/Q _3510_/X _3729_/X _3731_/X _3736_/X VGND VGND VPWR VPWR _3752_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_146_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6456_ _6578_/Q _6104_/X _6129_/D _6672_/Q _6455_/X VGND VGND VPWR VPWR _6456_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3668_ _6929_/Q _3533_/C _3902_/A3 _3434_/X _6820_/Q VGND VGND VPWR VPWR _3668_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5407_ _5404_/B _3919_/X _5412_/S hold948/X VGND VGND VPWR VPWR _5407_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6387_ _7266_/Q _6106_/X _6462_/B1 _6654_/Q _6386_/X VGND VGND VPWR VPWR _6387_/X
+ sky130_fd_sc_hd__a221o_1
X_3599_ _7266_/Q _6536_/A _4139_/C _3927_/B _6598_/Q VGND VGND VPWR VPWR _3599_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5338_ _5334_/B _3922_/X _5340_/S hold844/X VGND VGND VPWR VPWR _5338_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5269_ _4718_/D _4786_/B _5263_/C _4939_/B VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__o211a_1
X_7008_ _7123_/CLK _7008_/D fanout606/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_141_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4640_ _4640_/A _4939_/B VGND VGND VPWR VPWR _4640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4571_ _4597_/C _4923_/A _4606_/D _4589_/C VGND VGND VPWR VPWR _4573_/B sky130_fd_sc_hd__nand4_1
X_6310_ _6989_/Q _6098_/X _6129_/B _6925_/Q VGND VGND VPWR VPWR _6310_/X sky130_fd_sc_hd__a22o_1
X_3522_ _6559_/Q _6536_/A _5311_/B _3521_/X _7167_/Q VGND VGND VPWR VPWR _3523_/D
+ sky130_fd_sc_hd__a32o_1
Xhold705 _5673_/X VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7290_ _7290_/A VGND VGND VPWR VPWR _7290_/X sky130_fd_sc_hd__clkbuf_2
Xhold716 _7037_/Q VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold727 _7093_/Q VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap435 _4484_/C VGND VGND VPWR VPWR _5060_/C sky130_fd_sc_hd__buf_4
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap446 wire447/X VGND VGND VPWR VPWR _3721_/A3 sky130_fd_sc_hd__clkbuf_2
Xhold738 _5355_/X VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6241_ _6874_/Q _6466_/A1 _5759_/A VGND VGND VPWR VPWR _6241_/X sky130_fd_sc_hd__o21a_1
Xhold749 _5661_/X VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3453_ _6530_/D _5666_/C _5575_/D VGND VGND VPWR VPWR _4187_/S sky130_fd_sc_hd__and3_4
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6172_ _7144_/Q _6113_/X _6115_/X _7136_/Q _6171_/X VGND VGND VPWR VPWR _6181_/B
+ sky130_fd_sc_hd__a221o_1
X_3384_ _6535_/A0 _3384_/A1 _3384_/S VGND VGND VPWR VPWR _3384_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5123_ _4650_/Y _4699_/Y _4881_/B _4999_/X _5122_/Y VGND VGND VPWR VPWR _5125_/B
+ sky130_fd_sc_hd__o2111a_1
Xhold1405 _6665_/Q VGND VGND VPWR VPWR hold975/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _4040_/X VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 _7016_/Q VGND VGND VPWR VPWR hold253/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1438 _6691_/Q VGND VGND VPWR VPWR hold554/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5054_ _5260_/B _5143_/C _4394_/X _5053_/X _5052_/X VGND VGND VPWR VPWR _5058_/A
+ sky130_fd_sc_hd__a311oi_1
XFILLER_38_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1449 _6735_/Q VGND VGND VPWR VPWR hold974/A sky130_fd_sc_hd__dlygate4sd3_1
X_4005_ _6536_/B _6548_/C _4127_/C _4158_/D VGND VGND VPWR VPWR _4010_/S sky130_fd_sc_hd__and4_2
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5956_ _7006_/Q _5795_/D _6010_/C _5815_/B VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__o211a_1
X_4907_ _4907_/A _4907_/B _5020_/D VGND VGND VPWR VPWR _4909_/B sky130_fd_sc_hd__nor3b_1
X_5887_ _7123_/Q _5965_/B _5911_/C VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__and3_1
XFILLER_21_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4838_ _4549_/D _4632_/B _4633_/B _4751_/A VGND VGND VPWR VPWR _4838_/X sky130_fd_sc_hd__a31o_1
XFILLER_193_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4769_ _5263_/C _4775_/B VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6508_ _6507_/X hold21/A _6511_/S VGND VGND VPWR VPWR _7235_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6439_ _6676_/Q _6129_/A _6436_/X _6438_/X VGND VGND VPWR VPWR _6440_/C sky130_fd_sc_hd__a211o_1
XFILLER_134_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__buf_12
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__buf_6
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_7 _6138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5810_ _7063_/Q _5723_/X _6003_/C _7031_/Q _5809_/X VGND VGND VPWR VPWR _5810_/X
+ sky130_fd_sc_hd__a221o_1
X_6790_ _7156_/CLK _6790_/D fanout602/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5741_ _7186_/Q _7185_/Q _6143_/D _6141_/B VGND VGND VPWR VPWR _5741_/Y sky130_fd_sc_hd__nand4_2
XFILLER_50_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5672_ _4049_/B hold314/X _5674_/S VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4623_ _4290_/Y _4409_/C _7258_/Q VGND VGND VPWR VPWR _4623_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4554_ _4554_/A _4554_/B _4554_/C _4554_/D VGND VGND VPWR VPWR _4556_/C sky130_fd_sc_hd__nand4_1
Xhold502 _6980_/Q VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _6666_/Q VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold524 _6557_/Q VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _6975_/Q _5494_/C _5281_/A2 _3504_/X input4/X VGND VGND VPWR VPWR _3505_/X
+ sky130_fd_sc_hd__a32o_1
X_7273_ _7273_/CLK _7273_/D fanout579/X VGND VGND VPWR VPWR _7273_/Q sky130_fd_sc_hd__dfrtp_2
Xhold535 hold535/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xhold546 _6751_/Q VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__dlygate4sd3_1
X_4485_ _4511_/A _4208_/Y _4244_/Y _4344_/Y _5146_/D VGND VGND VPWR VPWR _4485_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold557 hold557/A VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold568 _5417_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold579 hold579/A VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _7066_/Q _6138_/B _6102_/X _6129_/A _6898_/Q VGND VGND VPWR VPWR _6224_/X
+ sky130_fd_sc_hd__a32o_1
X_3436_ _6633_/Q _3969_/C _3432_/X _6602_/Q _3435_/X VGND VGND VPWR VPWR _3437_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7023_/Q _6136_/A wire392/X _6323_/B1 _6959_/Q VGND VGND VPWR VPWR _6155_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _5324_/B hold26/X hold71/X VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__and3_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _4199_/X VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5140_/C _5036_/A _4619_/X _4976_/D _4516_/Y VGND VGND VPWR VPWR _5180_/A
+ sky130_fd_sc_hd__a2111o_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _4087_/X VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _6658_/Q VGND VGND VPWR VPWR _4000_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6086_ _6815_/Q _6010_/C _5815_/B _6086_/B1 _7279_/Q VGND VGND VPWR VPWR _6086_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1235 hold1372/X VGND VGND VPWR VPWR _4104_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3298_ _6800_/Q _5694_/A _3297_/Y VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__a21bo_1
Xhold1246 hold1324/X VGND VGND VPWR VPWR _5396_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1257 _3964_/A1 VGND VGND VPWR VPWR hold577/A sky130_fd_sc_hd__dlygate4sd3_1
X_5037_ _4738_/B _4718_/D _4620_/B _4620_/A VGND VGND VPWR VPWR _5037_/X sky130_fd_sc_hd__o211a_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1268 _6474_/A1 VGND VGND VPWR VPWR hold649/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _7220_/Q VGND VGND VPWR VPWR hold1279/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_408 _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_419 _3918_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6988_ _7143_/CLK hold87/X fanout588/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5939_ _6885_/Q _5768_/X _5794_/X _6925_/Q _5938_/X VGND VGND VPWR VPWR _5939_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4229_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4747_/A sky130_fd_sc_hd__buf_8
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6495_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6501_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6506_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6482_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4270_ _4632_/A _4511_/A _4632_/C _4612_/C VGND VGND VPWR VPWR _4716_/A sky130_fd_sc_hd__and4bb_4
XFILLER_141_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6911_ _7087_/CLK _6911_/D fanout589/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_47_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6842_ _7265_/CLK _6842_/D fanout575/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6773_ _6827_/CLK _6773_/D fanout573/X VGND VGND VPWR VPWR _6773_/Q sky130_fd_sc_hd__dfrtp_4
X_3985_ hold667/X _6540_/A0 _3986_/S VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5724_ _5782_/C _5795_/C _5721_/X VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5655_ _5494_/A _3503_/X _4051_/X _5656_/S hold807/X VGND VGND VPWR VPWR _5655_/X
+ sky130_fd_sc_hd__a32o_1
X_4606_ _4620_/A _4606_/B _4786_/B _4606_/D VGND VGND VPWR VPWR _4607_/C sky130_fd_sc_hd__and4_1
XFILLER_129_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5586_ _3915_/B hold274/X hold44/X VGND VGND VPWR VPWR _5586_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold310 _6897_/Q VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold321 _4050_/X VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _4523_/C _4523_/A _4509_/C _4522_/Y VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__a211o_1
Xhold332 _6905_/Q VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold343 hold343/A VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _6690_/Q VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _6873_/Q VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlygate4sd3_1
X_7256_ _7256_/CLK _7256_/D _6472_/A VGND VGND VPWR VPWR _7256_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4468_ _5060_/B _5060_/C _5044_/A _4738_/B VGND VGND VPWR VPWR _4469_/C sky130_fd_sc_hd__nand4_1
Xhold376 _7002_/Q VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _6960_/Q VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold398 hold398/A VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6207_ _6969_/Q _6097_/X _6098_/X _6985_/Q _6206_/X VGND VGND VPWR VPWR _6214_/A
+ sky130_fd_sc_hd__a221o_2
X_3419_ _3563_/A _6530_/D _5476_/C VGND VGND VPWR VPWR _5566_/B sky130_fd_sc_hd__and3_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7187_ _7259_/CLK _7187_/D fanout594/X VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_4
X_4399_ _4859_/C _5260_/B _4399_/C VGND VGND VPWR VPWR _4451_/A sky130_fd_sc_hd__and3_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6138_/A _6138_/B _6425_/B VGND VGND VPWR VPWR _6138_/X sky130_fd_sc_hd__and3_4
Xhold1010 _6906_/Q VGND VGND VPWR VPWR _3281_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1021 _6685_/Q VGND VGND VPWR VPWR _4032_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _6535_/X VGND VGND VPWR VPWR _7264_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1043 hold1380/X VGND VGND VPWR VPWR _5276_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6069_ _6090_/A2 _5761_/X _6068_/X VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__o21a_1
XFILLER_100_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1054 _5394_/X VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 _7166_/Q VGND VGND VPWR VPWR _5683_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 _5543_/X VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _6731_/Q VGND VGND VPWR VPWR _4101_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 _3934_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_205 _5795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_216 _6511_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_227 _3919_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 hold2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 hold89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3770_ _7099_/Q _3510_/X _6542_/B _7274_/Q _3769_/X VGND VGND VPWR VPWR _3770_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5440_ _5494_/A _5494_/C _5440_/C VGND VGND VPWR VPWR _5448_/S sky130_fd_sc_hd__and3_4
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ hold322/X _3919_/C _5376_/S VGND VGND VPWR VPWR _5371_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7110_ _7163_/CLK _7110_/D fanout610/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_1
X_4322_ _4246_/Y _4301_/Y _4662_/B VGND VGND VPWR VPWR _4322_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7041_ _7167_/CLK _7041_/D fanout604/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_2
X_4253_ _4657_/C _4698_/A VGND VGND VPWR VPWR _4777_/A sky130_fd_sc_hd__and2b_4
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4184_ _4184_/A0 _4183_/X _4188_/S VGND VGND VPWR VPWR _4184_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7219_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6825_ _6827_/CLK _6825_/D fanout573/X VGND VGND VPWR VPWR _6825_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6756_ _7241_/CLK _6756_/D fanout575/X VGND VGND VPWR VPWR _6756_/Q sky130_fd_sc_hd__dfrtp_4
X_3968_ _3905_/Y _3968_/A1 _3968_/S VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5707_ _7177_/Q _7176_/Q _5706_/D _7178_/Q VGND VGND VPWR VPWR _5708_/C sky130_fd_sc_hd__a31o_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6687_ _6687_/CLK _6687_/D fanout580/X VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3899_ _6950_/Q _3544_/X _3571_/X _6732_/Q _3898_/X VGND VGND VPWR VPWR _3904_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_164_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5638_ _5692_/A1 hold903/X hold29/X VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5569_ hold2/X hold155/X _5574_/S VGND VGND VPWR VPWR _5569_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold140 _6847_/Q VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlygate4sd3_1
X_7308_ _7308_/A VGND VGND VPWR VPWR _7308_/X sky130_fd_sc_hd__buf_2
XFILLER_104_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold151 _7029_/Q VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _5475_/X VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold173 _5565_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _7021_/Q VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold195 _5385_/X VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7239_ _7239_/CLK _7239_/D fanout574/X VGND VGND VPWR VPWR _7239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout620 _4494_/C VGND VGND VPWR VPWR _4632_/C sky130_fd_sc_hd__buf_12
XFILLER_104_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4940_ _4940_/A _4970_/D _4940_/C _4940_/D VGND VGND VPWR VPWR _4940_/Y sky130_fd_sc_hd__nand4_1
XFILLER_45_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4871_ _4853_/C _4640_/A _4945_/C _5255_/C _4878_/A VGND VGND VPWR VPWR _4872_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6610_ _7273_/CLK _6610_/D fanout579/X VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_4
X_3822_ _7052_/Q _5548_/C _3540_/B _3515_/X _7028_/Q VGND VGND VPWR VPWR _3822_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6541_ _3925_/C hold392/X _6541_/S VGND VGND VPWR VPWR _6541_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6671_/Q _3513_/X _3696_/X _3699_/X _3752_/Y VGND VGND VPWR VPWR _3753_/X
+ sky130_fd_sc_hd__a2111o_4
X_6472_ _6472_/A _7250_/Q VGND VGND VPWR VPWR _6480_/S sky130_fd_sc_hd__nand2_4
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3684_ _7097_/Q _3510_/X _5557_/B _7057_/Q VGND VGND VPWR VPWR _3684_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5423_ _5649_/A0 _5423_/A1 _5430_/S VGND VGND VPWR VPWR _5423_/X sky130_fd_sc_hd__mux2_1
Xoutput201 _3252_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3276_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
XFILLER_173_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput223 _7295_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
XFILLER_160_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput234 _7305_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
X_5354_ hold24/X hold234/X _5358_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
Xoutput245 _3334_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput256 _7313_/X VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput267 _6816_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
X_4305_ _4307_/A _4307_/B _4310_/D VGND VGND VPWR VPWR _4313_/A sky130_fd_sc_hd__nand3_4
Xoutput278 _6829_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
X_5285_ hold971/X _6539_/A0 _5287_/S VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__mux2_1
Xoutput289 _6735_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7024_ _7097_/CLK _7024_/D fanout600/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfstp_1
X_4236_ _4747_/A _4284_/C _4310_/B _4236_/D VGND VGND VPWR VPWR _4243_/B sky130_fd_sc_hd__nand4_4
X_4167_ _7254_/Q _7250_/Q VGND VGND VPWR VPWR _4167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4098_ _6546_/A0 hold465/X _4102_/S VGND VGND VPWR VPWR _4098_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_4_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7263_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6808_ _7254_/CLK _6808_/D _6472_/A VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_4
X_6739_ _6843_/CLK _6739_/D fanout584/X VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_139_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout461 _3409_/X VGND VGND VPWR VPWR _5331_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout472 _5449_/B VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__buf_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout483 _5667_/A0 VGND VGND VPWR VPWR _5649_/A0 sky130_fd_sc_hd__buf_6
XFILLER_101_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout494 hold1388/X VGND VGND VPWR VPWR _5620_/A sky130_fd_sc_hd__buf_12
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold909 _7070_/Q VGND VGND VPWR VPWR hold909/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_182_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5070_ _4722_/A _4674_/D _4950_/X _5066_/X _5069_/X VGND VGND VPWR VPWR _5070_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4021_ _6540_/A0 hold775/X _4021_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5972_ _7118_/Q _5767_/X _5780_/X _7102_/Q _5971_/X VGND VGND VPWR VPWR _5972_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4923_ _4923_/A _4923_/B _4923_/C VGND VGND VPWR VPWR _4923_/X sky130_fd_sc_hd__and3_1
XFILLER_33_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4854_ _4859_/C _4987_/A _4987_/B _4903_/B _4718_/D VGND VGND VPWR VPWR _4854_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3805_ _7163_/Q _3509_/X _3801_/X _3802_/X _3804_/X VGND VGND VPWR VPWR _3805_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4785_ _4613_/Y _4709_/Y _4745_/Y _4707_/Y _4784_/X VGND VGND VPWR VPWR _4785_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6524_ _6524_/A _6524_/B _6530_/C _6530_/D VGND VGND VPWR VPWR _6529_/S sky130_fd_sc_hd__nand4_4
X_3736_ _6832_/Q wire447/X _3457_/X _3733_/X _3735_/X VGND VGND VPWR VPWR _3736_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3667_ _6825_/Q _6524_/A _5331_/C _6536_/D _3666_/X VGND VGND VPWR VPWR _3667_/X
+ sky130_fd_sc_hd__a41o_1
X_6455_ _6637_/Q _6113_/X _6116_/X _6573_/Q _6444_/X VGND VGND VPWR VPWR _6455_/X
+ sky130_fd_sc_hd__a221o_1
X_5406_ _3540_/B _5422_/D _3916_/X _5412_/S hold854/X VGND VGND VPWR VPWR _5406_/X
+ sky130_fd_sc_hd__a32o_1
X_6386_ _6588_/Q _6138_/A _6110_/C _6107_/X _6812_/Q VGND VGND VPWR VPWR _6386_/X
+ sky130_fd_sc_hd__a32o_1
X_3598_ _6976_/Q _5273_/D _5281_/A2 _3531_/X _6754_/Q VGND VGND VPWR VPWR _3598_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5337_ _3918_/B hold240/X _5340_/S VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5268_ _5226_/Y _5258_/X _5267_/Y VGND VGND VPWR VPWR _5268_/Y sky130_fd_sc_hd__o21ai_1
X_7007_ _7007_/CLK _7007_/D fanout590/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4219_ _4219_/A _4219_/B VGND VGND VPWR VPWR _4307_/A sky130_fd_sc_hd__nor2_2
X_5199_ _4675_/A _5128_/A _4732_/C _4737_/B _4894_/X VGND VGND VPWR VPWR _5200_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4570_ _4570_/A _4570_/B _4570_/C VGND VGND VPWR VPWR _4573_/A sky130_fd_sc_hd__nor3_1
X_3521_ _5620_/A _5684_/B hold28/A VGND VGND VPWR VPWR _3521_/X sky130_fd_sc_hd__and3_4
XFILLER_128_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap414 _6139_/X VGND VGND VPWR VPWR _6425_/C sky130_fd_sc_hd__buf_12
Xhold706 hold706/A VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold717 _5537_/X VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold728 _5600_/X VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ _6221_/X _6240_/B _6240_/C VGND VGND VPWR VPWR _6240_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_155_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3452_ _4127_/C _5494_/C _5575_/D VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__and3_4
Xhold739 _7165_/Q VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6171_ _7000_/Q _6465_/A2 wire392/X _6462_/B1 _6936_/Q VGND VGND VPWR VPWR _6171_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_131_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3383_ _6540_/A0 hold733/X _3384_/S VGND VGND VPWR VPWR _3383_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5122_ _4704_/B _4375_/X _4738_/B _4705_/B _4884_/B VGND VGND VPWR VPWR _5122_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_69_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1406 _4008_/X VGND VGND VPWR VPWR _6665_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1417 _7254_/Q VGND VGND VPWR VPWR _7259_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5053_ _4738_/B _4597_/C _4838_/X _5260_/B _4460_/B VGND VGND VPWR VPWR _5053_/X
+ sky130_fd_sc_hd__o311a_1
Xhold1428 _5514_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 _4039_/X VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4004_ _4003_/S hold792/X _3447_/X _3925_/X VGND VGND VPWR VPWR _4004_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5955_ _5955_/A1 _5761_/X _5954_/X _5953_/X VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__o22a_1
X_4906_ _4522_/Y _4601_/Y _4658_/Y _4535_/Y _4558_/Y VGND VGND VPWR VPWR _5020_/D
+ sky130_fd_sc_hd__o32a_1
X_5886_ _5886_/A1 _5761_/X _5885_/X VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_84_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7007_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4837_ _4815_/A _5260_/B _4394_/X _4399_/C _4449_/B VGND VGND VPWR VPWR _4837_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4768_ _4923_/B _4641_/B _4767_/Y VGND VGND VPWR VPWR _4768_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6507_ _7258_/Q _6507_/A2 _6507_/B1 _4164_/Y _6506_/X VGND VGND VPWR VPWR _6507_/X
+ sky130_fd_sc_hd__a221o_1
X_3719_ _7106_/Q _6536_/A _5684_/C _3470_/X _7247_/Q VGND VGND VPWR VPWR _3719_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4699_ _4777_/A _4699_/B VGND VGND VPWR VPWR _4699_/Y sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_99_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6761_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6438_ _6605_/Q _6105_/X _6110_/X _6557_/Q _6437_/X VGND VGND VPWR VPWR _6438_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6369_ _7261_/Q _6425_/B _6425_/C _6097_/X _6759_/Q VGND VGND VPWR VPWR _6369_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_136_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_csclk _7277_/CLK VGND VGND VPWR VPWR _7072_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold11/A VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__buf_6
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold97/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7120_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _6444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5740_ _6143_/D _7187_/Q _6136_/A VGND VGND VPWR VPWR _6446_/B sky130_fd_sc_hd__and3_4
XFILLER_188_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5674_/S hold832/X _3550_/X _3925_/X VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__a22o_1
X_4622_ _4721_/C _4683_/C _4668_/C _4878_/B VGND VGND VPWR VPWR _4859_/D sky130_fd_sc_hd__o211a_2
X_4553_ _5090_/A _5090_/B _4620_/B _4923_/B VGND VGND VPWR VPWR _4554_/D sky130_fd_sc_hd__nand4_1
XFILLER_190_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold503 _5473_/X VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold514 _4009_/X VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold525 _3365_/X VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _6536_/C _4127_/C _3528_/C VGND VGND VPWR VPWR _3504_/X sky130_fd_sc_hd__and3_2
X_7272_ _7274_/CLK _7272_/D fanout579/X VGND VGND VPWR VPWR _7272_/Q sky130_fd_sc_hd__dfstp_2
Xhold536 _7273_/Q VGND VGND VPWR VPWR hold536/X sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _5060_/B _4801_/B _4484_/C _4484_/D VGND VGND VPWR VPWR _5146_/D sky130_fd_sc_hd__nand4_2
Xhold547 _4125_/X VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 hold558/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
X_3435_ _6818_/Q _5327_/D _5440_/C _3433_/X _6935_/Q VGND VGND VPWR VPWR _3435_/X
+ sky130_fd_sc_hd__a32o_1
X_6223_ _6962_/Q _6323_/B1 _6136_/X _7026_/Q _6222_/X VGND VGND VPWR VPWR _6230_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold569 _6703_/Q VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _7039_/Q _6444_/C _6465_/A3 _6099_/X VGND VGND VPWR VPWR _6154_/X sky130_fd_sc_hd__a31o_1
X_3366_ _3925_/C hold454/X _3366_/S VGND VGND VPWR VPWR _3366_/X sky130_fd_sc_hd__mux2_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _6857_/Q VGND VGND VPWR VPWR _5335_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5105_ _4620_/A _4595_/A _5263_/B _5104_/X VGND VGND VPWR VPWR _5105_/X sky130_fd_sc_hd__a31o_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6762_/Q _5771_/X _5788_/X _6747_/Q _6084_/X VGND VGND VPWR VPWR _6085_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1214 _6785_/Q VGND VGND VPWR VPWR _4176_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 _4000_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3297_ _7176_/Q _5757_/C _6803_/Q _7177_/Q VGND VGND VPWR VPWR _3297_/Y sky130_fd_sc_hd__nand4b_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 _6768_/Q VGND VGND VPWR VPWR _4146_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 _3947_/A1 VGND VGND VPWR VPWR hold469/A sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _5036_/A _5036_/B _5036_/C VGND VGND VPWR VPWR _5036_/X sky130_fd_sc_hd__and3_1
XFILLER_38_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1258 _3951_/A1 VGND VGND VPWR VPWR hold595/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _3961_/A1 VGND VGND VPWR VPWR hold637/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_409 _6935_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6987_ _7135_/CLK _6987_/D fanout588/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5938_ _6965_/Q _5770_/X _5793_/X _6989_/Q _5937_/X VGND VGND VPWR VPWR _5938_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5869_ _5869_/A _5869_/B _5869_/C _5869_/D VGND VGND VPWR VPWR _5869_/Y sky130_fd_sc_hd__nor4_1
XFILLER_181_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4229_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4637_/A sky130_fd_sc_hd__buf_6
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6497_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6504_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6509_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6483_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _3340_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6910_ _7053_/CLK _6910_/D fanout601/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6841_ _6967_/CLK _6841_/D fanout585/X VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6772_ _7248_/CLK _6772_/D fanout590/X VGND VGND VPWR VPWR _6772_/Q sky130_fd_sc_hd__dfrtp_1
X_3984_ hold998/X _6539_/A0 _3986_/S VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5723_ _7182_/Q _5782_/C _7183_/Q VGND VGND VPWR VPWR _5723_/X sky130_fd_sc_hd__and3b_4
X_5654_ _4049_/B hold256/X _5656_/S VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4605_ _4620_/B _4786_/B _4923_/A VGND VGND VPWR VPWR _4607_/B sky130_fd_sc_hd__and3_1
XFILLER_191_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5585_ _6549_/A0 hold994/X hold44/X VGND VGND VPWR VPWR _5585_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold300 _5388_/X VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _5380_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4536_ _5090_/A _5090_/B _4597_/B VGND VGND VPWR VPWR _4575_/B sky130_fd_sc_hd__and3_1
Xhold322 _6889_/Q VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _5389_/X VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold344 _6849_/Q VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold355 _4038_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _5353_/X VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7255_ _3340_/A1 _7255_/D fanout613/X VGND VGND VPWR VPWR _7255_/Q sky130_fd_sc_hd__dfrtp_4
X_4467_ _5060_/B _5060_/C _5044_/A _5128_/B VGND VGND VPWR VPWR _4469_/B sky130_fd_sc_hd__nand4_1
Xhold377 _5498_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _5451_/X VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6206_ _6897_/Q _6129_/A _6122_/X _6889_/Q VGND VGND VPWR VPWR _6206_/X sky130_fd_sc_hd__a22o_1
Xhold399 _6779_/Q VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ _5476_/B _6536_/C _5273_/D VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__and3_2
XFILLER_132_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7186_ _7256_/CLK _7186_/D fanout594/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfstp_4
X_4398_ _4848_/A _4356_/A _4295_/A _4348_/X VGND VGND VPWR VPWR _4398_/X sky130_fd_sc_hd__a211o_2
Xhold1000 _6752_/Q VGND VGND VPWR VPWR _4126_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ _3349_/A _3349_/B VGND VGND VPWR VPWR _3349_/X sky130_fd_sc_hd__and2_2
X_6137_ _6143_/D _6141_/B _6138_/B _6425_/B VGND VGND VPWR VPWR _6137_/X sky130_fd_sc_hd__and4_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _5390_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _4032_/X VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1033 _6611_/Q VGND VGND VPWR VPWR _3944_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _6762_/Q VGND VGND VPWR VPWR _4138_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6068_ _6442_/S _7204_/Q _6443_/S _6067_/X VGND VGND VPWR VPWR _6068_/X sky130_fd_sc_hd__a211o_1
XFILLER_73_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1055 _6894_/Q VGND VGND VPWR VPWR _5376_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1066 _5683_/X VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1077 _7125_/Q VGND VGND VPWR VPWR _5637_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ _4597_/C _4786_/B _5263_/A _4606_/D _4561_/B VGND VGND VPWR VPWR _5222_/D
+ sky130_fd_sc_hd__o2111ai_1
Xhold1088 _4101_/X VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 _6729_/Q VGND VGND VPWR VPWR _4099_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _5795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_217 _4049_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _3918_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_239 hold2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5370_ hold380/X _3916_/C _5376_/S VGND VGND VPWR VPWR _5370_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4321_ _4754_/B _4255_/A _4698_/A _4970_/D _4722_/A VGND VGND VPWR VPWR _4321_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7040_ _7114_/CLK _7040_/D fanout604/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfstp_2
X_4252_ _4427_/D _4320_/A _4657_/C VGND VGND VPWR VPWR _4252_/Y sky130_fd_sc_hd__o21ai_1
X_4183_ hold320/X _4049_/X _4187_/S VGND VGND VPWR VPWR _4183_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6824_ _6828_/CLK _6824_/D fanout573/X VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_90_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6755_ _6768_/CLK _6755_/D fanout576/X VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3967_ _3875_/Y _3967_/A1 _3968_/S VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__mux2_1
X_5706_ _7177_/Q _7176_/Q _7178_/Q _5706_/D VGND VGND VPWR VPWR _5708_/B sky130_fd_sc_hd__nand4_1
X_6686_ _7278_/CLK _6686_/D fanout595/X VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3898_ _6836_/Q _5325_/C _5311_/C input10/X _3469_/X VGND VGND VPWR VPWR _3898_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_109_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5637_ _5637_/A0 _4051_/X _5637_/S VGND VGND VPWR VPWR _5637_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5568_ _3915_/B hold270/X _5574_/S VGND VGND VPWR VPWR _5568_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold130 _6841_/Q VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7307_ _7307_/A VGND VGND VPWR VPWR _7307_/X sky130_fd_sc_hd__clkbuf_2
Xhold141 _5320_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4519_ _4620_/A _4595_/A _4519_/C VGND VGND VPWR VPWR _4607_/A sky130_fd_sc_hd__and3_1
Xhold152 _5528_/X VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 hold163/A VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ hold91/X hold5/X _5502_/S VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__mux2_1
Xhold174 _6700_/Q VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _5519_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7238_ _3340_/A1 _7238_/D fanout613/X VGND VGND VPWR VPWR _7238_/Q sky130_fd_sc_hd__dfrtp_4
Xhold196 _7278_/Q VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout610 fanout611/X VGND VGND VPWR VPWR fanout610/X sky130_fd_sc_hd__buf_8
Xfanout621 input124/X VGND VGND VPWR VPWR _4494_/C sky130_fd_sc_hd__buf_4
X_7169_ _7170_/CLK hold3/X fanout605/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4870_ _4987_/B _4870_/B _4870_/C VGND VGND VPWR VPWR _5255_/C sky130_fd_sc_hd__and3_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3821_ _7156_/Q _3550_/X _3559_/X _6908_/Q VGND VGND VPWR VPWR _3821_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6540_ _6540_/A0 hold615/X _6541_/S VGND VGND VPWR VPWR _6540_/X sky130_fd_sc_hd__mux2_1
X_3752_ _3752_/A _3752_/B _3752_/C VGND VGND VPWR VPWR _3752_/Y sky130_fd_sc_hd__nand3_2
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6471_ _7256_/D _3321_/B _6470_/Y _6471_/B2 VGND VGND VPWR VPWR _7220_/D sky130_fd_sc_hd__a22o_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3683_ _6685_/Q _4029_/B _5350_/B _6873_/Q VGND VGND VPWR VPWR _3683_/X sky130_fd_sc_hd__a22o_1
X_5422_ _6524_/B _6530_/D _5548_/D _5422_/D VGND VGND VPWR VPWR _5430_/S sky130_fd_sc_hd__nand4_4
XFILLER_145_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 _3251_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 _3336_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
XFILLER_173_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput224 _7296_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
Xoutput235 _7306_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
X_5353_ _3918_/B hold365/X _5358_/S VGND VGND VPWR VPWR _5353_/X sky130_fd_sc_hd__mux2_1
Xoutput246 _7286_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
XFILLER_114_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput257 _6826_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
Xoutput268 _6823_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
X_4304_ _4754_/B _4255_/A _4494_/C _4557_/A _4647_/C VGND VGND VPWR VPWR _4304_/Y
+ sky130_fd_sc_hd__o2111ai_4
Xoutput279 _6830_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
X_5284_ hold405/X _6538_/A0 _5287_/S VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__mux2_1
X_7023_ _7072_/CLK _7023_/D fanout599/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4235_ _4235_/A _4235_/B VGND VGND VPWR VPWR _4310_/C sky130_fd_sc_hd__nor2_2
XFILLER_101_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4166_ _7255_/Q _4166_/B VGND VGND VPWR VPWR _4206_/B sky130_fd_sc_hd__nand2b_4
XFILLER_67_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4097_ _5494_/A _3571_/X _3918_/X _4102_/S _4097_/B2 VGND VGND VPWR VPWR _4097_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6807_ _7254_/CLK _6807_/D _6472_/A VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4999_ _4999_/A1 _4722_/A _4984_/A _4662_/C _4722_/Y VGND VGND VPWR VPWR _4999_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_149_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6738_ _6855_/CLK _6738_/D fanout584/X VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__dfstp_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6669_ _7244_/CLK _6669_/D fanout576/X VGND VGND VPWR VPWR _6669_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout462 _5273_/D VGND VGND VPWR VPWR _5494_/C sky130_fd_sc_hd__clkbuf_16
Xfanout473 _5630_/C VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__buf_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout484 _6543_/A0 VGND VGND VPWR VPWR _5667_/A0 sky130_fd_sc_hd__buf_6
Xfanout495 _3987_/A VGND VGND VPWR VPWR _6524_/A sky130_fd_sc_hd__buf_12
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4020_ _4017_/B _3919_/X _4021_/S hold967/X VGND VGND VPWR VPWR _4020_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5971_ _7078_/Q _5971_/A2 _5813_/X _7062_/Q _5970_/X VGND VGND VPWR VPWR _5971_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4922_ _4922_/A _4922_/B _4922_/C VGND VGND VPWR VPWR _4925_/D sky130_fd_sc_hd__nor3_1
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4853_ _4984_/B _4984_/C _4853_/C _4903_/B VGND VGND VPWR VPWR _4865_/D sky130_fd_sc_hd__nand4_1
XFILLER_60_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3804_ _6891_/Q _3445_/X _3550_/X _7155_/Q _3803_/X VGND VGND VPWR VPWR _3804_/X
+ sky130_fd_sc_hd__a221o_1
X_4784_ _4550_/Y _5248_/A3 _4707_/Y _4783_/X VGND VGND VPWR VPWR _4784_/X sky130_fd_sc_hd__o31a_1
XFILLER_165_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6523_ _3925_/C hold396/X _6523_/S VGND VGND VPWR VPWR _6523_/X sky130_fd_sc_hd__mux2_1
X_3735_ _6600_/Q _3927_/B _5593_/B _7090_/Q _3734_/X VGND VGND VPWR VPWR _3735_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6454_ _6662_/Q _6129_/B _6454_/B1 _6772_/Q _6453_/X VGND VGND VPWR VPWR _6454_/X
+ sky130_fd_sc_hd__a221o_1
X_3666_ _6735_/Q _5341_/A _5311_/C _3571_/X _6727_/Q VGND VGND VPWR VPWR _3666_/X
+ sky130_fd_sc_hd__a32o_1
X_5405_ _5649_/A0 hold917/X _5412_/S VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__mux2_1
X_6385_ _6749_/Q _6098_/X _6105_/X _6603_/Q VGND VGND VPWR VPWR _6385_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3597_ _6849_/Q _5323_/S _3544_/X _6944_/Q _3596_/X VGND VGND VPWR VPWR _3597_/X
+ sky130_fd_sc_hd__a221o_2
X_5336_ _6550_/A0 hold735/X _5340_/S VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5267_ _5217_/X _5266_/Y _5235_/X _5262_/Y VGND VGND VPWR VPWR _5267_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_85_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7006_ _7006_/CLK _7006_/D fanout603/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfrtp_2
X_4218_ _4229_/A _4229_/B _4698_/A _4657_/C VGND VGND VPWR VPWR _4219_/B sky130_fd_sc_hd__nand4_1
X_5198_ _4751_/A _4294_/B _5128_/A _5197_/Y VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__a31o_1
XFILLER_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4149_ hold639/X _6546_/A0 _4150_/S VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3520_ _6597_/Q _6530_/C _3466_/X _5377_/C _6895_/Q VGND VGND VPWR VPWR _3523_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_7_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap415 _6108_/X VGND VGND VPWR VPWR _6465_/A3 sky130_fd_sc_hd__buf_12
XFILLER_128_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold707 hold707/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
XFILLER_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold718 _6932_/Q VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _7240_/Q VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap437 _4804_/A VGND VGND VPWR VPWR _4801_/B sky130_fd_sc_hd__clkbuf_1
Xmax_cap448 _5295_/D VGND VGND VPWR VPWR _5279_/D sky130_fd_sc_hd__clkbuf_2
X_3451_ _6854_/Q _5311_/B _5327_/D _3907_/B _6587_/Q VGND VGND VPWR VPWR _3451_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3382_ _6539_/A0 hold979/X _3384_/S VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__mux2_1
X_6170_ _6984_/Q _6098_/X _6129_/C _7152_/Q _6169_/X VGND VGND VPWR VPWR _6181_/A
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_3_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7274_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _5194_/B _5258_/A _5121_/C _5121_/D VGND VGND VPWR VPWR _5125_/A sky130_fd_sc_hd__and4_1
Xhold1407 _7055_/Q VGND VGND VPWR VPWR hold1407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 _6835_/Q VGND VGND VPWR VPWR hold115/A sky130_fd_sc_hd__dlygate4sd3_1
X_5052_ _5060_/C _5260_/B _5260_/C _5051_/X VGND VGND VPWR VPWR _5052_/X sky130_fd_sc_hd__a31o_1
XFILLER_85_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1429 _6584_/Q VGND VGND VPWR VPWR _3845_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4003_ _6546_/A0 hold488/X _4003_/S VGND VGND VPWR VPWR _4003_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5954_ _6292_/S _5954_/A2 _6343_/S VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4905_ _4597_/B _5263_/A _4557_/X _4903_/B _4774_/B VGND VGND VPWR VPWR _4907_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5885_ _6292_/S _7196_/Q _6443_/S _5884_/X VGND VGND VPWR VPWR _5885_/X sky130_fd_sc_hd__a211o_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4836_ _4344_/Y _4349_/X _4466_/X _4299_/Y _4835_/X VGND VGND VPWR VPWR _4836_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4767_ _4598_/Y _4645_/Y _4743_/Y _4635_/Y _4766_/Y VGND VGND VPWR VPWR _4767_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_21_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6506_ _7259_/Q _6506_/A2 _6506_/B1 _7257_/Q VGND VGND VPWR VPWR _6506_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3718_ _6736_/Q _5341_/A _5311_/C _3531_/X _6756_/Q VGND VGND VPWR VPWR _3718_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4698_ _4698_/A _4699_/B _4870_/B VGND VGND VPWR VPWR _4923_/C sky130_fd_sc_hd__and3_4
X_6437_ _6651_/Q _6177_/A _6106_/C _6143_/X _6776_/Q VGND VGND VPWR VPWR _6437_/X
+ sky130_fd_sc_hd__a32o_1
X_3649_ _6594_/Q _3913_/B _3503_/X _7137_/Q _3573_/X VGND VGND VPWR VPWR _3649_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6368_ _6367_/X _6392_/B1 _6443_/S VGND VGND VPWR VPWR _6368_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5319_ _3919_/C hold284/X _5322_/S VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6299_ _7165_/Q _6444_/B _6138_/B _6137_/X _7101_/Q VGND VGND VPWR VPWR _6299_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold12 hold7/X VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__buf_6
XFILLER_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold23 hold49/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold34 hold34/A VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__buf_6
XFILLER_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__buf_8
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_9 _3368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7254_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5674_/S hold876/X _3550_/X _3922_/X VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4621_ _4620_/X _4619_/X _4618_/Y _4516_/A VGND VGND VPWR VPWR _4621_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4552_ _5263_/A _4923_/B VGND VGND VPWR VPWR _4552_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold504 _6689_/Q VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 _6681_/Q VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _5666_/C _5575_/C _5575_/D VGND VGND VPWR VPWR _3503_/X sky130_fd_sc_hd__and3_4
X_7271_ _7271_/CLK _7271_/D fanout597/X VGND VGND VPWR VPWR _7271_/Q sky130_fd_sc_hd__dfrtp_4
Xhold526 hold526/A VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4483_ _4600_/B _4860_/B _4801_/A _5128_/B VGND VGND VPWR VPWR _4484_/D sky130_fd_sc_hd__a31o_1
XFILLER_171_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold537 _6546_/X VGND VGND VPWR VPWR _7273_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold548 hold548/A VGND VGND VPWR VPWR hold548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _7074_/Q VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ _7162_/Q _6444_/B _6465_/A2 _6116_/X hold52/A VGND VGND VPWR VPWR _6222_/X
+ sky130_fd_sc_hd__a32o_1
X_3434_ _5476_/C _5327_/D _6536_/D VGND VGND VPWR VPWR _3434_/X sky130_fd_sc_hd__and3_1
XFILLER_143_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6153_ _7095_/Q _6138_/B _5750_/C _6150_/X _6152_/X VGND VGND VPWR VPWR _6153_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _6546_/A0 hold524/X _3366_/S VGND VGND VPWR VPWR _3365_/X sky130_fd_sc_hd__mux2_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5104_ _4333_/A _4786_/B _5036_/X _4549_/D _4615_/X VGND VGND VPWR VPWR _5104_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6601_/Q _6025_/B _6028_/B _5789_/X _6782_/Q VGND VGND VPWR VPWR _6084_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _5335_/X VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _7176_/Q _5757_/C _7177_/Q VGND VGND VPWR VPWR _3296_/Y sky130_fd_sc_hd__nand3b_1
Xhold1215 _4176_/X VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _6717_/Q VGND VGND VPWR VPWR _4079_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _4146_/X VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _3569_/A1 VGND VGND VPWR VPWR hold526/A sky130_fd_sc_hd__dlygate4sd3_1
X_5035_ _5089_/A _5263_/B _5089_/B _4333_/A _5034_/Y VGND VGND VPWR VPWR _5035_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1259 _3633_/A1 VGND VGND VPWR VPWR hold585/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6986_ _7145_/CLK _6986_/D fanout600/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5937_ _6981_/Q _6073_/B2 _5774_/X _6909_/Q _5935_/X VGND VGND VPWR VPWR _5937_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5868_ _6962_/Q _5770_/X _5794_/X _6922_/Q _5867_/X VGND VGND VPWR VPWR _5869_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4819_ _4738_/B _4597_/C _5143_/A _5260_/A _5260_/B VGND VGND VPWR VPWR _4832_/B
+ sky130_fd_sc_hd__o2111ai_1
X_5799_ _6975_/Q _6073_/B2 _5771_/X _6967_/Q VGND VGND VPWR VPWR _5799_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4228_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4747_/C sky130_fd_sc_hd__buf_4
XFILLER_49_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR input124/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6500_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6506_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6498_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6514_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _6976_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6751_/CLK sky130_fd_sc_hd__clkbuf_16
X_6840_ _7071_/CLK hold41/X fanout585/X VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6771_ _6812_/CLK _6771_/D fanout580/X VGND VGND VPWR VPWR _6771_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_16_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3983_ hold789/X _6550_/A0 _3986_/S VGND VGND VPWR VPWR _3983_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5722_ _7182_/Q _7183_/Q VGND VGND VPWR VPWR _6010_/D sky130_fd_sc_hd__and2b_4
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_csclk _7277_/CLK VGND VGND VPWR VPWR _7245_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5653_ hold13/X _3503_/X _3924_/X _5656_/S hold809/X VGND VGND VPWR VPWR _5653_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_136_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4604_ _4604_/A _4604_/B _4604_/C VGND VGND VPWR VPWR _4607_/D sky130_fd_sc_hd__nand3_1
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5584_ _5630_/A _6548_/B _5675_/D _5657_/D VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__nand4_4
XFILLER_163_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7163_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold301 _6695_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4535_ _4544_/A _4544_/B _4606_/D _4544_/D VGND VGND VPWR VPWR _4535_/Y sky130_fd_sc_hd__nand4_2
Xhold312 _6839_/Q VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _5371_/X VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _6561_/Q VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold345 _5322_/X VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7254_ _7254_/CLK _7254_/D fanout613/X VGND VGND VPWR VPWR _7254_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4466_ _4356_/A _4848_/A _4259_/Y _4295_/A _4348_/X VGND VGND VPWR VPWR _4466_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_144_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold356 _6882_/Q VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _7092_/Q VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _6556_/Q VGND VGND VPWR VPWR hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 _6609_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ _6205_/A _6205_/B _6205_/C _6205_/D VGND VGND VPWR VPWR _6215_/B sky130_fd_sc_hd__nor4_4
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3417_ _6778_/Q _5311_/B _4158_/D VGND VGND VPWR VPWR _3417_/X sky130_fd_sc_hd__and3_1
X_7185_ _7251_/CLK _7185_/D fanout594/X VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfstp_4
X_4397_ _5042_/A _5060_/C _5042_/B VGND VGND VPWR VPWR _4399_/C sky130_fd_sc_hd__and3_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6136_/A _6425_/B _6177_/C VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__and3_4
X_3348_ _6851_/Q _6898_/Q _3346_/D _6882_/Q VGND VGND VPWR VPWR _3348_/Y sky130_fd_sc_hd__o31ai_2
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _4126_/X VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1012 _6683_/Q VGND VGND VPWR VPWR _4030_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _6559_/Q VGND VGND VPWR VPWR _3373_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ _6691_/Q _5726_/Y _6056_/X _6066_/X _5759_/A VGND VGND VPWR VPWR _6067_/X
+ sky130_fd_sc_hd__o221a_1
Xhold1034 _3944_/X VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 _4138_/X VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3279_ _6922_/Q VGND VGND VPWR VPWR _3279_/Y sky130_fd_sc_hd__inv_2
Xhold1056 _5376_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 _7078_/Q VGND VGND VPWR VPWR _5583_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5018_ _4620_/B _5263_/A _5017_/X _4900_/X VGND VGND VPWR VPWR _5020_/C sky130_fd_sc_hd__a31oi_2
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1078 _5637_/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 _7123_/Q VGND VGND VPWR VPWR _5635_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_207 _5313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _6535_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _6538_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _7067_/CLK hold36/X fanout582/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold890 _7260_/Q VGND VGND VPWR VPWR hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4320_ _4320_/A _4320_/B _4940_/C VGND VGND VPWR VPWR _4320_/Y sky130_fd_sc_hd__nor3_2
XFILLER_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4251_ _4427_/D _4320_/A _4249_/Y VGND VGND VPWR VPWR _4427_/A sky130_fd_sc_hd__o21ai_1
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4182_ _4182_/A0 _4181_/X _4188_/S VGND VGND VPWR VPWR _4182_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6823_ _6828_/CLK _6823_/D fanout573/X VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6754_ _7244_/CLK _6754_/D fanout581/X VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3966_ _3844_/Y _3966_/A1 _3968_/S VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5705_ _3307_/Y _5703_/Y _5704_/X _5697_/Y _7177_/Q VGND VGND VPWR VPWR _7177_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_188_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6685_ _7241_/CLK _6685_/D fanout576/X VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_2
X_3897_ _7078_/Q _3488_/X _5404_/B _6926_/Q _3896_/X VGND VGND VPWR VPWR _3904_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5636_ _6505_/A1 hold818/X hold29/X VGND VGND VPWR VPWR _5636_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5567_ _5667_/A0 _5567_/A1 _5574_/S VGND VGND VPWR VPWR _5567_/X sky130_fd_sc_hd__mux2_1
X_7306_ _7306_/A VGND VGND VPWR VPWR _7306_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold120 _5294_/X VGND VGND VPWR VPWR _6828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _5310_/X VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _4312_/A _4544_/D _4317_/Y _4388_/Y _4510_/Y VGND VGND VPWR VPWR _4518_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold142 _7035_/Q VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _7173_/Q VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ hold376/X _3921_/B _5502_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold164 _6972_/Q VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _4054_/X VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7237_ _7237_/CLK _7237_/D input164/X VGND VGND VPWR VPWR _7237_/Q sky130_fd_sc_hd__dfrtp_2
X_4449_ _4449_/A _4449_/B VGND VGND VPWR VPWR _4450_/B sky130_fd_sc_hd__nand2_1
Xhold186 _7041_/Q VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _6552_/X VGND VGND VPWR VPWR _7278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 input75/X VGND VGND VPWR VPWR fanout600/X sky130_fd_sc_hd__buf_6
Xfanout611 input75/X VGND VGND VPWR VPWR fanout611/X sky130_fd_sc_hd__buf_6
Xfanout622 _4729_/A VGND VGND VPWR VPWR _4612_/C sky130_fd_sc_hd__buf_12
X_7168_ _7168_/CLK _7168_/D fanout608/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfstp_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6119_ _6177_/A _6130_/A _6425_/B VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__and3_4
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7099_ _7099_/CLK _7099_/D fanout598/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _7084_/Q _3413_/X _5404_/B _6924_/Q _3819_/X VGND VGND VPWR VPWR _3825_/C
+ sky130_fd_sc_hd__a221o_1
X_3751_ _3751_/A _3751_/B _3751_/C _3751_/D VGND VGND VPWR VPWR _3752_/C sky130_fd_sc_hd__nor4_2
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ _7250_/Q _6470_/A2 _7249_/Q _7256_/Q _3321_/B VGND VGND VPWR VPWR _6470_/Y
+ sky130_fd_sc_hd__o41ai_1
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3682_ _6556_/Q _3359_/B _6542_/B _7272_/Q _3681_/X VGND VGND VPWR VPWR _3682_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5421_ _6511_/A1 hold428/X _5421_/S VGND VGND VPWR VPWR _5421_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput203 _3330_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_145_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput214 _7288_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
X_5352_ _6550_/A0 hold767/X _5358_/S VGND VGND VPWR VPWR _5352_/X sky130_fd_sc_hd__mux2_1
Xoutput225 _7297_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
XFILLER_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput236 _3331_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput247 _7287_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput258 _6827_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
X_4303_ _4549_/D _4255_/A _4600_/B _4557_/A _4647_/C VGND VGND VPWR VPWR _4310_/D
+ sky130_fd_sc_hd__o2111a_2
Xoutput269 _6824_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
X_5283_ _5283_/A0 _4152_/B _5287_/S VGND VGND VPWR VPWR _5283_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7022_ _7132_/CLK _7022_/D fanout611/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_114_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4234_ _4747_/A _4416_/A VGND VGND VPWR VPWR _4243_/A sky130_fd_sc_hd__nand2b_4
XFILLER_101_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4165_ _7255_/Q _7257_/Q _7258_/Q _7259_/Q VGND VGND VPWR VPWR _4165_/Y sky130_fd_sc_hd__nor4_2
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ _5494_/A _3571_/X _3915_/X _4102_/S _4096_/B2 VGND VGND VPWR VPWR _4096_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6806_ _3340_/A1 _6806_/D _6472_/A VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4998_ _4675_/A _4689_/A _4719_/B _4778_/C _4879_/C VGND VGND VPWR VPWR _5194_/A
+ sky130_fd_sc_hd__a221oi_2
X_6737_ _7239_/CLK _6737_/D fanout576/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfstp_2
X_3949_ _3753_/X _3949_/A1 _3953_/S VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6668_ _6780_/CLK _6668_/D fanout575/X VGND VGND VPWR VPWR _6668_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5619_ _5692_/A1 hold862/X _5619_/S VGND VGND VPWR VPWR _5619_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6599_ _6751_/CLK _6599_/D _3291_/A VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout430 _5714_/Y VGND VGND VPWR VPWR _5782_/C sky130_fd_sc_hd__buf_12
Xfanout452 hold28/X VGND VGND VPWR VPWR _5575_/D sky130_fd_sc_hd__buf_12
Xfanout463 _5485_/B VGND VGND VPWR VPWR _5273_/D sky130_fd_sc_hd__buf_12
XFILLER_59_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout474 _3385_/X VGND VGND VPWR VPWR _5630_/C sky130_fd_sc_hd__buf_12
Xfanout485 _6543_/A0 VGND VGND VPWR VPWR _6549_/A0 sky130_fd_sc_hd__buf_8
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout496 _3987_/A VGND VGND VPWR VPWR _5304_/A sky130_fd_sc_hd__buf_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5970_ _7046_/Q _5826_/B _5959_/B _5970_/B1 _6934_/Q VGND VGND VPWR VPWR _5970_/X
+ sky130_fd_sc_hd__a32o_1
X_4921_ _4746_/A _4939_/B _4778_/C _4582_/B VGND VGND VPWR VPWR _4922_/C sky130_fd_sc_hd__a31o_1
X_4852_ _5255_/A _5128_/B _4982_/D VGND VGND VPWR VPWR _4852_/X sky130_fd_sc_hd__and3_1
XANTENNA_390 _6446_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3803_ _7316_/A _5684_/B _3446_/X _3503_/X _7139_/Q VGND VGND VPWR VPWR _3803_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4783_ _4598_/Y _4701_/Y _4707_/Y _4743_/Y _4782_/Y VGND VGND VPWR VPWR _4783_/X
+ sky130_fd_sc_hd__o221a_1
X_6522_ _6540_/A0 hold664/X _6523_/S VGND VGND VPWR VPWR _6522_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3734_ _6572_/Q _6548_/A _5341_/A _3565_/X _6651_/Q VGND VGND VPWR VPWR _3734_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6453_ _6762_/Q _6097_/X _6143_/X _6777_/Q _6452_/X VGND VGND VPWR VPWR _6453_/X
+ sky130_fd_sc_hd__a221o_1
X_3665_ _6755_/Q _3531_/X _3663_/X _3664_/X VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__a211o_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5404_ _6542_/A _5404_/B VGND VGND VPWR VPWR _5412_/S sky130_fd_sc_hd__nand2_8
XFILLER_106_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6384_ _7245_/Q _6103_/X _6454_/B1 _6769_/Q _6383_/X VGND VGND VPWR VPWR _6389_/B
+ sky130_fd_sc_hd__a221o_1
X_3596_ _6968_/Q _5449_/B _5476_/C _5494_/C _3595_/X VGND VGND VPWR VPWR _3596_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5335_ _6549_/A0 _5335_/A1 _5340_/S VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5266_ _5266_/A _5266_/B _5266_/C VGND VGND VPWR VPWR _5266_/Y sky130_fd_sc_hd__nand3_1
XFILLER_87_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7005_ _7088_/CLK _7005_/D fanout590/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_1
X_4217_ _4662_/B _4870_/B VGND VGND VPWR VPWR _4363_/A sky130_fd_sc_hd__nor2_1
X_5197_ _5191_/Y _5197_/B _5197_/C VGND VGND VPWR VPWR _5197_/Y sky130_fd_sc_hd__nand3b_1
X_4148_ hold417/X _3919_/C _4150_/S VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4079_ _4079_/A0 _4078_/X _4093_/S VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7259_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap416 _6102_/X VGND VGND VPWR VPWR _6106_/C sky130_fd_sc_hd__buf_8
XFILLER_156_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold708 _7115_/Q VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold719 _5419_/X VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3450_ _3987_/A _5620_/A _5512_/B VGND VGND VPWR VPWR _3907_/B sky130_fd_sc_hd__and3_4
Xmax_cap449 _3528_/C VGND VGND VPWR VPWR _5295_/D sky130_fd_sc_hd__buf_2
XFILLER_143_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3381_ hold89/X _3381_/A1 _3384_/S VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__mux2_1
X_5120_ _5120_/A _5120_/B _5120_/C VGND VGND VPWR VPWR _5258_/B sky130_fd_sc_hd__and3_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5051_ _4460_/B _5143_/C _5140_/B _5050_/X _5049_/Y VGND VGND VPWR VPWR _5051_/X
+ sky130_fd_sc_hd__a311o_1
Xhold1408 _5558_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1419 _6577_/Q VGND VGND VPWR VPWR hold239/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4002_ _4003_/S hold791/X _3447_/X _3919_/X VGND VGND VPWR VPWR _4002_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5953_ _6877_/Q _5726_/Y _5939_/X _5952_/X _3246_/Y VGND VGND VPWR VPWR _5953_/X
+ sky130_fd_sc_hd__o221a_1
X_4904_ _5040_/C _4529_/X _4535_/Y _4552_/Y _4663_/Y VGND VGND VPWR VPWR _4907_/A
+ sky130_fd_sc_hd__o32ai_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5884_ _5726_/Y _6874_/Q _5759_/A _5883_/Y VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__o211a_1
XFILLER_178_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4835_ _4259_/Y _4358_/X _5040_/A _4814_/Y _4834_/X VGND VGND VPWR VPWR _4835_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_178_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4766_ _4923_/B _4682_/B _4765_/Y VGND VGND VPWR VPWR _4766_/Y sky130_fd_sc_hd__a21oi_1
X_3717_ _3717_/A _3717_/B _3717_/C _3717_/D VGND VGND VPWR VPWR _3717_/Y sky130_fd_sc_hd__nor4_1
X_6505_ _6504_/X _6505_/A1 _6511_/S VGND VGND VPWR VPWR _7234_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _4879_/A _4697_/B _4697_/C VGND VGND VPWR VPWR _4697_/Y sky130_fd_sc_hd__nor3_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6436_ _6681_/Q _6122_/X _6126_/X _6766_/Q VGND VGND VPWR VPWR _6436_/X sky130_fd_sc_hd__a22o_1
X_3648_ _6576_/Q _3397_/B _3969_/C _6635_/Q _3647_/X VGND VGND VPWR VPWR _3648_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6367_ _6366_/X _7214_/Q _6442_/S VGND VGND VPWR VPWR _6367_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3579_ _6575_/Q _3397_/B _3539_/X input53/X _3578_/X VGND VGND VPWR VPWR _3579_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5318_ _5323_/S _3922_/X _5322_/S hold932/X VGND VGND VPWR VPWR _5318_/X sky130_fd_sc_hd__a22o_1
X_6298_ _7157_/Q _6129_/C _6112_/X _7109_/Q _6297_/X VGND VGND VPWR VPWR _6305_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__buf_12
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__buf_6
X_5249_ _5249_/A _5249_/B _5249_/C VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__and3_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold35 hold1/X VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold46 hold46/A VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _4620_/A _4620_/B _4620_/C VGND VGND VPWR VPWR _4620_/X sky130_fd_sc_hd__and3_1
XFILLER_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4551_ _5090_/A _5090_/B _4923_/B VGND VGND VPWR VPWR _4903_/A sky130_fd_sc_hd__and3_2
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3502_ _5304_/A _5630_/C _5422_/D VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__and3_4
X_7270_ _7270_/CLK _7270_/D fanout579/X VGND VGND VPWR VPWR _7270_/Q sky130_fd_sc_hd__dfrtp_4
Xhold505 _4037_/X VGND VGND VPWR VPWR _6689_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _4027_/X VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4482_/A _4482_/B _4482_/C VGND VGND VPWR VPWR _4482_/Y sky130_fd_sc_hd__nand3_1
Xhold527 hold527/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
Xhold538 hold538/A VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6906_/Q _6129_/D _6138_/X _7034_/Q _6220_/X VGND VGND VPWR VPWR _6221_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3433_ _6530_/D _5476_/C _5422_/D VGND VGND VPWR VPWR _3433_/X sky130_fd_sc_hd__and3_4
Xhold549 hold549/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XFILLER_103_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _7159_/Q _6104_/X _6130_/X _6927_/Q _6151_/X VGND VGND VPWR VPWR _6152_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3919_/C hold378/X _3366_/S VGND VGND VPWR VPWR _3364_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _4333_/A _5089_/B _5102_/Y _5089_/X _5101_/Y VGND VGND VPWR VPWR _5103_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6657_/Q _5782_/X _6081_/X _6028_/C _6082_/X VGND VGND VPWR VPWR _6083_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _7178_/Q _7179_/Q VGND VGND VPWR VPWR _5757_/C sky130_fd_sc_hd__nor2_1
Xhold1205 _7290_/A VGND VGND VPWR VPWR _4182_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _6790_/Q VGND VGND VPWR VPWR _4186_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _4079_/X VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5034_ _5034_/A _5102_/A _5034_/C VGND VGND VPWR VPWR _5034_/Y sky130_fd_sc_hd__nand3_1
Xhold1238 _6818_/Q VGND VGND VPWR VPWR _5283_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1249 _3754_/A1 VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6985_ _7067_/CLK _6985_/D fanout582/X VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5936_ _5934_/C _6072_/C _6893_/Q _5776_/X _6957_/Q VGND VGND VPWR VPWR _5936_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5867_ _7026_/Q _5784_/X _5813_/X _7058_/Q VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4818_ _4349_/X _4356_/Y _4382_/Y _4398_/X _4815_/Y VGND VGND VPWR VPWR _5261_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_193_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5798_ _6959_/Q _5770_/X _5794_/X _6919_/Q _5797_/X VGND VGND VPWR VPWR _5798_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4799_/A _4748_/B _4747_/Y _4945_/C VGND VGND VPWR VPWR _4749_/X sky130_fd_sc_hd__a31o_1
XFILLER_107_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6419_ _6686_/Q _6101_/X _6454_/B1 _6771_/Q VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__a22o_1
XFILLER_122_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4228_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4747_/B sky130_fd_sc_hd__buf_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4706_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6503_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6510_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6501_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_stb_i VGND VGND VPWR VPWR _3313_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7270_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6770_ _6843_/CLK _6770_/D fanout581/X VGND VGND VPWR VPWR _6770_/Q sky130_fd_sc_hd__dfstp_2
X_3982_ hold874/X _6543_/A0 _3986_/S VGND VGND VPWR VPWR _3982_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5721_ _7181_/Q _7180_/Q _7182_/Q _7183_/Q VGND VGND VPWR VPWR _5721_/X sky130_fd_sc_hd__o31a_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5652_ hold13/X _3503_/X _3921_/X _5656_/S hold750/X VGND VGND VPWR VPWR _5652_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4603_ _4620_/C _4603_/B VGND VGND VPWR VPWR _4604_/C sky130_fd_sc_hd__nand2_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5583_ _5583_/A0 _5692_/A1 hold18/X VGND VGND VPWR VPWR _5583_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4534_ _4815_/A _4584_/B _5263_/A _4561_/B VGND VGND VPWR VPWR _4560_/C sky130_fd_sc_hd__nand4_1
Xhold302 _4046_/X VGND VGND VPWR VPWR _6695_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold313 _5308_/X VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _7106_/Q VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _3375_/X VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold346 _6864_/Q VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__dlygate4sd3_1
X_7253_ _7256_/CLK _7253_/D _6472_/A VGND VGND VPWR VPWR _7253_/Q sky130_fd_sc_hd__dfrtp_2
X_4465_ _4465_/A _4465_/B _4465_/C VGND VGND VPWR VPWR _4469_/A sky130_fd_sc_hd__nor3_1
Xhold357 _5363_/X VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _5599_/X VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ _6921_/Q _6129_/B _6129_/D _6905_/Q _6203_/X VGND VGND VPWR VPWR _6205_/D
+ sky130_fd_sc_hd__a221o_2
Xhold379 _3364_/X VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ hold54/X hold75/X hold16/X _5324_/B VGND VGND VPWR VPWR _3542_/B sky130_fd_sc_hd__and4bb_4
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7184_ _7256_/CLK _7184_/D fanout594/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4396_ _5055_/D _5143_/A _4449_/B VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__and3_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6141_/B _6138_/B _6143_/C _6143_/D VGND VGND VPWR VPWR _6135_/X sky130_fd_sc_hd__and4b_4
X_3347_ hold64/A _3347_/A2 _3346_/Y _3347_/B2 VGND VGND VPWR VPWR _3347_/X sky130_fd_sc_hd__a22o_2
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _6750_/Q VGND VGND VPWR VPWR _4124_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 _4030_/X VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 _3373_/X VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6066_ _6656_/Q _5782_/X _6058_/X _6060_/X _6065_/X VGND VGND VPWR VPWR _6066_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1035 hold1279/X VGND VGND VPWR VPWR hold1035/X sky130_fd_sc_hd__dlygate4sd3_1
X_3278_ _6930_/Q VGND VGND VPWR VPWR _3278_/Y sky130_fd_sc_hd__inv_2
Xhold1046 _7158_/Q VGND VGND VPWR VPWR _5674_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 _7006_/Q VGND VGND VPWR VPWR _5502_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _4494_/C _4801_/A _4860_/B _4923_/B VGND VGND VPWR VPWR _5017_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1068 _5583_/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 _6863_/Q VGND VGND VPWR VPWR _5342_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _5313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 _3925_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6968_ _7071_/CLK _6968_/D fanout586/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfstp_2
X_5919_ _7012_/Q _5965_/B _5815_/B _5783_/C _5918_/X VGND VGND VPWR VPWR _5919_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_179_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6899_ _7073_/CLK _6899_/D fanout585/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 _6595_/Q VGND VGND VPWR VPWR hold880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _6531_/X VGND VGND VPWR VPWR _7260_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4250_ _4761_/C _4209_/Y _4320_/A _4249_/Y VGND VGND VPWR VPWR _4383_/A sky130_fd_sc_hd__o31a_4
XFILLER_4_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4181_ hold369/X _3924_/X _4187_/S VGND VGND VPWR VPWR _4181_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6822_ _7265_/CLK _6822_/D fanout575/X VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6753_ _6828_/CLK _6753_/D fanout573/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfrtp_2
X_3965_ _3965_/A0 _3965_/A1 _3968_/S VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__mux2_1
X_5704_ _6803_/Q _6442_/S _7177_/Q _7176_/Q VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6684_ _7248_/CLK _6684_/D fanout580/X VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_2
X_3896_ _7110_/Q _6548_/A _5684_/C _3413_/X _7086_/Q VGND VGND VPWR VPWR _3896_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5635_ _5635_/A0 _3924_/X _5637_/S VGND VGND VPWR VPWR _5635_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5566_ _6542_/A _5566_/B VGND VGND VPWR VPWR _5574_/S sky130_fd_sc_hd__nand2_8
Xhold110 _6922_/Q VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _6866_/Q VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7305_ _7305_/A VGND VGND VPWR VPWR _7305_/X sky130_fd_sc_hd__clkbuf_2
Xhold132 _7101_/Q VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4517_ _4620_/B _4517_/B _5090_/B VGND VGND VPWR VPWR _5036_/A sky130_fd_sc_hd__and3_2
X_5497_ hold81/X hold2/X _5502_/S VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold143 _5535_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _5691_/X VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _5464_/X VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _7013_/Q VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlygate4sd3_1
X_7236_ _3340_/A1 _7236_/D input164/X VGND VGND VPWR VPWR _7236_/Q sky130_fd_sc_hd__dfrtp_2
X_4448_ _4860_/C _4449_/A _5260_/B _4447_/Y VGND VGND VPWR VPWR _4450_/A sky130_fd_sc_hd__a31oi_1
Xfanout601 fanout603/X VGND VGND VPWR VPWR fanout601/X sky130_fd_sc_hd__buf_8
XFILLER_120_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold187 _5542_/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _6974_/Q VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 input164/X VGND VGND VPWR VPWR _6472_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout623 _4557_/A VGND VGND VPWR VPWR _4729_/A sky130_fd_sc_hd__buf_8
X_4379_ _5042_/A _5143_/D _5042_/B VGND VGND VPWR VPWR _4460_/B sky130_fd_sc_hd__and3_1
X_7167_ _7167_/CLK _7167_/D fanout604/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfstp_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6118_ _6130_/A _6136_/A _6425_/B VGND VGND VPWR VPWR _6118_/X sky130_fd_sc_hd__and3_4
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7130_/CLK hold51/X fanout600/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6776_/Q _5779_/X _5793_/X _6751_/Q _6048_/X VGND VGND VPWR VPWR _6049_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_97_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6781_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7096_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7117_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ _6676_/Q _4017_/B _5334_/B input64/X _3749_/X VGND VGND VPWR VPWR _3751_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3681_ _7262_/Q _6530_/C _5325_/C _5611_/B _7105_/Q VGND VGND VPWR VPWR _3681_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5420_ _5413_/B _4073_/X _5421_/S hold814/X VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput204 _3328_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
X_5351_ _5667_/A0 hold625/X _5358_/S VGND VGND VPWR VPWR _5351_/X sky130_fd_sc_hd__mux2_1
Xoutput215 _7289_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
Xoutput226 _7298_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
XFILLER_154_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput237 _3332_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
Xoutput248 _7309_/A VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
XFILLER_153_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4302_ _4494_/C _4557_/A _4647_/C VGND VGND VPWR VPWR _4320_/B sky130_fd_sc_hd__nand3_2
X_5282_ _6536_/B _5476_/C _5327_/D _6536_/D VGND VGND VPWR VPWR _5287_/S sky130_fd_sc_hd__and4_2
Xoutput259 _6828_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
XFILLER_153_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7021_ _7165_/CLK _7021_/D fanout601/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_2
X_4233_ _4427_/D _4235_/B VGND VGND VPWR VPWR _4236_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4164_ _7257_/Q _7258_/Q _7259_/Q VGND VGND VPWR VPWR _4164_/Y sky130_fd_sc_hd__nor3_4
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4095_ _4152_/B _4095_/A1 _4102_/S VGND VGND VPWR VPWR _4095_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6805_ _7254_/CLK _6805_/D _6472_/A VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4997_ _4997_/A _5257_/B _5109_/B VGND VGND VPWR VPWR _5003_/A sky130_fd_sc_hd__and3_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6736_ _7239_/CLK _6736_/D fanout574/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfstp_2
X_3948_ _3693_/Y _3948_/A1 _3953_/S VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6667_ _7239_/CLK _6667_/D fanout576/X VGND VGND VPWR VPWR _6667_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3879_ _7054_/Q _3548_/X _3550_/X _7158_/Q _3878_/X VGND VGND VPWR VPWR _3889_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5618_ hold21/X _5618_/A1 _5619_/S VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__mux2_1
X_6598_ _6761_/CLK _6598_/D fanout572/X VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5549_ _6549_/A0 _5549_/A1 _5556_/S VGND VGND VPWR VPWR _5549_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7251_/CLK sky130_fd_sc_hd__clkbuf_16
X_7219_ _7219_/CLK _7219_/D fanout577/X VGND VGND VPWR VPWR _7219_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout431 _5714_/Y VGND VGND VPWR VPWR _6010_/C sky130_fd_sc_hd__buf_8
Xfanout453 hold27/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__buf_12
Xfanout464 hold1436/X VGND VGND VPWR VPWR _5485_/B sky130_fd_sc_hd__buf_12
Xfanout475 hold76/X VGND VGND VPWR VPWR _6530_/C sky130_fd_sc_hd__buf_12
Xfanout486 _3361_/X VGND VGND VPWR VPWR _6543_/A0 sky130_fd_sc_hd__buf_8
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout497 hold1441/X VGND VGND VPWR VPWR _3987_/A sky130_fd_sc_hd__buf_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4920_ _4211_/X _4575_/B _4589_/C _4778_/C _4903_/A VGND VGND VPWR VPWR _4922_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ _4377_/X _4987_/A _4987_/B _4903_/B _4708_/A VGND VGND VPWR VPWR _4851_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_380 hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_391 _5773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3802_ _6606_/Q hold56/A _4139_/C _5458_/B hold61/A VGND VGND VPWR VPWR _3802_/X
+ sky130_fd_sc_hd__a32o_2
X_4782_ _4923_/C _4775_/B _4781_/X _4780_/Y VGND VGND VPWR VPWR _4782_/Y sky130_fd_sc_hd__a211oi_1
X_6521_ _6539_/A0 _6521_/A1 _6523_/S VGND VGND VPWR VPWR _6521_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3733_ _7010_/Q _5512_/B _5657_/D hold28/A _3732_/X VGND VGND VPWR VPWR _3733_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_159_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6452_ _6682_/Q _6122_/X _6452_/B1 _6757_/Q _6451_/X VGND VGND VPWR VPWR _6452_/X
+ sky130_fd_sc_hd__a221o_1
X_3664_ input97/X _5331_/C _3540_/B _5323_/S _6846_/Q VGND VGND VPWR VPWR _3664_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5403_ hold178/X _4053_/B _5403_/S VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3595_ _6774_/Q _5422_/D _5325_/C _3452_/X _6960_/Q VGND VGND VPWR VPWR _3595_/X
+ sky130_fd_sc_hd__a32o_1
X_6383_ _6593_/Q _6130_/A _6114_/X _6177_/X _6639_/Q VGND VGND VPWR VPWR _6383_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5334_ _6548_/B _5334_/B VGND VGND VPWR VPWR _5340_/S sky130_fd_sc_hd__nand2_4
X_5265_ _5265_/A _5265_/B _5265_/C _5265_/D VGND VGND VPWR VPWR _5266_/C sky130_fd_sc_hd__and4_1
XFILLER_87_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7004_ _7157_/CLK _7004_/D fanout592/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_4
X_4216_ _4229_/C _4229_/D _4228_/A _4228_/B VGND VGND VPWR VPWR _4219_/A sky130_fd_sc_hd__nand4_1
X_5196_ _4409_/C _4376_/Y _5225_/B wire358/X _5225_/C VGND VGND VPWR VPWR _5197_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_96_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4147_ hold528/X _6538_/A0 _4150_/S VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4078_ _5342_/A0 _5649_/A0 _4092_/S VGND VGND VPWR VPWR _4078_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6719_ _7143_/CLK _6719_/D fanout587/X VGND VGND VPWR VPWR _7282_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_165_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold709 _5625_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap439 _4799_/B VGND VGND VPWR VPWR _4792_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3380_ _3370_/B _3380_/A1 _3384_/S VGND VGND VPWR VPWR _3380_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5050_ _4738_/B _4597_/C _4838_/X _5260_/B _4449_/A VGND VGND VPWR VPWR _5050_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1409 _7252_/Q VGND VGND VPWR VPWR _7258_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4001_ _4003_/S hold884/X _3447_/X _3916_/X VGND VGND VPWR VPWR _4001_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3347_/B2
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5952_ _7101_/Q _5780_/X _5944_/X _5948_/X _5951_/X VGND VGND VPWR VPWR _5952_/X
+ sky130_fd_sc_hd__a2111o_1
X_4903_ _4903_/A _4903_/B VGND VGND VPWR VPWR _4903_/Y sky130_fd_sc_hd__nand2_1
X_5883_ _5883_/A _5883_/B VGND VGND VPWR VPWR _5883_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4834_ _4380_/X _4382_/Y _5040_/A _4816_/X _4833_/X VGND VGND VPWR VPWR _4834_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4765_ _4765_/A _4765_/B _4765_/C VGND VGND VPWR VPWR _4765_/Y sky130_fd_sc_hd__nand3_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6504_ _7257_/Q _6504_/A2 _6504_/B1 _4164_/Y _6503_/X VGND VGND VPWR VPWR _6504_/X
+ sky130_fd_sc_hd__a221o_1
X_3716_ _6610_/Q _3558_/X _3712_/X _3715_/X VGND VGND VPWR VPWR _3717_/D sky130_fd_sc_hd__a211o_1
X_4696_ _4939_/A _5255_/A _4878_/B _4878_/C VGND VGND VPWR VPWR _4697_/B sky130_fd_sc_hd__and4_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _7268_/Q _6106_/X _6119_/X _6590_/Q _6434_/X VGND VGND VPWR VPWR _6440_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3647_ _7145_/Q _5684_/B _3412_/X _3539_/X input54/X VGND VGND VPWR VPWR _3647_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6366_ _6356_/Y wire352/X _6688_/Q _6466_/A1 VGND VGND VPWR VPWR _6366_/X sky130_fd_sc_hd__o2bb2a_1
X_3578_ _6654_/Q _5341_/A _3542_/B _5377_/C _6896_/Q VGND VGND VPWR VPWR _3578_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5317_ hold5/X _5317_/A1 _5322_/S VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__mux2_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6297_ _7093_/Q _6136_/A _6106_/C _6144_/X _7085_/Q VGND VGND VPWR VPWR _6297_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__buf_6
X_5248_ _4344_/Y _5153_/X _5248_/A3 _4965_/X _5079_/C VGND VGND VPWR VPWR _5249_/C
+ sky130_fd_sc_hd__o311a_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold47 hold4/X VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5179_ _4208_/Y _4970_/A _4333_/Y _5178_/X VGND VGND VPWR VPWR _5180_/B sky130_fd_sc_hd__o31a_1
XFILLER_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4550_ _5036_/C _4755_/D VGND VGND VPWR VPWR _4550_/Y sky130_fd_sc_hd__nand2_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3501_ _6991_/Q _3496_/X _3497_/X _6823_/Q _3500_/X VGND VGND VPWR VPWR _3507_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold506 _6562_/Q VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlygate4sd3_1
X_4481_ _5040_/C _4244_/Y _4259_/Y _4356_/Y _5165_/C VGND VGND VPWR VPWR _4482_/C
+ sky130_fd_sc_hd__o41a_1
Xhold517 _6776_/Q VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 _6769_/Q VGND VGND VPWR VPWR hold528/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6220_ _6922_/Q _6129_/B _6451_/B1 _6914_/Q _6219_/X VGND VGND VPWR VPWR _6220_/X
+ sky130_fd_sc_hd__a221o_1
Xhold539 hold539/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
X_3432_ _6548_/C _5666_/C _5575_/C VGND VGND VPWR VPWR _3432_/X sky130_fd_sc_hd__and3_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ hold89/X _3363_/A1 _3366_/S VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__mux2_1
X_6151_ _7167_/Q _6130_/A _6114_/X _6107_/X _6999_/Q VGND VGND VPWR VPWR _6151_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A _5102_/B VGND VGND VPWR VPWR _5102_/Y sky130_fd_sc_hd__nand2_1
X_6082_ _6028_/C _5782_/C _5795_/C _5813_/X _6568_/Q VGND VGND VPWR VPWR _6082_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _7192_/Q _6844_/Q _6849_/Q VGND VGND VPWR VPWR _3307_/B sky130_fd_sc_hd__mux2_8
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _4182_/X VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _4186_/X VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _6663_/Q VGND VGND VPWR VPWR _4006_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5033_ _5033_/A _5033_/B VGND VGND VPWR VPWR _5034_/C sky130_fd_sc_hd__nor2_1
Xhold1239 _5283_/X VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6984_ _7163_/CLK _6984_/D fanout610/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_25_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5935_ _7037_/Q _6072_/B _6003_/C _5934_/X VGND VGND VPWR VPWR _5935_/X sky130_fd_sc_hd__a31o_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5866_ _7106_/Q _5764_/X _5776_/X _6954_/Q _5865_/X VGND VGND VPWR VPWR _5869_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4817_ _4299_/Y _4382_/Y _4395_/Y _4456_/B VGND VGND VPWR VPWR _4817_/X sky130_fd_sc_hd__o31a_1
XFILLER_166_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5797_ _7079_/Q _5826_/B _6009_/C _5796_/X VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__a31o_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4748_ _4799_/A _4748_/B VGND VGND VPWR VPWR _4752_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4679_ _4359_/Y _4372_/Y _4408_/X _4848_/B _4667_/Y VGND VGND VPWR VPWR _4681_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_135_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6418_ _6417_/X _6442_/A1 _6443_/S VGND VGND VPWR VPWR _6418_/X sky130_fd_sc_hd__mux2_1
X_6349_ _6663_/Q _6451_/B1 _6452_/B1 _6753_/Q VGND VGND VPWR VPWR _6349_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4228_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3316_/C sky130_fd_sc_hd__clkbuf_1
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR input126/X sky130_fd_sc_hd__clkbuf_1
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6507_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6488_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6504_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ _6542_/A _5273_/D _5325_/C VGND VGND VPWR VPWR _3986_/S sky130_fd_sc_hd__and3_4
X_5720_ _7183_/Q _7182_/Q VGND VGND VPWR VPWR _5720_/Y sky130_fd_sc_hd__nor2_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5651_ hold13/X _3503_/X _3918_/X _5656_/S hold756/X VGND VGND VPWR VPWR _5651_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_175_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4602_ _4214_/A _4214_/B _4517_/B _4544_/A _4510_/Y VGND VGND VPWR VPWR _4603_/B
+ sky130_fd_sc_hd__a2111oi_4
X_5582_ hold607/X _4051_/B hold18/X VGND VGND VPWR VPWR _5582_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4533_ _4597_/C _4561_/B _4581_/B VGND VGND VPWR VPWR _4562_/B sky130_fd_sc_hd__and3_1
XFILLER_144_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold303 hold303/A VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _7156_/Q VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold325 _5615_/X VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7252_ _7259_/CLK _7252_/D _6472_/A VGND VGND VPWR VPWR _7252_/Q sky130_fd_sc_hd__dfrtp_2
X_4464_ _4464_/A _4464_/B _4464_/C VGND VGND VPWR VPWR _4465_/C sky130_fd_sc_hd__nand3_1
Xhold336 _7122_/Q VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _5343_/X VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _6939_/Q VGND VGND VPWR VPWR hold358/X sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6913_/Q _6451_/B1 _6462_/B1 _6937_/Q VGND VGND VPWR VPWR _6203_/X sky130_fd_sc_hd__a22o_1
Xhold369 _6697_/Q VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlygate4sd3_1
X_3415_ _6838_/Q _3406_/X _4133_/B _6758_/Q _3414_/X VGND VGND VPWR VPWR _3415_/X
+ sky130_fd_sc_hd__a221o_1
X_7183_ _7259_/CLK _7183_/D fanout594/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_4
X_4395_ _5055_/D _5143_/A VGND VGND VPWR VPWR _4395_/Y sky130_fd_sc_hd__nand2_2
XFILLER_131_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6132_/Y _6121_/X _6134_/C _6134_/D VGND VGND VPWR VPWR _6134_/Y sky130_fd_sc_hd__nand4bb_4
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ hold64/A _6851_/Q _6898_/Q _3346_/D VGND VGND VPWR VPWR _3346_/Y sky130_fd_sc_hd__nor4_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1003 _4124_/X VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _7263_/Q _5777_/X _6061_/X _6062_/X _6064_/X VGND VGND VPWR VPWR _6065_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1014 _7298_/A VGND VGND VPWR VPWR _4205_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 _6554_/Q VGND VGND VPWR VPWR _3362_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3277_ _6938_/Q VGND VGND VPWR VPWR _3277_/Y sky130_fd_sc_hd__inv_2
Xhold1036 hold1036/A VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
Xhold1047 _5674_/X VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _5502_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5016_ _4549_/D _4600_/B _4860_/B _4298_/X VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__a31o_1
XFILLER_66_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1069 _7150_/Q VGND VGND VPWR VPWR _5665_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_209 _4127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _6967_/CLK _6967_/D fanout586/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5918_ _7084_/Q _5965_/B _6009_/C _5788_/X _6996_/Q VGND VGND VPWR VPWR _5918_/X
+ sky130_fd_sc_hd__a32o_1
X_6898_ _7143_/CLK _6898_/D fanout589/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5849_ _6881_/Q _5768_/X _5845_/X _5846_/X _5848_/X VGND VGND VPWR VPWR _5849_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold870 _7304_/A VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold881 _3923_/X VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold892 _6701_/Q VGND VGND VPWR VPWR hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__1184_ clkbuf_0__1184_/X VGND VGND VPWR VPWR _3965_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4180_ _4180_/A0 _4179_/X _4188_/S VGND VGND VPWR VPWR _4180_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6821_ _6827_/CLK _6821_/D fanout573/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6752_ _7269_/CLK _6752_/D fanout576/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3964_ _3753_/X _3964_/A1 _3968_/S VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5703_ _7177_/Q _7176_/Q VGND VGND VPWR VPWR _5703_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6683_ _7241_/CLK _6683_/D fanout576/X VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfrtp_2
X_3895_ _6894_/Q _3445_/X _3890_/X _3892_/X _3894_/X VGND VGND VPWR VPWR _3905_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_149_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5634_ _3921_/B hold336/X hold29/X VGND VGND VPWR VPWR _5634_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5565_ _4053_/B hold172/X _5565_/S VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__mux2_1
Xhold100 _7076_/Q VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__dlygate4sd3_1
X_7304_ _7304_/A VGND VGND VPWR VPWR _7304_/X sky130_fd_sc_hd__clkbuf_1
Xhold111 _5408_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4516_/A VGND VGND VPWR VPWR _4516_/Y sky130_fd_sc_hd__inv_2
Xhold122 _5345_/X VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ hold458/X _3916_/C _5502_/S VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold133 _5609_/X VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _6637_/Q VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _7065_/Q VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlygate4sd3_1
X_7235_ _3340_/A1 _7235_/D input164/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfrtp_2
Xhold166 _7049_/Q VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _4358_/X _4392_/Y _4435_/X _4380_/X _4446_/Y VGND VGND VPWR VPWR _4447_/Y
+ sky130_fd_sc_hd__o221ai_1
Xhold177 _5510_/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _6926_/Q VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _5466_/X VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 fanout603/X VGND VGND VPWR VPWR fanout602/X sky130_fd_sc_hd__buf_8
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout613 input164/X VGND VGND VPWR VPWR fanout613/X sky130_fd_sc_hd__buf_4
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7166_ _7173_/CLK _7166_/D fanout603/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout624 _4632_/B VGND VGND VPWR VPWR _4511_/A sky130_fd_sc_hd__buf_12
XFILLER_144_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4378_ _4859_/C _4704_/B _4862_/A VGND VGND VPWR VPWR _4465_/B sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_1_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7273_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6117_ _6117_/A _6130_/A _6117_/C VGND VGND VPWR VPWR _6117_/X sky130_fd_sc_hd__and3_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3329_/A _3350_/A VGND VGND VPWR VPWR _3329_/Y sky130_fd_sc_hd__nand2_2
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7097_/CLK _7097_/D fanout596/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6048_ _6766_/Q wire398/X _6028_/C _6557_/Q _5767_/X VGND VGND VPWR VPWR _6048_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3680_ _6561_/Q _3372_/B _3671_/X _3672_/X _3679_/X VGND VGND VPWR VPWR _3692_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5350_ hold12/X _5350_/B VGND VGND VPWR VPWR _5358_/S sky130_fd_sc_hd__nand2_8
Xoutput205 _3326_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput216 _7290_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
Xoutput227 _7299_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
Xoutput238 _7307_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
X_4301_ _4754_/B _4255_/A _4494_/C _4557_/A VGND VGND VPWR VPWR _4301_/Y sky130_fd_sc_hd__o211ai_4
Xoutput249 _7308_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
X_5281_ _5279_/D _5281_/A2 _3916_/X _5280_/S hold882/X VGND VGND VPWR VPWR _5281_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_99_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7020_ _7132_/CLK _7020_/D fanout610/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_4
X_4232_ _4698_/A _4657_/C _4656_/C VGND VGND VPWR VPWR _4235_/B sky130_fd_sc_hd__nand3_1
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4163_ _5311_/B _4158_/D _3925_/X _4162_/S hold915/X VGND VGND VPWR VPWR _4163_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4094_ _5311_/C _5476_/C _5630_/C _6524_/B VGND VGND VPWR VPWR _4102_/S sky130_fd_sc_hd__nand4_4
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6804_ _7254_/CLK _6804_/D _6472_/A VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfrtp_4
X_4996_ _5263_/C _4719_/B _5255_/C _4987_/C _4874_/X VGND VGND VPWR VPWR _5109_/B
+ sky130_fd_sc_hd__a221oi_1
X_6735_ _6828_/CLK _6735_/D fanout573/X VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3947_ _3632_/Y _3947_/A1 _3953_/S VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6666_ _7241_/CLK _6666_/D fanout575/X VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3878_ _7070_/Q _5566_/B _3499_/X _7022_/Q _3877_/X VGND VGND VPWR VPWR _3878_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5617_ _6505_/A1 hold805/X _5619_/S VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6597_ _6781_/CLK _6597_/D _3291_/A VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5548_ _5620_/A _6548_/B _5548_/C _5548_/D VGND VGND VPWR VPWR _5556_/S sky130_fd_sc_hd__nand4_4
XFILLER_145_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5479_ _3919_/C hold293/X _5484_/S VGND VGND VPWR VPWR _5479_/X sky130_fd_sc_hd__mux2_1
X_7218_ _7218_/CLK _7218_/D fanout577/X VGND VGND VPWR VPWR _7218_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout421 _5959_/B VGND VGND VPWR VPWR _6028_/B sky130_fd_sc_hd__buf_12
Xfanout432 _4638_/Y VGND VGND VPWR VPWR _5248_/A3 sky130_fd_sc_hd__clkbuf_8
Xfanout454 _3533_/C VGND VGND VPWR VPWR _4158_/D sky130_fd_sc_hd__buf_8
X_7149_ _7157_/CLK _7149_/D fanout593/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout465 _5548_/D VGND VGND VPWR VPWR _5476_/C sky130_fd_sc_hd__clkbuf_16
Xfanout476 hold76/A VGND VGND VPWR VPWR _3563_/A sky130_fd_sc_hd__buf_6
XFILLER_171_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout487 _6524_/B VGND VGND VPWR VPWR _6536_/B sky130_fd_sc_hd__buf_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4751_/A _4730_/D _4945_/B _4862_/A VGND VGND VPWR VPWR _4850_/X sky130_fd_sc_hd__o211a_1
XFILLER_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_370 _5815_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_381 hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 _5776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3801_ _6578_/Q _3987_/A _6548_/D _5684_/B _3757_/X VGND VGND VPWR VPWR _3801_/X
+ sky130_fd_sc_hd__a41o_1
X_4781_ _4923_/B _4939_/B _4923_/C VGND VGND VPWR VPWR _4781_/X sky130_fd_sc_hd__and3_1
XFILLER_33_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6520_ _6538_/A0 hold729/X _6523_/S VGND VGND VPWR VPWR _6520_/X sky130_fd_sc_hd__mux2_1
X_3732_ _7050_/Q _5512_/B _3540_/B _3562_/X _6641_/Q VGND VGND VPWR VPWR _3732_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6451_ _7264_/Q _6446_/C _6425_/C _6451_/B1 _6667_/Q VGND VGND VPWR VPWR _6451_/X
+ sky130_fd_sc_hd__a32o_1
X_3663_ _6750_/Q _5494_/C _3446_/X _5458_/B _6969_/Q VGND VGND VPWR VPWR _3663_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5402_ hold696/X _4051_/B _5403_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
X_6382_ _6555_/Q _6110_/X _6113_/X _6634_/Q _6381_/X VGND VGND VPWR VPWR _6389_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3594_ input96/X _5331_/C _3540_/B _5359_/B _6880_/Q VGND VGND VPWR VPWR _3594_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5333_ _6538_/A0 hold413/X _5333_/S VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5264_ _4576_/A _5263_/X _5264_/C _5264_/D VGND VGND VPWR VPWR _5265_/D sky130_fd_sc_hd__and4bb_1
XFILLER_141_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7003_ _7119_/CLK hold92/X fanout590/X VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__dfrtp_2
XFILLER_102_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4215_ _4637_/A _4747_/B _4747_/C VGND VGND VPWR VPWR _4742_/C sky130_fd_sc_hd__nor3_2
X_5195_ _4290_/Y _5040_/B _4715_/Y _4726_/Y _5127_/C VGND VGND VPWR VPWR _5225_/C
+ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_81_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _6843_/CLK sky130_fd_sc_hd__clkbuf_16
X_4146_ _4146_/A0 _4152_/B _4150_/S VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4077_ _4092_/S _3539_/X _4056_/Y _3387_/Y _4076_/X VGND VGND VPWR VPWR _4093_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_96_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7267_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4979_ _4516_/Y _4976_/Y _4978_/X _4896_/Y VGND VGND VPWR VPWR _4979_/X sky130_fd_sc_hd__o211a_1
XFILLER_149_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6718_ _7152_/CLK _6718_/D fanout587/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6649_ _7096_/CLK _6649_/D fanout596/X VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7170_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7133_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4000_ _4152_/B _4000_/A1 _4003_/S VGND VGND VPWR VPWR _4000_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5951_ _6973_/Q _5771_/X _5933_/X _5936_/X _5950_/X VGND VGND VPWR VPWR _5951_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4902_ _4620_/B _5263_/A _4901_/X _4900_/X VGND VGND VPWR VPWR _4909_/A sky130_fd_sc_hd__a31oi_1
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5882_ _5871_/X _5874_/X _5881_/X VGND VGND VPWR VPWR _5883_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4833_ _4382_/Y _4395_/Y _5040_/A _4817_/X _4832_/X VGND VGND VPWR VPWR _4833_/X
+ sky130_fd_sc_hd__o311a_1
X_4764_ _4730_/D _4939_/B _4755_/B _4763_/Y VGND VGND VPWR VPWR _4765_/C sky130_fd_sc_hd__a31oi_1
XFILLER_193_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6503_ _7259_/Q _6503_/A2 _6503_/B1 _7258_/Q VGND VGND VPWR VPWR _6503_/X sky130_fd_sc_hd__a22o_1
X_3715_ _6978_/Q _5485_/B _5281_/A2 _3714_/X VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__a31o_1
X_4695_ _4862_/A _4791_/B _4778_/C VGND VGND VPWR VPWR _4879_/A sky130_fd_sc_hd__and3_1
X_6434_ _6610_/Q _6138_/B _6465_/A3 _6107_/X _6814_/Q VGND VGND VPWR VPWR _6434_/X
+ sky130_fd_sc_hd__a32o_1
X_3646_ input5/X _4127_/C _5476_/C _5311_/C _3645_/X VGND VGND VPWR VPWR _3646_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6365_ _6365_/A _6365_/B _6440_/D _6365_/D VGND VGND VPWR VPWR _6365_/Y sky130_fd_sc_hd__nor4_1
XFILLER_127_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3577_ _7136_/Q _3503_/X _3521_/X _7168_/Q VGND VGND VPWR VPWR _3577_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5316_ _6524_/B _5323_/S VGND VGND VPWR VPWR _5322_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6296_ _7173_/Q _6117_/X _6177_/X _7021_/Q _6295_/X VGND VGND VPWR VPWR _6296_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5247_ _5247_/A _5247_/B _5247_/C VGND VGND VPWR VPWR _5247_/Y sky130_fd_sc_hd__nand3_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5178_/A _5266_/A _5220_/A VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__and3_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4129_ _6538_/A0 hold486/X _4132_/S VGND VGND VPWR VPWR _4129_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3500_ _6763_/Q _5494_/C _4139_/C _3499_/X _7015_/Q VGND VGND VPWR VPWR _3500_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4480_ _4689_/C _4480_/B VGND VGND VPWR VPWR _5165_/C sky130_fd_sc_hd__nand2_1
Xhold507 _3376_/X VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _4156_/X VGND VGND VPWR VPWR _6776_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _4147_/X VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3431_ _5324_/B hold26/X hold71/X _5657_/D VGND VGND VPWR VPWR _4139_/C sky130_fd_sc_hd__and4_4
XFILLER_143_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6150_ _7063_/Q _6103_/X _6110_/X _7111_/Q _6149_/X VGND VGND VPWR VPWR _6150_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _3370_/B _3362_/A1 _3366_/S VGND VGND VPWR VPWR _3362_/X sky130_fd_sc_hd__mux2_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5101_ _5101_/A _5220_/C VGND VGND VPWR VPWR _5101_/Y sky130_fd_sc_hd__nand2_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6682_/Q _5795_/C _5815_/C _6028_/B _6667_/Q VGND VGND VPWR VPWR _6081_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _7313_/A VGND VGND VPWR VPWR _3293_/Y sky130_fd_sc_hd__inv_2
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1207 _7288_/A VGND VGND VPWR VPWR _4178_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _4786_/B _4600_/Y _4606_/D _4620_/A _4606_/B VGND VGND VPWR VPWR _5033_/A
+ sky130_fd_sc_hd__o2111a_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 hold1366/X VGND VGND VPWR VPWR _4113_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1229 _4006_/X VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6983_ _7035_/CLK _6983_/D fanout590/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5934_ _6917_/Q _6028_/B _5934_/C VGND VGND VPWR VPWR _5934_/X sky130_fd_sc_hd__and3_1
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5865_ _7114_/Q _5965_/B _5842_/C _5814_/X _7050_/Q VGND VGND VPWR VPWR _5865_/X
+ sky130_fd_sc_hd__a32o_1
X_4816_ _4277_/Y _4382_/Y _4395_/Y _4815_/Y _4380_/X VGND VGND VPWR VPWR _4816_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_166_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5796_ _6999_/Q _5795_/D _6010_/C _5795_/C VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__o211a_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4747_ _4747_/A _4747_/B _4747_/C _4637_/A VGND VGND VPWR VPWR _4747_/Y sky130_fd_sc_hd__nor4b_2
XFILLER_193_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4678_ _4678_/A _4678_/B _4678_/C VGND VGND VPWR VPWR _4681_/A sky130_fd_sc_hd__nor3_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6417_ _6442_/S _7216_/Q _6415_/Y _6416_/X VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3629_ _6984_/Q _5485_/B _3540_/B _3628_/X VGND VGND VPWR VPWR _3629_/X sky130_fd_sc_hd__a31o_1
X_6348_ _6643_/Q _6177_/C _6112_/C _6462_/B1 _6653_/Q VGND VGND VPWR VPWR _6348_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4228_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6279_ _6972_/Q _6097_/X _6143_/X _6948_/Q _6278_/X VGND VGND VPWR VPWR _6279_/X
+ sky130_fd_sc_hd__a221o_1
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR _3317_/A sky130_fd_sc_hd__clkbuf_1
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4999_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6509_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6491_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ _3980_/A0 _6535_/A0 _3980_/S VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5650_ hold13/X _3503_/X _3915_/X _5656_/S hold744/X VGND VGND VPWR VPWR _5650_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4601_ _4754_/B _4633_/B _5036_/B VGND VGND VPWR VPWR _4601_/Y sky130_fd_sc_hd__nand3_4
X_5581_ hold100/X hold83/X hold18/X VGND VGND VPWR VPWR _5581_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _5090_/A _5090_/B _4584_/B VGND VGND VPWR VPWR _4581_/B sky130_fd_sc_hd__and3_2
XFILLER_129_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold304 hold304/A VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__dlygate4sd3_1
X_7251_ _7251_/CLK _7251_/D _6472_/A VGND VGND VPWR VPWR _7251_/Q sky130_fd_sc_hd__dfrtp_2
Xhold315 _5672_/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _6774_/Q VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _5060_/B _5044_/A _5260_/A _4738_/B VGND VGND VPWR VPWR _4464_/C sky130_fd_sc_hd__nand4_1
XFILLER_144_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold337 _5634_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _6936_/Q VGND VGND VPWR VPWR hold348/X sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _7049_/Q _6119_/X _6454_/B1 _6953_/Q _6201_/X VGND VGND VPWR VPWR _6205_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold359 _5427_/X VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ input98/X _5331_/C _3540_/B _3413_/X _7079_/Q VGND VGND VPWR VPWR _3414_/X
+ sky130_fd_sc_hd__a32o_2
X_7182_ _7259_/CLK _7182_/D fanout594/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_4
X_4394_ _5042_/A _5055_/D _5042_/B VGND VGND VPWR VPWR _4394_/X sky130_fd_sc_hd__and3_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6132_/Y _6121_/X _6134_/C _6134_/D VGND VGND VPWR VPWR _6339_/D sky130_fd_sc_hd__and4bb_4
X_3345_ _7219_/Q _6848_/Q _6849_/Q VGND VGND VPWR VPWR _3345_/X sky130_fd_sc_hd__mux2_4
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1004 hold1375/X VGND VGND VPWR VPWR _6539_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6686_/Q _5768_/X _5814_/X _6590_/Q _6063_/X VGND VGND VPWR VPWR _6064_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3276_ _6946_/Q VGND VGND VPWR VPWR _3276_/Y sky130_fd_sc_hd__inv_2
Xhold1015 _4205_/X VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _3362_/X VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 _6563_/Q VGND VGND VPWR VPWR _3377_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5015_ _4561_/B _4575_/B _5012_/X _4907_/B VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__a31o_1
Xhold1048 _6568_/Q VGND VGND VPWR VPWR _3384_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1059 _6647_/Q VGND VGND VPWR VPWR _3986_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _7160_/CLK _6966_/D fanout592/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5917_ _6964_/Q _5770_/X _5793_/X _6988_/Q _5916_/X VGND VGND VPWR VPWR _5917_/X
+ sky130_fd_sc_hd__a221o_2
X_6897_ _7073_/CLK _6897_/D fanout585/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_4
X_5848_ _6953_/Q _5776_/X _5793_/X _6985_/Q _5847_/X VGND VGND VPWR VPWR _5848_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5779_ _6010_/D _5783_/C _5795_/D VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__and3_4
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold860 _6605_/Q VGND VGND VPWR VPWR hold860/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold871 _4072_/X VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 _6817_/Q VGND VGND VPWR VPWR hold882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _4058_/X VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6820_ _7265_/CLK _6820_/D fanout575/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6751_ _6751_/CLK _6751_/D _3291_/A VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_4
X_3963_ _3693_/Y _3963_/A1 _3968_/S VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5702_ _5706_/D _5698_/Y _5710_/D _5701_/Y VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__a211oi_1
XFILLER_149_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6682_ _7239_/CLK _6682_/D fanout576/X VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfrtp_2
X_3894_ _6878_/Q _5350_/B _5359_/B _6886_/Q _3893_/X VGND VGND VPWR VPWR _3894_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_176_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5633_ hold2/X _5633_/A1 hold29/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__mux2_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5564_ hold21/X hold190/X _5565_/S VGND VGND VPWR VPWR _5564_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold101 _5581_/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4515_ _4319_/X _4510_/Y _4514_/Y _7259_/Q VGND VGND VPWR VPWR _4516_/A sky130_fd_sc_hd__o31a_1
XFILLER_156_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7303_ _7303_/A VGND VGND VPWR VPWR _7303_/X sky130_fd_sc_hd__clkbuf_1
Xhold112 hold112/A VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _6964_/Q VGND VGND VPWR VPWR hold123/X sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ hold573/X _6543_/A0 _5502_/S VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold134 _6560_/Q VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold145 _3974_/X VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _5569_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7234_ _3340_/A1 _7234_/D fanout613/X VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__dfrtp_2
X_4446_ _4446_/A _4446_/B VGND VGND VPWR VPWR _4446_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold167 _5551_/X VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold178 _6918_/Q VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 input75/X VGND VGND VPWR VPWR fanout603/X sky130_fd_sc_hd__buf_8
Xhold189 _5412_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ _7165_/CLK _7165_/D fanout601/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout614 _4662_/C VGND VGND VPWR VPWR _4657_/C sky130_fd_sc_hd__buf_12
X_4377_ _4984_/B _4984_/C _4859_/C VGND VGND VPWR VPWR _4377_/X sky130_fd_sc_hd__and3_2
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout625 _4255_/A VGND VGND VPWR VPWR _4632_/B sky130_fd_sc_hd__buf_6
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6117_/A _6138_/B _6177_/C VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__and3_4
XFILLER_100_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3328_ _3327_/A _7162_/Q _3327_/Y VGND VGND VPWR VPWR _3328_/Y sky130_fd_sc_hd__o21ai_4
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/CLK _7096_/D fanout596/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfstp_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6047_/A1 _5761_/X _6046_/X _6045_/X VGND VGND VPWR VPWR _7204_/D sky130_fd_sc_hd__o22a_1
X_3259_ _7082_/Q VGND VGND VPWR VPWR _3259_/Y sky130_fd_sc_hd__inv_2
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6949_ _7143_/CLK _6949_/D fanout588/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold690 _6957_/Q VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1390 _5550_/X VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput206 _3249_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
XFILLER_114_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput217 _3341_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
XFILLER_5_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4300_ _4632_/A _4511_/A _4632_/C _4612_/C VGND VGND VPWR VPWR _4308_/D sky130_fd_sc_hd__o211a_2
Xoutput228 _7300_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
XFILLER_154_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput239 _3333_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
X_5280_ _4152_/B _5280_/A1 _5280_/S VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4231_ _4698_/A _4656_/C VGND VGND VPWR VPWR _4320_/A sky130_fd_sc_hd__nand2_8
XFILLER_141_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4162_ _6546_/A0 hold476/X _4162_/S VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4093_ hold980/X _4092_/X _4093_/S VGND VGND VPWR VPWR _4093_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6803_ _7256_/CLK _6803_/D fanout594/X VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4995_ _4640_/A _4719_/B _4683_/X _4987_/C _4872_/C VGND VGND VPWR VPWR _5257_/B
+ sky130_fd_sc_hd__a221oi_2
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6734_ _7239_/CLK _6734_/D fanout574/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfstp_2
X_3946_ _3568_/Y _3946_/A1 _3953_/S VGND VGND VPWR VPWR _6612_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6665_ _6828_/CLK _6665_/D fanout573/X VGND VGND VPWR VPWR _6665_/Q sky130_fd_sc_hd__dfstp_1
X_3877_ _6958_/Q _5485_/B _5440_/C _3536_/X _6990_/Q VGND VGND VPWR VPWR _3877_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5616_ _3924_/B hold246/X _5619_/S VGND VGND VPWR VPWR _5616_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6596_ _7161_/CLK _6596_/D fanout599/X VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_191_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5547_ _5692_/A1 hold927/X hold77/X VGND VGND VPWR VPWR _5547_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5478_ _3915_/B hold342/X _5484_/S VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7217_ _7219_/CLK _7217_/D fanout577/X VGND VGND VPWR VPWR _7217_/Q sky130_fd_sc_hd__dfrtp_1
X_4429_ _4429_/A _5143_/D _4815_/A _4429_/D VGND VGND VPWR VPWR _5044_/B sky130_fd_sc_hd__and4_1
Xfanout422 _6446_/C VGND VGND VPWR VPWR _6425_/B sky130_fd_sc_hd__buf_12
XFILLER_132_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout433 _4474_/X VGND VGND VPWR VPWR _4597_/C sky130_fd_sc_hd__buf_6
X_7148_ _7148_/CLK _7148_/D fanout592/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout455 _3533_/C VGND VGND VPWR VPWR _5422_/D sky130_fd_sc_hd__buf_8
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout466 _5548_/D VGND VGND VPWR VPWR _5675_/D sky130_fd_sc_hd__buf_12
Xfanout477 hold76/X VGND VGND VPWR VPWR _5512_/B sky130_fd_sc_hd__buf_12
Xfanout488 hold66/A VGND VGND VPWR VPWR _6524_/B sky130_fd_sc_hd__buf_12
XFILLER_74_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7079_ _7117_/CLK _7079_/D fanout608/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout499 _5959_/C VGND VGND VPWR VPWR _6028_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_360 _6452_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _5575_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_382 _3969_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_393 _5779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3800_ input48/X _4204_/S _3913_/B _6596_/Q _3799_/X VGND VGND VPWR VPWR _3800_/X
+ sky130_fd_sc_hd__a221o_2
X_4780_ _4692_/Y _4745_/Y _4779_/Y VGND VGND VPWR VPWR _4780_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3731_ _6646_/Q _5485_/B _3457_/X _3730_/X VGND VGND VPWR VPWR _3731_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_0_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7260_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3662_ _6977_/Q _5485_/B _5281_/A2 _3452_/X _6961_/Q VGND VGND VPWR VPWR _3662_/X
+ sky130_fd_sc_hd__a32o_1
X_6450_ _6782_/Q _6130_/X _6144_/X _6652_/Q _6449_/X VGND VGND VPWR VPWR _6450_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5401_ hold180/X hold83/X _5403_/S VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6381_ _6744_/Q _6446_/B _6347_/C _6136_/X _6621_/Q VGND VGND VPWR VPWR _6381_/X
+ sky130_fd_sc_hd__a32o_1
X_3593_ _7000_/Q hold39/A _5273_/D _5593_/B _7088_/Q VGND VGND VPWR VPWR _3593_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5332_ _5649_/A0 _5332_/A1 _5333_/S VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5263_ _5263_/A _5263_/B _5263_/C VGND VGND VPWR VPWR _5263_/X sky130_fd_sc_hd__and3_1
XFILLER_87_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7002_ _7170_/CLK _7002_/D fanout605/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_4
X_4214_ _4214_/A _4214_/B VGND VGND VPWR VPWR _4670_/D sky130_fd_sc_hd__nand2_4
X_5194_ _5194_/A _5194_/B _5194_/C VGND VGND VPWR VPWR _5197_/B sky130_fd_sc_hd__and3_1
X_4145_ _5304_/A _6524_/B _5494_/C _6536_/D VGND VGND VPWR VPWR _4150_/S sky130_fd_sc_hd__and4_2
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ _6851_/Q _6898_/Q _3346_/D _3540_/Y hold66/A VGND VGND VPWR VPWR _4076_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4978_ _4623_/Y _5200_/C _4805_/X _4974_/X _4206_/B VGND VGND VPWR VPWR _4978_/X
+ sky130_fd_sc_hd__o221a_1
X_6717_ _7067_/CLK _6717_/D fanout582/X VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfrtp_1
X_3929_ _6538_/A0 hold433/X _3932_/S VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6648_ _6812_/CLK _6648_/D fanout580/X VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6579_ _7219_/CLK _6579_/D VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5950_ _6949_/Q _5779_/X _5782_/X _6941_/Q _5949_/X VGND VGND VPWR VPWR _5950_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4901_ _4754_/B _4255_/A _5036_/C _4939_/A VGND VGND VPWR VPWR _4901_/X sky130_fd_sc_hd__a31o_1
XFILLER_33_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5881_ _6938_/Q _5782_/X _5876_/X _5878_/X _5880_/X VGND VGND VPWR VPWR _5881_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_61_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4832_ _5261_/D _4832_/B _4832_/C _4832_/D VGND VGND VPWR VPWR _4832_/X sky130_fd_sc_hd__and4_1
XANTENNA_190 _5325_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4763_ _4601_/Y _4638_/Y _4658_/Y _4663_/Y _4743_/Y VGND VGND VPWR VPWR _4763_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_147_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6502_ _6501_/X _3924_/B _6511_/S VGND VGND VPWR VPWR _7233_/D sky130_fd_sc_hd__mux2_1
X_3714_ _6761_/Q _4133_/B _4121_/B _6751_/Q _3713_/X VGND VGND VPWR VPWR _3714_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4694_ _4650_/Y _4692_/Y _4693_/Y _4690_/Y VGND VGND VPWR VPWR _4697_/C sky130_fd_sc_hd__o211ai_1
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6433_ _6577_/Q _6104_/X _6118_/X _6567_/Q _6432_/X VGND VGND VPWR VPWR _6440_/A
+ sky130_fd_sc_hd__a221o_1
X_3645_ _6780_/Q _5311_/B _5422_/D _3528_/X input13/X VGND VGND VPWR VPWR _3645_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6364_ _6597_/Q _6109_/X _6361_/X _6363_/X VGND VGND VPWR VPWR _6365_/D sky130_fd_sc_hd__a211o_1
X_3576_ _6659_/Q _3447_/X _3913_/B _6593_/Q _3575_/X VGND VGND VPWR VPWR _3576_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5315_ _5313_/X _5315_/B _5494_/A hold64/X VGND VGND VPWR VPWR _5315_/X sky130_fd_sc_hd__and4b_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6295_ _7133_/Q _6116_/X _6122_/X _6893_/Q _6294_/X VGND VGND VPWR VPWR _6295_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5246_ _4973_/B _5064_/X _5246_/C _5246_/D VGND VGND VPWR VPWR _5247_/C sky130_fd_sc_hd__and4bb_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _5177_/A _5177_/B _5177_/C _5177_/D VGND VGND VPWR VPWR _5220_/A sky130_fd_sc_hd__nor4_1
XFILLER_69_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4128_ _4152_/B _4128_/A1 _4132_/S VGND VGND VPWR VPWR _4128_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4059_ _3915_/X hold613/X _4065_/S VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6855_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire450 _5313_/D VGND VGND VPWR VPWR _3528_/C sky130_fd_sc_hd__buf_2
XFILLER_156_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold508 _6756_/Q VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3430_ _5304_/A _5666_/C _5575_/C VGND VGND VPWR VPWR _3969_/C sky130_fd_sc_hd__and3_4
Xhold519 hold519/A VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3361_ input58/X hold211/X hold65/X VGND VGND VPWR VPWR _3361_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_95_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7241_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5100_/A _5100_/B _5100_/C VGND VGND VPWR VPWR _5220_/C sky130_fd_sc_hd__and3_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _7248_/Q _5723_/X wire398/X _7269_/Q _6079_/X VGND VGND VPWR VPWR _6080_/X
+ sky130_fd_sc_hd__a221o_1
X_3292_ _7311_/A VGND VGND VPWR VPWR _3292_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _4595_/A _4774_/B _4596_/B _5030_/X VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__a211oi_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _4178_/X VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 _6975_/Q VGND VGND VPWR VPWR _5468_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6982_ _7157_/CLK _6982_/D fanout592/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfrtp_4
X_5933_ _7005_/Q _5934_/C _5782_/C _5795_/C VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7122_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5864_ _7122_/Q _5826_/B _5911_/C _5779_/X _6946_/Q VGND VGND VPWR VPWR _5869_/B
+ sky130_fd_sc_hd__a32o_1
X_4815_ _4815_/A _5260_/B VGND VGND VPWR VPWR _4815_/Y sky130_fd_sc_hd__nand2_1
X_5795_ _7181_/Q _7180_/Q _5795_/C _5795_/D VGND VGND VPWR VPWR _5795_/X sky130_fd_sc_hd__and4_4
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_48_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7006_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4746_ _4746_/A _4939_/B _4923_/C VGND VGND VPWR VPWR _4746_/X sky130_fd_sc_hd__and3_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4677_ _4748_/B _4945_/C _4755_/B VGND VGND VPWR VPWR _4678_/B sky130_fd_sc_hd__and3_1
X_6416_ _6690_/Q _6466_/A1 _5759_/A VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__o21a_1
X_3628_ _7276_/Q _5630_/A _3466_/X _3499_/X _7016_/Q VGND VGND VPWR VPWR _3628_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6347_ _6743_/Q _6446_/B _6347_/C VGND VGND VPWR VPWR _6347_/X sky130_fd_sc_hd__and3_1
XFILLER_143_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3559_ _5449_/B _5476_/C _5422_/D VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__and3_4
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6278_ _6916_/Q _6451_/B1 _6122_/X _6892_/Q _6277_/X VGND VGND VPWR VPWR _6278_/X
+ sky130_fd_sc_hd__a221o_1
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4227_/B sky130_fd_sc_hd__clkbuf_2
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _3312_/D sky130_fd_sc_hd__clkbuf_1
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4662_/C sky130_fd_sc_hd__clkbuf_2
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6487_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5229_ _5255_/B _5128_/B _4987_/A _4987_/B _4862_/A VGND VGND VPWR VPWR _5231_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_56_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _5788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4600_ _4632_/B _4600_/B _4612_/C _4549_/D VGND VGND VPWR VPWR _4600_/Y sky130_fd_sc_hd__nor4b_2
X_5580_ _5580_/A0 hold5/X hold18/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4531_ _4815_/A _4589_/B _4561_/B VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__and3_1
Xhold305 _6886_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _6961_/Q VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_7250_ _7259_/CLK _7250_/D _6472_/A VGND VGND VPWR VPWR _7250_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4462_ _4409_/C _4654_/B _4391_/Y _4870_/C _4358_/X VGND VGND VPWR VPWR _4464_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_171_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold327 _4154_/X VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _7012_/Q VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold349 _5424_/X VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _7137_/Q _6145_/C _6114_/X _6129_/C _7153_/Q VGND VGND VPWR VPWR _6201_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3413_ _6548_/A _5675_/D _5657_/D VGND VGND VPWR VPWR _3413_/X sky130_fd_sc_hd__and3_4
X_7181_ _7256_/CLK _7181_/D fanout594/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfstp_4
X_4393_ _5143_/A _5260_/B _5128_/B _5143_/D VGND VGND VPWR VPWR _4459_/B sky130_fd_sc_hd__nand4_1
X_3344_ _7206_/Q _6847_/Q _6849_/Q VGND VGND VPWR VPWR _3344_/X sky130_fd_sc_hd__mux2_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _6127_/X _6132_/B _6132_/C VGND VGND VPWR VPWR _6132_/Y sky130_fd_sc_hd__nand3b_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6761_/Q _5771_/X _5795_/X _6676_/Q VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__a22o_1
X_3275_ _6954_/Q VGND VGND VPWR VPWR _3275_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _6927_/Q VGND VGND VPWR VPWR _5414_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 hold1368/X VGND VGND VPWR VPWR _3957_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _6755_/Q VGND VGND VPWR VPWR _4130_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1038 _3377_/X VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5014_ _5263_/A _4606_/D _4589_/C _5012_/X _4898_/X VGND VGND VPWR VPWR _5264_/C
+ sky130_fd_sc_hd__a41oi_2
Xhold1049 _3384_/X VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7015_/CLK _6965_/D fanout588/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5916_ _6980_/Q _6073_/B2 _5774_/X _6908_/Q _5915_/X VGND VGND VPWR VPWR _5916_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6896_ _7148_/CLK _6896_/D fanout591/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _7041_/Q _6059_/S _6028_/B _5815_/X _7017_/Q VGND VGND VPWR VPWR _5847_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5778_ _7181_/Q _7183_/Q _7182_/Q _7180_/Q VGND VGND VPWR VPWR _5959_/B sky130_fd_sc_hd__and4bb_4
XFILLER_154_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4729_ _4729_/A _5128_/A _4860_/C _4729_/D VGND VGND VPWR VPWR _4729_/X sky130_fd_sc_hd__and4_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold850 _7058_/Q VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _3937_/X VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold872 _7244_/Q VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _5281_/X VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold894 hold894/A VGND VGND VPWR VPWR hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1550 _7207_/Q VGND VGND VPWR VPWR _6192_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6750_ _6781_/CLK _6750_/D _3291_/A VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3962_ _3632_/Y _3962_/A1 _3968_/S VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__mux2_1
X_5701_ _7176_/Q _5706_/D VGND VGND VPWR VPWR _5701_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6681_ _7265_/CLK _6681_/D fanout575/X VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3893_ _7046_/Q _5512_/B _5684_/C _3428_/X _7014_/Q VGND VGND VPWR VPWR _3893_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5632_ _5632_/A0 _3915_/X _5637_/S VGND VGND VPWR VPWR _5632_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5563_ _4049_/B hold251/X _5565_/S VGND VGND VPWR VPWR _5563_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7302_ _7302_/A VGND VGND VPWR VPWR _7302_/X sky130_fd_sc_hd__clkbuf_1
X_4514_ _4970_/D _4755_/D VGND VGND VPWR VPWR _4514_/Y sky130_fd_sc_hd__nand2_4
Xhold102 _6868_/Q VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _5494_/A hold39/X _5494_/C VGND VGND VPWR VPWR _5502_/S sky130_fd_sc_hd__and3_4
Xhold113 _7004_/Q VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _5455_/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _3374_/X VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7233_ _7254_/CLK _7233_/D fanout613/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfrtp_1
XFILLER_132_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold146 _6914_/Q VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4859_/C _4460_/B _5140_/B VGND VGND VPWR VPWR _4446_/A sky130_fd_sc_hd__and3_1
XFILLER_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold157 _7236_/Q VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _6924_/Q VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold179 _5403_/X VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7164_ _7174_/CLK _7164_/D fanout608/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout604 fanout607/X VGND VGND VPWR VPWR fanout604/X sky130_fd_sc_hd__buf_8
Xfanout615 _4999_/A1 VGND VGND VPWR VPWR _4698_/A sky130_fd_sc_hd__buf_12
X_4376_ _4285_/A _4346_/A _4667_/D _4859_/A VGND VGND VPWR VPWR _4376_/Y sky130_fd_sc_hd__o211ai_4
Xfanout626 input110/X VGND VGND VPWR VPWR _4255_/A sky130_fd_sc_hd__buf_8
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6115_ _6117_/A _6444_/C _6177_/C VGND VGND VPWR VPWR _6115_/X sky130_fd_sc_hd__and3_4
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3327_ _3327_/A _3327_/B VGND VGND VPWR VPWR _3327_/Y sky130_fd_sc_hd__nand2_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7159_/CLK _7095_/D fanout599/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_113_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6046_ _6442_/S _7203_/Q _6443_/S VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3258_ _7090_/Q VGND VGND VPWR VPWR _3258_/Y sky130_fd_sc_hd__inv_2
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _7154_/CLK _6948_/D fanout592/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6879_ _7151_/CLK _6879_/D fanout585/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_167_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold680 _6965_/Q VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _5447_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1380 _6813_/Q VGND VGND VPWR VPWR hold1380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1391 _6888_/Q VGND VGND VPWR VPWR hold380/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput207 _3281_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
Xoutput218 _7291_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
Xoutput229 _7301_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ _4230_/A _4230_/B VGND VGND VPWR VPWR _4310_/B sky130_fd_sc_hd__nor2_8
XFILLER_99_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4161_ _5311_/B _4158_/D _3919_/X _4162_/S hold936/X VGND VGND VPWR VPWR _4161_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ hold128/X _4053_/X _4092_/S VGND VGND VPWR VPWR _4092_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6802_ _7256_/CLK _6802_/D fanout594/X VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4994_ _4408_/X _4722_/Y _4867_/C _4681_/C _4992_/X VGND VGND VPWR VPWR _4997_/A
+ sky130_fd_sc_hd__o2111a_1
X_6733_ _6827_/CLK _6733_/D fanout574/X VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfstp_2
X_3945_ _3945_/A _6472_/A VGND VGND VPWR VPWR _3953_/S sky130_fd_sc_hd__nand2_4
X_6664_ _6976_/CLK _6664_/D fanout590/X VGND VGND VPWR VPWR _6664_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3876_ _3875_/Y _3876_/A1 _3906_/S VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5615_ _3921_/B hold324/X _5619_/S VGND VGND VPWR VPWR _5615_/X sky130_fd_sc_hd__mux2_1
X_6595_ _7111_/CLK _6595_/D fanout599/X VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5546_ hold21/X _5546_/A1 hold77/X VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__mux2_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5477_ _5667_/A0 _5477_/A1 _5484_/S VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7216_ _7219_/CLK _7216_/D fanout577/X VGND VGND VPWR VPWR _7216_/Q sky130_fd_sc_hd__dfrtp_1
X_4428_ _4271_/Y _4423_/Y _4427_/Y VGND VGND VPWR VPWR _4428_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout412 _3386_/X VGND VGND VPWR VPWR _5341_/A sky130_fd_sc_hd__buf_12
XFILLER_120_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout423 _5747_/X VGND VGND VPWR VPWR _6446_/C sky130_fd_sc_hd__buf_8
XFILLER_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7147_ _7157_/CLK _7147_/D fanout593/X VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout434 _4519_/C VGND VGND VPWR VPWR _5128_/B sky130_fd_sc_hd__buf_6
Xfanout445 wire447/X VGND VGND VPWR VPWR _5311_/C sky130_fd_sc_hd__buf_12
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4359_ _4722_/A _4984_/A VGND VGND VPWR VPWR _4359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout456 hold1499/X VGND VGND VPWR VPWR _3533_/C sky130_fd_sc_hd__buf_8
Xfanout467 _3404_/X VGND VGND VPWR VPWR _5548_/D sky130_fd_sc_hd__buf_12
XFILLER_100_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout478 hold76/X VGND VGND VPWR VPWR _5548_/C sky130_fd_sc_hd__buf_6
Xfanout489 hold66/A VGND VGND VPWR VPWR _6548_/B sky130_fd_sc_hd__buf_12
X_7078_ _7173_/CLK _7078_/D fanout603/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6029_ _6609_/Q _6025_/B _6003_/C _6028_/X VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__a31o_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _6805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_361 _6129_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_372 _5657_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_383 _3969_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_394 _5815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _6590_/Q _5512_/B _3446_/X _5639_/B hold52/A VGND VGND VPWR VPWR _3730_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_159_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3661_ _6852_/Q _5311_/B _5327_/D _4133_/B _6760_/Q VGND VGND VPWR VPWR _3661_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_158_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5400_ hold500/X _3925_/C _5403_/S VGND VGND VPWR VPWR _5400_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6380_ _6380_/A _6380_/B _6380_/C _6380_/D VGND VGND VPWR VPWR _6390_/C sky130_fd_sc_hd__nor4_1
X_3592_ _6634_/Q _3969_/C _3587_/X _3590_/X _3591_/X VGND VGND VPWR VPWR _3592_/Y
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5331_ _6536_/B _6530_/D _5331_/C _5575_/D VGND VGND VPWR VPWR _5333_/S sky130_fd_sc_hd__nand4_2
XFILLER_141_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5262_ _5184_/C _5262_/B _5262_/C VGND VGND VPWR VPWR _5262_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_141_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7001_ _7067_/CLK _7001_/D fanout582/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4213_ _4637_/A _4747_/A _4747_/B _4747_/C VGND VGND VPWR VPWR _4214_/B sky130_fd_sc_hd__nand4_4
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5193_ _4862_/A _4791_/B _4778_/C _4879_/B _5192_/X VGND VGND VPWR VPWR _5194_/C
+ sky130_fd_sc_hd__a311oi_1
X_4144_ hold996/X _6535_/A0 _4144_/S VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4075_ _6511_/A1 hold272/X hold57/X VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7277_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4977_ _4290_/Y _4423_/Y _4501_/Y _4740_/Y VGND VGND VPWR VPWR _5200_/C sky130_fd_sc_hd__o31a_1
X_6716_ _7132_/CLK _6716_/D fanout610/X VGND VGND VPWR VPWR _7306_/A sky130_fd_sc_hd__dfrtp_1
X_3928_ _3370_/B hold986/X _3932_/S VGND VGND VPWR VPWR _3928_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6647_ _6676_/CLK _6647_/D fanout579/X VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3859_ _3345_/X _5331_/C _4139_/C _3433_/X _6941_/Q VGND VGND VPWR VPWR _3859_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6578_ _7017_/CLK _6578_/D fanout604/X VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_124_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5529_ hold905/X _5692_/A1 _5529_/S VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap409 _5629_/C VGND VGND VPWR VPWR _3902_/A3 sky130_fd_sc_hd__buf_12
XFILLER_40_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4900_ _4540_/Y _4541_/Y _4774_/B _4620_/B VGND VGND VPWR VPWR _4900_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5880_ _6978_/Q _6073_/B2 _5780_/X _7098_/Q _5879_/X VGND VGND VPWR VPWR _5880_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4831_ _4738_/B _4597_/C _5060_/C _5143_/A _5260_/B VGND VGND VPWR VPWR _4832_/D
+ sky130_fd_sc_hd__o2111ai_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_180 _6734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_191 _3902_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4762_ _4777_/C _4761_/X _4750_/B VGND VGND VPWR VPWR _4765_/B sky130_fd_sc_hd__o21ai_1
X_6501_ _7257_/Q _6501_/A2 _6501_/B1 _4164_/Y _6500_/X VGND VGND VPWR VPWR _6501_/X
+ sky130_fd_sc_hd__a221o_1
X_3713_ _6814_/Q _5341_/A _5485_/B _3538_/X _7042_/Q VGND VGND VPWR VPWR _3713_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4693_ _4708_/A _4778_/C VGND VGND VPWR VPWR _4693_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6432_ _7278_/Q _6444_/C _5750_/C _6137_/X _7273_/Q VGND VGND VPWR VPWR _6432_/X
+ sky130_fd_sc_hd__a32o_1
X_3644_ input26/X _3504_/X _3553_/X _6680_/Q _3643_/X VGND VGND VPWR VPWR _3644_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6363_ _6602_/Q _6105_/X _6106_/X _7265_/Q _6362_/X VGND VGND VPWR VPWR _6363_/X
+ sky130_fd_sc_hd__a221o_1
X_3575_ _6779_/Q _5311_/B _3533_/C _4092_/S input47/X VGND VGND VPWR VPWR _3575_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5314_ _5476_/B _5476_/C _5311_/C _5314_/B1 VGND VGND VPWR VPWR _5315_/B sky130_fd_sc_hd__a31o_1
XFILLER_161_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6294_ _7077_/Q _6446_/C _6425_/C _6109_/X _7045_/Q VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5245_ _4480_/B _4799_/C _4843_/A _5085_/X _5244_/X VGND VGND VPWR VPWR _5246_/D
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__buf_6
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__buf_6
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5176_ _4923_/A _5263_/B _4923_/C _4587_/A VGND VGND VPWR VPWR _5177_/D sky130_fd_sc_hd__a31o_1
XFILLER_56_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4127_ _6536_/B _6536_/C _4127_/C _5273_/D VGND VGND VPWR VPWR _4132_/S sky130_fd_sc_hd__nand4_4
XFILLER_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4058_ _4065_/S hold892/X _3370_/X _4055_/X VGND VGND VPWR VPWR _4058_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire440 _4263_/Y VGND VGND VPWR VPWR _5143_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_143_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold509 _4131_/X VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3360_ hold13/A hold65/X VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__and2_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3291_/A VGND VGND VPWR VPWR _7309_/A sky130_fd_sc_hd__inv_2
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _4595_/A _4597_/C _4923_/A _4923_/B _4603_/B VGND VGND VPWR VPWR _5030_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1209 hold1483/X VGND VGND VPWR VPWR _5432_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6981_ _7015_/CLK _6981_/D fanout591/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5932_ _5954_/A2 _5761_/X _5931_/X VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5863_ _7002_/Q _5795_/D _6010_/C _5815_/B VGND VGND VPWR VPWR _5869_/A sky130_fd_sc_hd__o211a_1
XFILLER_34_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4814_ _5060_/B _4815_/A _4449_/A _4461_/A VGND VGND VPWR VPWR _4814_/Y sky130_fd_sc_hd__a31oi_2
X_5794_ _5815_/C _5814_/C _5934_/C VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__and3_4
X_4745_ _4761_/A _4939_/B VGND VGND VPWR VPWR _4745_/Y sky130_fd_sc_hd__nand2_4
XFILLER_119_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4676_ _5036_/C _4633_/B _4674_/D _4940_/C _4722_/A VGND VGND VPWR VPWR _4676_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6415_ _6396_/X _6415_/B _6415_/C VGND VGND VPWR VPWR _6415_/Y sky130_fd_sc_hd__nand3b_2
X_3627_ _6570_/Q _6548_/A _5341_/A _3525_/X _7120_/Q VGND VGND VPWR VPWR _3627_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6346_ _7275_/Q _6112_/X _6118_/X _6564_/Q _6345_/X VGND VGND VPWR VPWR _6356_/A
+ sky130_fd_sc_hd__a221o_1
X_3558_ _3987_/A _6530_/C _6548_/D VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__and3_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6277_ _7076_/Q _6425_/B _6425_/C _6452_/B1 _6980_/Q VGND VGND VPWR VPWR _6277_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3489_ _5476_/B _5422_/D _5575_/D VGND VGND VPWR VPWR _3489_/X sky130_fd_sc_hd__and3_1
XFILLER_88_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4227_/A sky130_fd_sc_hd__clkbuf_2
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__clkbuf_1
X_5228_ _5228_/A _5228_/B _5228_/C VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__and3_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4229_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5159_ _5159_/A _5270_/B _5159_/C VGND VGND VPWR VPWR _5164_/A sky130_fd_sc_hd__and3_1
XFILLER_57_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_80 _5776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _5793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4530_ _4597_/C _4586_/B _5263_/A _4561_/B VGND VGND VPWR VPWR _4565_/D sky130_fd_sc_hd__nand4_1
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4461_ _4461_/A _4461_/B _4461_/C VGND VGND VPWR VPWR _4464_/A sky130_fd_sc_hd__nor3_1
Xhold306 _5367_/X VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_100_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7268_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold317 _5452_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _7272_/Q VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _6881_/Q _6101_/X _6143_/X _6945_/Q _6199_/X VGND VGND VPWR VPWR _6205_/B
+ sky130_fd_sc_hd__a221o_1
Xhold339 _5509_/X VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ hold26/X hold71/X _5657_/D hold65/A VGND VGND VPWR VPWR _3412_/X sky130_fd_sc_hd__and4b_4
X_7180_ _7251_/CLK _7180_/D fanout594/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4392_ _5260_/B _5128_/B VGND VGND VPWR VPWR _4392_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6145_/C _6114_/X _6116_/X _6130_/X _6101_/X VGND VGND VPWR VPWR _6132_/C
+ sky130_fd_sc_hd__a2111oi_1
X_3343_ _7193_/Q _6845_/Q _6849_/Q VGND VGND VPWR VPWR _3343_/X sky130_fd_sc_hd__mux2_2
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6814_/Q _6028_/C _5782_/C _5795_/C VGND VGND VPWR VPWR _6062_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _6962_/Q VGND VGND VPWR VPWR _3274_/Y sky130_fd_sc_hd__inv_2
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _5414_/X VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 _6881_/Q VGND VGND VPWR VPWR _5362_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _4589_/B _4589_/C _5012_/X _4897_/X VGND VGND VPWR VPWR _5100_/B sky130_fd_sc_hd__a31oi_1
Xhold1028 _4130_/X VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1039 _7262_/Q VGND VGND VPWR VPWR _6533_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6964_ _7151_/CLK _6964_/D fanout586/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5915_ _6884_/Q _5768_/X _5794_/X _6924_/Q _5913_/X VGND VGND VPWR VPWR _5915_/X
+ sky130_fd_sc_hd__a221o_1
X_6895_ _7073_/CLK _6895_/D fanout585/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5846_ _6977_/Q _6073_/B2 _5970_/B1 _6929_/Q VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5777_ _6059_/S _6010_/D _5783_/C VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__and3_4
X_4728_ _5128_/A _4740_/C _4738_/B _4987_/B VGND VGND VPWR VPWR _5009_/B sky130_fd_sc_hd__nand4_1
XFILLER_175_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4659_ _4708_/A _4659_/B VGND VGND VPWR VPWR _4659_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold840 _5411_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold851 _5561_/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 _7110_/Q VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _6525_/X VGND VGND VPWR VPWR _7244_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold884 _6659_/Q VGND VGND VPWR VPWR hold884/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6329_ _7110_/Q _6112_/X _6119_/X _7054_/Q _6328_/X VGND VGND VPWR VPWR _6330_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold895 _6923_/Q VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1540 _7219_/Q VGND VGND VPWR VPWR _6468_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1551 _6804_/Q VGND VGND VPWR VPWR _4206_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_94_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6780_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7123_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7053_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ _3568_/Y _3961_/A1 _3968_/S VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5700_ _6803_/Q _6292_/S _5759_/B _7176_/Q _3307_/Y VGND VGND VPWR VPWR _5710_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_188_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6680_ _6828_/CLK _6680_/D fanout574/X VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3892_ _3352_/B _4092_/S _3452_/X _6966_/Q _3891_/X VGND VGND VPWR VPWR _3892_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_176_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5631_ _6543_/A0 hold888/X hold29/X VGND VGND VPWR VPWR _5631_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5562_ _3924_/B hold552/X _5565_/S VGND VGND VPWR VPWR _5562_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7301_ _7301_/A VGND VGND VPWR VPWR _7301_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4513_ _4255_/A _4600_/B _4612_/C _4549_/D VGND VGND VPWR VPWR _4730_/D sky130_fd_sc_hd__and4b_4
XFILLER_144_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold103 _5347_/X VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ hold262/X _6511_/A1 _5493_/S VGND VGND VPWR VPWR _5493_/X sky130_fd_sc_hd__mux2_1
Xhold114 _5500_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7232_ _7254_/CLK _7232_/D fanout613/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfrtp_2
Xhold125 hold157/X VGND VGND VPWR VPWR hold158/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _6699_/Q VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4444_ _4444_/A _4444_/B _4444_/C VGND VGND VPWR VPWR _4446_/B sky130_fd_sc_hd__nand3_1
Xhold147 _5399_/X VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold158 hold158/A VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _5410_/X VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _7163_/CLK _7163_/D fanout608/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4375_ _4859_/A _4667_/C _4667_/D VGND VGND VPWR VPWR _4375_/X sky130_fd_sc_hd__and3_2
Xfanout605 fanout607/X VGND VGND VPWR VPWR fanout605/X sky130_fd_sc_hd__buf_4
Xfanout616 _4848_/A VGND VGND VPWR VPWR _4656_/C sky130_fd_sc_hd__buf_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _7186_/Q _7189_/Q _7190_/Q _7185_/Q VGND VGND VPWR VPWR _6114_/X sky130_fd_sc_hd__and4bb_4
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3327_/A _7170_/Q _3325_/Y VGND VGND VPWR VPWR _3326_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7094_ _7156_/CLK _7094_/D fanout603/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6690_/Q _5726_/Y _6032_/X _6044_/X _5759_/A VGND VGND VPWR VPWR _6045_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _7098_/Q VGND VGND VPWR VPWR _3257_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6947_ _7152_/CLK _6947_/D fanout586/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6878_ _7108_/CLK _6878_/D fanout606/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5829_ _6992_/Q _5959_/C _5911_/C _5825_/X _5828_/X VGND VGND VPWR VPWR _5829_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_155_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold670 _5393_/X VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 _5456_/X VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _6588_/Q VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1370 _6737_/Q VGND VGND VPWR VPWR hold940/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1381 _5276_/X VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1392 _5370_/X VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput208 _3280_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput219 _7292_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ _6538_/A0 hold399/X _4162_/S VGND VGND VPWR VPWR _4160_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4091_ _4091_/A0 _4090_/X _4093_/S VGND VGND VPWR VPWR _4091_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6801_ _7256_/CLK _6801_/D fanout577/X VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4993_ _4643_/Y _4650_/Y _4722_/Y _4254_/Y _4867_/C VGND VGND VPWR VPWR _5257_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6732_ _6889_/CLK _6732_/D fanout582/X VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfstp_2
X_3944_ _6535_/A0 _3944_/A1 _3944_/S VGND VGND VPWR VPWR _3944_/X sky130_fd_sc_hd__mux2_1
X_6663_ _6828_/CLK _6663_/D fanout573/X VGND VGND VPWR VPWR _6663_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3875_ _3875_/A _3875_/B VGND VGND VPWR VPWR _3875_/Y sky130_fd_sc_hd__nand2_4
XFILLER_149_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5614_ _3918_/B hold627/X _5619_/S VGND VGND VPWR VPWR _5614_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6594_ _7114_/CLK _6594_/D fanout604/X VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5545_ _6505_/A1 hold856/X hold77/X VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5476_ _5494_/A _5476_/B _5476_/C _5494_/C VGND VGND VPWR VPWR _5476_/Y sky130_fd_sc_hd__nand4_1
Xclkbuf_3_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_144_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7215_ _7218_/CLK _7215_/D fanout594/X VGND VGND VPWR VPWR _7215_/Q sky130_fd_sc_hd__dfrtp_1
X_4427_ _4427_/A _4427_/B _4427_/C _4427_/D VGND VGND VPWR VPWR _4427_/Y sky130_fd_sc_hd__nand4_1
Xfanout413 _3368_/X VGND VGND VPWR VPWR _5311_/B sky130_fd_sc_hd__buf_12
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7146_ _7156_/CLK _7146_/D fanout602/X VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout424 _6117_/C VGND VGND VPWR VPWR _6444_/C sky130_fd_sc_hd__buf_12
X_4358_ _4243_/A _4243_/B _4346_/Y _4356_/Y VGND VGND VPWR VPWR _4358_/X sky130_fd_sc_hd__a211o_4
XFILLER_98_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout457 _5657_/D VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__buf_8
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout468 hold56/X VGND VGND VPWR VPWR _5666_/C sky130_fd_sc_hd__buf_12
X_3309_ _6292_/S _3307_/B _3308_/X VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__a21o_1
X_7077_ _7077_/CLK _7077_/D fanout587/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout479 _6548_/C VGND VGND VPWR VPWR _6536_/C sky130_fd_sc_hd__buf_12
X_4289_ _4637_/A _4747_/B _4747_/C _4984_/B VGND VGND VPWR VPWR _4730_/C sky130_fd_sc_hd__nor4_1
XFILLER_58_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6028_ _6665_/Q _6028_/B _6028_/C VGND VGND VPWR VPWR _6028_/X sky130_fd_sc_hd__and3_1
XFILLER_74_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_340 _7160_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 _5970_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_373 _4127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 _3969_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 _6098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ _6937_/Q _3433_/X _3657_/X _3658_/X _3659_/X VGND VGND VPWR VPWR _3692_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_186_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3591_ _6912_/Q _4158_/D _5281_/A2 _3513_/X _6669_/Q VGND VGND VPWR VPWR _3591_/X
+ sky130_fd_sc_hd__a32o_1
X_5330_ _6549_/A0 _5330_/A1 _5330_/S VGND VGND VPWR VPWR _5330_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5261_ _5260_/X _5259_/X _5261_/C _5261_/D VGND VGND VPWR VPWR _5262_/C sky130_fd_sc_hd__and4bb_1
XFILLER_141_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7000_ _7151_/CLK _7000_/D fanout586/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_142_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4212_ _4689_/B _4511_/A _4632_/C _4612_/C VGND VGND VPWR VPWR _5040_/C sky130_fd_sc_hd__nand4_4
X_5192_ _4862_/A _4738_/B _4878_/B _4878_/C _4697_/B VGND VGND VPWR VPWR _5192_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4143_ hold540/X _6546_/A0 _4144_/S VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4074_ hold8/X _3539_/X _4051_/X hold57/X hold510/X VGND VGND VPWR VPWR _4074_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4976_ _4976_/A _4976_/B _4976_/C _4976_/D VGND VGND VPWR VPWR _4976_/Y sky130_fd_sc_hd__nor4_1
X_6715_ _7163_/CLK _6715_/D fanout610/X VGND VGND VPWR VPWR _7305_/A sky130_fd_sc_hd__dfrtp_1
X_3927_ _6542_/A _3927_/B VGND VGND VPWR VPWR _3932_/S sky130_fd_sc_hd__nand2_4
XFILLER_177_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3858_ input27/X _3471_/X _3488_/X _7077_/Q _3857_/X VGND VGND VPWR VPWR _3874_/A
+ sky130_fd_sc_hd__a221o_1
X_6646_ _7263_/CLK _6646_/D fanout577/X VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3789_ _7083_/Q _6548_/A _3412_/X _3907_/B _6591_/Q VGND VGND VPWR VPWR _3789_/X
+ sky130_fd_sc_hd__a32o_1
X_6577_ _7099_/CLK _6577_/D fanout604/X VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_133_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5528_ hold151/X hold21/X _5529_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5459_ _5649_/A0 _5459_/A1 _5466_/S VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7129_ _7129_/CLK _7129_/D fanout598/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4830_ _4380_/X _4403_/X _5040_/A _4820_/X _4829_/X VGND VGND VPWR VPWR _4832_/C
+ sky130_fd_sc_hd__o311a_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _7317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_181 _6466_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_192 _5311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _4761_/A _4939_/B _4761_/C VGND VGND VPWR VPWR _4761_/X sky130_fd_sc_hd__and3_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6500_ _7259_/Q _6500_/A2 _6500_/B1 _7258_/Q VGND VGND VPWR VPWR _6500_/X sky130_fd_sc_hd__a22o_1
X_3712_ input95/X _5331_/C _3540_/B _3536_/X _6986_/Q VGND VGND VPWR VPWR _3712_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4692_ _4777_/A _4777_/B VGND VGND VPWR VPWR _4692_/Y sky130_fd_sc_hd__nand2_2
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3643_ _6921_/Q _3540_/B _5422_/D _3471_/X input22/X VGND VGND VPWR VPWR _3643_/X
+ sky130_fd_sc_hd__a32o_1
X_6431_ _6431_/A _6431_/B _6431_/C _6431_/D VGND VGND VPWR VPWR _6431_/Y sky130_fd_sc_hd__nor4_1
XFILLER_162_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6362_ _6607_/Q _6465_/A2 _6465_/A3 _6110_/X _6554_/Q VGND VGND VPWR VPWR _6362_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3574_ _6742_/Q _5327_/D _5575_/C _5575_/D VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__and4_1
XFILLER_127_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5313_ hold211/X _5476_/B _5548_/D _5313_/D VGND VGND VPWR VPWR _5313_/X sky130_fd_sc_hd__and4b_1
X_6293_ _6292_/X _6293_/A1 _6343_/S VGND VGND VPWR VPWR _7212_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5244_ _4689_/C _4792_/A _4788_/A _4970_/B _4984_/A VGND VGND VPWR VPWR _5244_/X
+ sky130_fd_sc_hd__a32o_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__buf_8
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _5094_/A _5175_/B _5175_/C VGND VGND VPWR VPWR _5266_/A sky130_fd_sc_hd__and3b_1
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4126_ _6535_/A0 _4126_/A1 _4126_/S VGND VGND VPWR VPWR _4126_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4057_ _4204_/S _5341_/C VGND VGND VPWR VPWR _4065_/S sky130_fd_sc_hd__nand2_8
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4959_ _4601_/Y _4629_/Y _5248_/A3 _4692_/Y _4939_/Y VGND VGND VPWR VPWR _4959_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_184_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6629_ _7237_/CLK _6629_/D VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3290_ _4647_/C VGND VGND VPWR VPWR _4761_/C sky130_fd_sc_hd__clkinv_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6980_ _7150_/CLK _6980_/D fanout602/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5931_ _6292_/S _7198_/Q _6443_/S _5930_/X VGND VGND VPWR VPWR _5931_/X sky130_fd_sc_hd__a211o_1
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5862_ _5862_/A1 _5761_/X _5861_/X VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4813_ _5060_/B _4815_/A _5060_/C _5143_/A _4465_/A VGND VGND VPWR VPWR _4813_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_61_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5793_ _7183_/Q _7182_/Q _5815_/C _5795_/D VGND VGND VPWR VPWR _5793_/X sky130_fd_sc_hd__and4_4
XFILLER_178_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4744_ _4761_/A _4760_/B _4760_/C VGND VGND VPWR VPWR _4774_/B sky130_fd_sc_hd__and3_2
XFILLER_193_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4675_ _4675_/A _4675_/B VGND VGND VPWR VPWR _4675_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6414_ _6414_/A _6414_/B _6414_/C _6440_/D VGND VGND VPWR VPWR _6415_/C sky130_fd_sc_hd__nor4_1
X_3626_ _6769_/Q _3482_/X _3621_/X _3622_/X _3625_/X VGND VGND VPWR VPWR _3626_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_135_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3557_ _6678_/Q _5304_/A _6536_/D _4158_/D _3556_/X VGND VGND VPWR VPWR _3557_/X
+ sky130_fd_sc_hd__a41o_1
X_6345_ _6574_/Q _6104_/X _6122_/X _6678_/Q _6344_/X VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6276_ _6932_/Q _6130_/X _6144_/X _7084_/Q _6275_/X VGND VGND VPWR VPWR _6276_/X
+ sky130_fd_sc_hd__a221o_1
X_3488_ hold17/A _5575_/C _5575_/D VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__and3_4
XFILLER_130_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4227_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_88_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5227_ _4939_/A _4738_/B _4729_/D _4859_/A _4984_/C VGND VGND VPWR VPWR _5228_/C
+ sky130_fd_sc_hd__o2111ai_1
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5158_ _5248_/A3 _5153_/X _4692_/Y _4959_/X _5076_/B VGND VGND VPWR VPWR _5159_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4109_ hold83/X hold93/X _4111_/S VGND VGND VPWR VPWR _4109_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5089_ _5089_/A _5089_/B _5089_/C VGND VGND VPWR VPWR _5089_/X sky130_fd_sc_hd__and3_1
XFILLER_16_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_70 _5574_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _5779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_92 _5793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4460_ _4859_/C _4460_/B _4460_/C VGND VGND VPWR VPWR _4461_/B sky130_fd_sc_hd__and3_1
Xhold307 _6953_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold318 _6977_/Q VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _6545_/X VGND VGND VPWR VPWR _7272_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ hold37/X hold42/X _5324_/B VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__o21ai_2
X_4391_ _4860_/B _4632_/C _4511_/A _4632_/A VGND VGND VPWR VPWR _4391_/Y sky130_fd_sc_hd__nand4_4
XFILLER_171_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6130_ _6130_/A _6136_/A _6143_/C VGND VGND VPWR VPWR _6130_/X sky130_fd_sc_hd__and3_4
X_3342_ _7191_/Q _6846_/Q _6849_/Q VGND VGND VPWR VPWR _3342_/X sky130_fd_sc_hd__mux2_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _7268_/Q _6072_/B wire398/X _5763_/X _6756_/Q VGND VGND VPWR VPWR _6061_/X
+ sky130_fd_sc_hd__a32o_1
X_3273_ _6970_/Q VGND VGND VPWR VPWR _3273_/Y sky130_fd_sc_hd__inv_2
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1007 _6601_/Q VGND VGND VPWR VPWR _3932_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5012_ _4689_/B _4255_/A _4633_/B _4786_/B VGND VGND VPWR VPWR _5012_/X sky130_fd_sc_hd__a31o_2
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _5362_/X VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 _6599_/Q VGND VGND VPWR VPWR _3930_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6963_ _7063_/CLK _6963_/D fanout590/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_4
X_5914_ _5934_/C _6072_/C _6892_/Q _5776_/X _6956_/Q VGND VGND VPWR VPWR _5914_/X
+ sky130_fd_sc_hd__a32o_1
X_6894_ _7053_/CLK _6894_/D fanout601/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5845_ _6945_/Q _5779_/X _5841_/X _5842_/X _5844_/X VGND VGND VPWR VPWR _5845_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5776_ _6010_/D _5815_/C _5795_/D VGND VGND VPWR VPWR _5776_/X sky130_fd_sc_hd__and3_4
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4290_/Y _4391_/Y _4669_/X _4293_/Y _4280_/A VGND VGND VPWR VPWR _4731_/B
+ sky130_fd_sc_hd__o32a_1
X_4658_ _4722_/A _4674_/D VGND VGND VPWR VPWR _4658_/Y sky130_fd_sc_hd__nand2_4
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR _3327_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3609_ _7056_/Q _5512_/B _5630_/C hold28/A _3608_/X VGND VGND VPWR VPWR _3609_/X
+ sky130_fd_sc_hd__a41o_1
Xhold830 _7084_/Q VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 hold841/A VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold852 _6884_/Q VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4589_ _4751_/A _4589_/B _4589_/C VGND VGND VPWR VPWR _4591_/A sky130_fd_sc_hd__and3_1
XFILLER_89_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold863 _5619_/X VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _6643_/Q VGND VGND VPWR VPWR hold874/X sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _7030_/Q _6136_/A _6328_/A3 _6141_/X _6982_/Q VGND VGND VPWR VPWR _6328_/X
+ sky130_fd_sc_hd__a32o_1
Xhold885 _4001_/X VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _5409_/X VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6259_ _7131_/Q _6116_/X _6136_/X _7027_/Q _6258_/X VGND VGND VPWR VPWR _6264_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1530 hold75/A VGND VGND VPWR VPWR _5272_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1541 _6616_/Q VGND VGND VPWR VPWR _3950_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3960_ _6472_/A _7252_/Q VGND VGND VPWR VPWR _3968_/S sky130_fd_sc_hd__nand2_4
XFILLER_189_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3891_ _6934_/Q _3542_/B _3902_/A3 _5458_/B _6974_/Q VGND VGND VPWR VPWR _3891_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5630_ _5630_/A _6548_/B _5630_/C hold28/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__nand4_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5561_ _5557_/B _3922_/X _5565_/S hold850/X VGND VGND VPWR VPWR _5561_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7300_ _7300_/A VGND VGND VPWR VPWR _7300_/X sky130_fd_sc_hd__clkbuf_2
X_4512_ _5036_/B _4549_/D VGND VGND VPWR VPWR _4512_/Y sky130_fd_sc_hd__nand2_1
X_5492_ hold79/X hold21/X _5493_/S VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__mux2_1
Xhold104 _7067_/Q VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 hold115/A VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold126/A VGND VGND VPWR VPWR _4053_/B sky130_fd_sc_hd__buf_8
X_7231_ _3340_/A1 _7231_/D fanout613/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfrtp_1
X_4443_ _4349_/X _4412_/Y _4413_/Y _4442_/Y VGND VGND VPWR VPWR _4444_/A sky130_fd_sc_hd__a2bb2oi_1
Xhold137 _4052_/X VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold148/A VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold159 _4102_/X VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7162_ _7162_/CLK _7162_/D fanout600/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfrtp_4
X_4374_ _4656_/C _4740_/C _4848_/B VGND VGND VPWR VPWR _4704_/B sky130_fd_sc_hd__and3_2
XFILLER_171_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout606 fanout607/X VGND VGND VPWR VPWR fanout606/X sky130_fd_sc_hd__buf_8
Xfanout617 input126/X VGND VGND VPWR VPWR _4848_/A sky130_fd_sc_hd__buf_8
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6177_/A _6117_/A _6177_/C VGND VGND VPWR VPWR _6113_/X sky130_fd_sc_hd__and3_4
X_3325_ _3327_/A _3325_/B VGND VGND VPWR VPWR _3325_/Y sky130_fd_sc_hd__nand2_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7093_/CLK _7093_/D fanout591/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6044_ _5782_/C _6026_/X _6036_/X _6039_/X _6043_/X VGND VGND VPWR VPWR _6044_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _7106_/Q VGND VGND VPWR VPWR _3256_/Y sky130_fd_sc_hd__inv_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6946_ _7161_/CLK _6946_/D fanout599/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6877_ _7017_/CLK _6877_/D fanout606/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5828_ _7048_/Q _5814_/X _5815_/X _7016_/Q _5827_/X VGND VGND VPWR VPWR _5828_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5759_ _5759_/A _5759_/B VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__and2_2
XFILLER_182_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold660 _6994_/Q VGND VGND VPWR VPWR hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold671 hold671/A VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap390 _6101_/X VGND VGND VPWR VPWR _6325_/A2 sky130_fd_sc_hd__buf_8
Xhold682 _7097_/Q VGND VGND VPWR VPWR hold682/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold693 _3909_/X VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1360 _7023_/Q VGND VGND VPWR VPWR hold1360/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1371 _4108_/X VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1382 _7010_/Q VGND VGND VPWR VPWR hold894/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 _6983_/Q VGND VGND VPWR VPWR hold1393/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput209 _3279_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_175_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4090_ hold530/X _4051_/X _4092_/S VGND VGND VPWR VPWR _4090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6800_ _7218_/CLK _6800_/D fanout577/X VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_36_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4992_ _5120_/B _5231_/A _4992_/C VGND VGND VPWR VPWR _4992_/X sky130_fd_sc_hd__and3_1
X_6731_ _6889_/CLK _6731_/D fanout582/X VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3943_ _6540_/A0 hold678/X _3944_/S VGND VGND VPWR VPWR _3943_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6662_ _6855_/CLK _6662_/D fanout584/X VGND VGND VPWR VPWR _6662_/Q sky130_fd_sc_hd__dfrtp_2
X_3874_ _3874_/A _3874_/B _3874_/C _3873_/Y VGND VGND VPWR VPWR _3874_/Y sky130_fd_sc_hd__nor4b_1
XFILLER_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5613_ _3915_/B hold762/X _5619_/S VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__mux2_1
X_6593_ _7114_/CLK _6593_/D fanout604/X VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5544_ _3924_/B hold260/X hold77/X VGND VGND VPWR VPWR _5544_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5475_ _4053_/B hold161/X _5475_/S VGND VGND VPWR VPWR _5475_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7214_ _7251_/CLK _7214_/D fanout594/X VGND VGND VPWR VPWR _7214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4426_ _4848_/A _5040_/C VGND VGND VPWR VPWR _4427_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout403 _4574_/C VGND VGND VPWR VPWR _4589_/C sky130_fd_sc_hd__buf_4
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7145_ _7145_/CLK _7145_/D fanout600/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_93_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7265_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout425 _6465_/A2 VGND VGND VPWR VPWR _6138_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4357_ _5042_/A _5042_/B _5260_/A VGND VGND VPWR VPWR _4449_/A sky130_fd_sc_hd__and3_1
XFILLER_99_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout436 _4298_/X VGND VGND VPWR VPWR _4815_/A sky130_fd_sc_hd__buf_6
Xfanout458 _5657_/D VGND VGND VPWR VPWR _5575_/C sky130_fd_sc_hd__buf_8
X_3308_ _3300_/B _6442_/S _5759_/B VGND VGND VPWR VPWR _3308_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7076_ _7077_/CLK _7076_/D fanout588/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout469 hold56/A VGND VGND VPWR VPWR _5684_/B sky130_fd_sc_hd__buf_12
X_4288_ _4670_/D _4667_/C _4288_/C VGND VGND VPWR VPWR _4984_/C sky130_fd_sc_hd__and3_4
XFILLER_58_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6027_ _6028_/C _6072_/C _6680_/Q _5776_/X _6770_/Q VGND VGND VPWR VPWR _6027_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _7130_/CLK _6929_/D fanout599/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7108_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7150_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold490 _7018_/Q VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1190 _5685_/X VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_330 _7036_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 _6907_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_352 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_363 _5971_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 _3918_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 _4092_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_396 _6098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3590_ _6817_/Q _3528_/C _5281_/A2 _3588_/X _3589_/X VGND VGND VPWR VPWR _3590_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_139_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5260_ _5260_/A _5260_/B _5260_/C VGND VGND VPWR VPWR _5260_/X sky130_fd_sc_hd__and3_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4211_ _4549_/D _4632_/B _4600_/B _4612_/C VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__and4b_2
X_5191_ _5258_/A _5258_/B VGND VGND VPWR VPWR _5191_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4142_ hold982/X _6539_/A0 _4144_/S VGND VGND VPWR VPWR _4142_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4073_ _5494_/A hold64/X hold21/X VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__and3_2
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4975_ _4620_/A _4597_/C _4620_/B _4620_/X VGND VGND VPWR VPWR _4976_/D sky130_fd_sc_hd__a31o_1
X_6714_ _7120_/CLK _6714_/D fanout610/X VGND VGND VPWR VPWR _7304_/A sky130_fd_sc_hd__dfrtp_1
X_3926_ hold13/X _3913_/B _3924_/X _3914_/S hold760/X VGND VGND VPWR VPWR _3926_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6645_ _7274_/CLK _6645_/D fanout577/X VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_149_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3857_ _6917_/Q _3533_/C _5281_/A2 _5566_/B _7069_/Q VGND VGND VPWR VPWR _3857_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6576_ _7129_/CLK _6576_/D fanout598/X VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3788_ _6563_/Q _3372_/B _3954_/B _6624_/Q _3787_/X VGND VGND VPWR VPWR _3788_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_152_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5527_ hold848/X _6505_/A1 _5529_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5458_ _5494_/A _5458_/B VGND VGND VPWR VPWR _5466_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4409_ _4878_/B _4654_/B _4409_/C _4668_/C VGND VGND VPWR VPWR _4411_/B sky130_fd_sc_hd__and4_1
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5389_ hold332/X _3919_/C _5394_/S VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7128_ _7161_/CLK _7128_/D fanout599/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7059_ _7072_/CLK _7059_/D fanout596/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_160 _7191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _3349_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _6466_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_193 _5911_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4923_/B _4760_/B _4760_/C VGND VGND VPWR VPWR _4777_/C sky130_fd_sc_hd__and3_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3711_ _6691_/Q _3481_/X _6542_/B _7273_/Q _3710_/X VGND VGND VPWR VPWR _3717_/C
+ sky130_fd_sc_hd__a221o_1
X_4691_ _4777_/A _4691_/B _4706_/B VGND VGND VPWR VPWR _4778_/C sky130_fd_sc_hd__and3_4
XFILLER_119_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6430_ _6751_/Q _6098_/X _6113_/X _6636_/Q _6429_/X VGND VGND VPWR VPWR _6431_/D
+ sky130_fd_sc_hd__a221o_1
X_3642_ _7161_/Q _3509_/X _3521_/X _7169_/Q _3641_/X VGND VGND VPWR VPWR _3652_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6361_ _7239_/Q _6177_/C _6114_/X _6113_/X _6633_/Q VGND VGND VPWR VPWR _6361_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3573_ _5675_/D _5657_/D _3757_/D VGND VGND VPWR VPWR _3573_/X sky130_fd_sc_hd__and3_2
X_5312_ _5312_/A0 _4152_/B _5312_/S VGND VGND VPWR VPWR _5312_/X sky130_fd_sc_hd__mux2_1
X_6292_ _6291_/X _7211_/Q _6292_/S VGND VGND VPWR VPWR _6292_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5243_ _5243_/A _5243_/B _5243_/C VGND VGND VPWR VPWR _5243_/Y sky130_fd_sc_hd__nand3_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _4562_/A _5173_/X _5174_/C _5174_/D VGND VGND VPWR VPWR _5175_/C sky130_fd_sc_hd__and4bb_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4125_ _6546_/A0 hold546/X _4126_/S VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4056_ _5326_/A0 _6898_/Q _3346_/D _5666_/C VGND VGND VPWR VPWR _4056_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4958_ _4246_/Y _4254_/Y _4951_/X _4957_/X _5270_/D VGND VGND VPWR VPWR _4958_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3909_ _6550_/A0 hold692/X _3912_/S VGND VGND VPWR VPWR _3909_/X sky130_fd_sc_hd__mux2_1
X_4889_ _4670_/D _4859_/A _4721_/C _4626_/X VGND VGND VPWR VPWR _5225_/A sky130_fd_sc_hd__a31oi_1
XFILLER_177_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6628_ _7219_/CLK _6628_/D VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6559_ _6781_/CLK _6559_/D _3291_/A VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire442 _4170_/B VGND VGND VPWR VPWR wire442/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ _6876_/Q _5726_/Y _5917_/X _5929_/X _5759_/A VGND VGND VPWR VPWR _5930_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_34_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5861_ _6442_/S _5861_/A2 _6443_/S _5860_/X VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__a211o_1
XFILLER_178_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4812_ _5089_/C _4753_/B _4729_/A _4473_/Y VGND VGND VPWR VPWR _5040_/A sky130_fd_sc_hd__o22a_4
X_5792_ _7119_/Q _6072_/B _6025_/C VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__and3_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4743_ _4786_/B _4939_/B VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__nand2_2
XFILLER_187_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4674_ _4940_/C _5036_/C _4674_/C _4674_/D VGND VGND VPWR VPWR _4674_/X sky130_fd_sc_hd__and4_1
X_6413_ _6556_/Q _6110_/X _6410_/X _6412_/X VGND VGND VPWR VPWR _6414_/C sky130_fd_sc_hd__a211o_1
X_3625_ _7080_/Q _3413_/X _3463_/X _7112_/Q _3624_/X VGND VGND VPWR VPWR _3625_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6344_ _7260_/Q _6446_/C _6425_/C _6144_/X _6648_/Q VGND VGND VPWR VPWR _6344_/X
+ sky130_fd_sc_hd__a32o_1
X_3556_ _6725_/Q hold38/A _5295_/D _3554_/X _3555_/X VGND VGND VPWR VPWR _3556_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_115_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6275_ _6996_/Q _6176_/B _6143_/C _6129_/A _6900_/Q VGND VGND VPWR VPWR _6275_/X
+ sky130_fd_sc_hd__a32o_1
X_3487_ _6816_/Q _3528_/C _5281_/A2 _5323_/S _7175_/Q VGND VGND VPWR VPWR _3487_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4227_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_130_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5226_ _5226_/A _5226_/B _5226_/C VGND VGND VPWR VPWR _5226_/Y sky130_fd_sc_hd__nand3_1
XFILLER_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5157_ _4635_/Y _5153_/X _5248_/A3 _4956_/X _5073_/B VGND VGND VPWR VPWR _5270_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_96_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4108_ _6535_/A0 hold940/X _4108_/S VGND VGND VPWR VPWR _4108_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5088_ _5087_/Y _5038_/X _5011_/X hold37/A _4206_/B VGND VGND VPWR VPWR _6806_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4039_ _6546_/A0 hold554/X _4040_/S VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_60 _3905_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_71 _5708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _5779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 _5813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold308 _5443_/X VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold319 _5470_/X VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3410_ hold26/X hold71/X _5620_/A _5324_/B VGND VGND VPWR VPWR _3540_/B sky130_fd_sc_hd__and4b_4
X_4390_ _4632_/A _4511_/A _5036_/C VGND VGND VPWR VPWR _4519_/C sky130_fd_sc_hd__and3_2
X_3341_ _6789_/Q input93/X _6854_/Q VGND VGND VPWR VPWR _3341_/X sky130_fd_sc_hd__mux2_4
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6060_ _6641_/Q _6025_/B _5781_/X _6059_/X _6009_/C VGND VGND VPWR VPWR _6060_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _6978_/Q VGND VGND VPWR VPWR _3272_/Y sky130_fd_sc_hd__inv_2
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 _3932_/X VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _4894_/X _5010_/X _5009_/Y _4981_/X VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__o31a_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1019 _6773_/Q VGND VGND VPWR VPWR _4153_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6962_ _7037_/CLK _6962_/D fanout591/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_4
X_5913_ _7036_/Q _6072_/B _5773_/X _5912_/X VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__a31o_1
X_6893_ _7037_/CLK _6893_/D fanout591/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5844_ _7097_/Q _5780_/X _5788_/X _6993_/Q _5843_/X VGND VGND VPWR VPWR _5844_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5775_ _7180_/Q _7182_/Q _7183_/Q _7181_/Q VGND VGND VPWR VPWR _6009_/C sky130_fd_sc_hd__and4bb_4
X_4726_ _4984_/A _4970_/B VGND VGND VPWR VPWR _4726_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4657_ _4722_/A _4662_/B _4657_/C VGND VGND VPWR VPWR _4659_/B sky130_fd_sc_hd__and3_2
XFILLER_174_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_2
X_3608_ _7128_/Q _6548_/A hold39/A _3563_/X _7024_/Q VGND VGND VPWR VPWR _3608_/X
+ sky130_fd_sc_hd__a32o_1
Xhold820 _7271_/Q VGND VGND VPWR VPWR hold820/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold831 _5590_/X VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4588_ _4473_/Y _4527_/X _4567_/Y _4587_/Y VGND VGND VPWR VPWR _4591_/C sky130_fd_sc_hd__o31ai_1
XFILLER_190_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap550 _4637_/Y VGND VGND VPWR VPWR _4645_/A sky130_fd_sc_hd__clkbuf_1
Xhold842 _7132_/Q VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 _5365_/X VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap561 _4304_/Y VGND VGND VPWR VPWR _4523_/C sky130_fd_sc_hd__buf_2
Xhold864 _7172_/Q VGND VGND VPWR VPWR hold864/X sky130_fd_sc_hd__dlygate4sd3_1
X_6327_ _6974_/Q _6097_/X _6120_/X _6918_/Q _6326_/X VGND VGND VPWR VPWR _6330_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold875 _3982_/X VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmgmt_gpio_15_buff_inst _3339_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
XFILLER_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3539_ _5620_/A _5684_/B _5675_/D VGND VGND VPWR VPWR _3539_/X sky130_fd_sc_hd__and3_4
Xhold886 _6931_/Q VGND VGND VPWR VPWR hold886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _6638_/Q VGND VGND VPWR VPWR hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6258_ _7019_/Q _6177_/C _6110_/C _6451_/B1 _6915_/Q VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5209_ _5209_/A _5246_/C _5209_/C VGND VGND VPWR VPWR _5210_/C sky130_fd_sc_hd__and3_1
XFILLER_190_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6189_ _7048_/Q _6130_/A _6110_/C _6186_/X _6188_/X VGND VGND VPWR VPWR _6190_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_130_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1520 _6851_/Q VGND VGND VPWR VPWR _4055_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1531 _6583_/Q VGND VGND VPWR VPWR _3813_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _6805_/Q VGND VGND VPWR VPWR _4980_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3890_ _6998_/Q _5485_/B _5629_/C _5639_/B _7134_/Q VGND VGND VPWR VPWR _3890_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_188_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5560_ _5557_/B _3919_/X _5565_/S _5560_/B2 VGND VGND VPWR VPWR _5560_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4511_ _4511_/A _4689_/B VGND VGND VPWR VPWR _4755_/D sky130_fd_sc_hd__nor2_4
X_5491_ hold803/X _6505_/A1 _5493_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
Xhold105 _5571_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7230_ _7254_/CLK _7230_/D fanout613/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__dfrtp_1
Xhold116 hold116/A VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4442_ _4442_/A _4442_/B _4442_/C _4442_/D VGND VGND VPWR VPWR _4442_/Y sky130_fd_sc_hd__nand4_1
Xhold127 _5303_/X VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _6812_/Q VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _6948_/Q VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlygate4sd3_1
X_7161_ _7161_/CLK _7161_/D fanout600/X VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_2
X_4373_ _4689_/B _4761_/C _4209_/Y _4369_/X _4848_/A VGND VGND VPWR VPWR _4849_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6143_/D _6141_/B _6112_/C VGND VGND VPWR VPWR _6112_/X sky130_fd_sc_hd__and3_4
Xfanout607 fanout611/X VGND VGND VPWR VPWR fanout607/X sky130_fd_sc_hd__buf_6
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3324_ _6861_/Q input89/X _3327_/A VGND VGND VPWR VPWR _3324_/X sky130_fd_sc_hd__mux2_2
Xfanout618 _4706_/B VGND VGND VPWR VPWR _4647_/C sky130_fd_sc_hd__buf_12
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7145_/CLK _7092_/D fanout602/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _7277_/Q _6086_/B1 _5784_/X _6622_/Q _6042_/X VGND VGND VPWR VPWR _6043_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _7114_/Q VGND VGND VPWR VPWR _3255_/Y sky130_fd_sc_hd__inv_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6945_/CLK hold68/X fanout583/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6876_ _7108_/CLK _6876_/D fanout606/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_4
X_5827_ _7008_/Q _5783_/X _5791_/X _7120_/Q _5826_/X VGND VGND VPWR VPWR _5827_/X
+ sky130_fd_sc_hd__a221o_1
X_5758_ _5758_/A0 _5757_/X _5758_/S VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4709_ _4945_/C _4792_/C VGND VGND VPWR VPWR _4709_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5689_ _5689_/A0 hold5/X _5692_/S VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__mux2_1
XFILLER_147_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold650 hold650/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xhold661 _5489_/X VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _7025_/Q VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold683 _5605_/X VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap391 _6096_/Y VGND VGND VPWR VPWR _6328_/A3 sky130_fd_sc_hd__buf_2
Xhold694 hold694/A VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1350 _5603_/X VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 _5522_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1372 _6733_/Q VGND VGND VPWR VPWR hold1372/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 _6829_/Q VGND VGND VPWR VPWR hold1383/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _6952_/Q VGND VGND VPWR VPWR hold401/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4991_ _4859_/C _4862_/A _4859_/D _4673_/X _4988_/X VGND VGND VPWR VPWR _4991_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6730_ _6855_/CLK hold95/X fanout583/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dfstp_2
XFILLER_189_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3942_ _3919_/C hold389/X _3944_/S VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__mux2_1
X_6661_ _6780_/CLK _6661_/D fanout575/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfrtp_4
X_3873_ _3873_/A _3873_/B _3873_/C _3873_/D VGND VGND VPWR VPWR _3873_/Y sky130_fd_sc_hd__nor4_1
X_5612_ _6549_/A0 _5612_/A1 _5619_/S VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__mux2_1
X_6592_ _7072_/CLK _6592_/D fanout599/X VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5543_ _3921_/X _5543_/A1 hold77/X VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__mux2_1
X_5474_ _4051_/B hold674/X _5475_/S VGND VGND VPWR VPWR _5474_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7213_ _7254_/CLK _7213_/D fanout595/X VGND VGND VPWR VPWR _7213_/Q sky130_fd_sc_hd__dfrtp_1
X_4425_ _4751_/A _4429_/A _5055_/D _4429_/D VGND VGND VPWR VPWR _4488_/C sky130_fd_sc_hd__and4_1
XFILLER_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7144_ _7160_/CLK _7144_/D fanout592/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfstp_2
Xfanout404 _5255_/B VGND VGND VPWR VPWR _4738_/B sky130_fd_sc_hd__buf_8
X_4356_ _4356_/A _4848_/A _4427_/D VGND VGND VPWR VPWR _4356_/Y sky130_fd_sc_hd__nand3_4
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout426 _5733_/Y VGND VGND VPWR VPWR _6465_/A2 sky130_fd_sc_hd__buf_12
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3307_ _6442_/S _3307_/B VGND VGND VPWR VPWR _3307_/Y sky130_fd_sc_hd__nand2_1
Xfanout459 hold43/X VGND VGND VPWR VPWR _5657_/D sky130_fd_sc_hd__buf_12
X_7075_ _7108_/CLK hold19/X fanout607/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_4
X_4287_ _4214_/A _4214_/B _4285_/A _4637_/A VGND VGND VPWR VPWR _4667_/D sky130_fd_sc_hd__a22oi_4
XFILLER_101_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6026_ _6813_/Q _6028_/C _5795_/C VGND VGND VPWR VPWR _6026_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _7114_/CLK _6928_/D fanout604/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6859_ _7122_/CLK _6859_/D fanout606/X VGND VGND VPWR VPWR _7307_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold480 _6973_/Q VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold491 _5516_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1180 _6854_/Q VGND VGND VPWR VPWR _5330_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _7287_/A VGND VGND VPWR VPWR _4174_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_320 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_331 _6598_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_342 _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 _3327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_364 _6086_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 hold65/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_386 _3915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _6098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4210_ _4632_/A _5036_/B VGND VGND VPWR VPWR _4801_/A sky130_fd_sc_hd__nor2_4
X_5190_ _5060_/A _4505_/B _4718_/D _4488_/X _5189_/Y VGND VGND VPWR VPWR _5190_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_141_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4141_ hold411/X _6538_/A0 _4144_/S VGND VGND VPWR VPWR _4141_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4072_ _6505_/A1 hold870/X hold57/X VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4974_ _4511_/A _4970_/D _4633_/B _4735_/Y _4973_/Y VGND VGND VPWR VPWR _4974_/X
+ sky130_fd_sc_hd__o41a_1
X_3925_ _5494_/A hold64/X _3925_/C VGND VGND VPWR VPWR _3925_/X sky130_fd_sc_hd__and3_4
X_6713_ _7120_/CLK _6713_/D fanout610/X VGND VGND VPWR VPWR _7303_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6644_ _7279_/CLK _6644_/D fanout597/X VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3856_ _3856_/A _3856_/B _3856_/C _3856_/D VGND VGND VPWR VPWR _3875_/A sky130_fd_sc_hd__nor4_4
XFILLER_137_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6575_ _7129_/CLK _6575_/D fanout598/X VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfrtp_4
X_3787_ _6827_/Q _3497_/X _3531_/X _6757_/Q VGND VGND VPWR VPWR _3787_/X sky130_fd_sc_hd__a22o_1
X_5526_ hold698/X _3924_/B _5529_/S VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5457_ hold218/X _4053_/B _5457_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4408_ _4363_/A _4722_/A _4675_/A _4870_/C _4683_/C VGND VGND VPWR VPWR _4408_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_182_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5388_ hold299/X _6550_/A0 _5394_/S VGND VGND VPWR VPWR _5388_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7127_ _7154_/CLK _7127_/D fanout593/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_113_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4339_ _4597_/B _4509_/D _4509_/A VGND VGND VPWR VPWR _4595_/A sky130_fd_sc_hd__and3_4
XFILLER_47_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7058_ _7170_/CLK _7058_/D fanout605/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6009_ _6649_/Q _6059_/S _6009_/C VGND VGND VPWR VPWR _6009_/X sky130_fd_sc_hd__and3_1
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 _6935_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _6440_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_194 _5911_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_92_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6827_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _6930_/Q _3533_/C _3902_/A3 _3497_/X _6826_/Q VGND VGND VPWR VPWR _3710_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4690_ _4712_/B _4687_/B _4689_/X _4688_/Y VGND VGND VPWR VPWR _4690_/Y sky130_fd_sc_hd__a211oi_1
X_3641_ _6840_/Q _5666_/C hold39/A _3432_/X _6604_/Q VGND VGND VPWR VPWR _3641_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6360_ _6658_/Q _6129_/B _6116_/X _6569_/Q _6359_/X VGND VGND VPWR VPWR _6365_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3572_ _6839_/Q _5666_/C hold39/A _3492_/X _6664_/Q VGND VGND VPWR VPWR _3572_/X
+ sky130_fd_sc_hd__a32o_2
X_5311_ _6536_/B _5311_/B _5311_/C VGND VGND VPWR VPWR _5312_/S sky130_fd_sc_hd__and3_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6291_ _6285_/Y _6290_/Y _6876_/Q _6134_/Y VGND VGND VPWR VPWR _6291_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_142_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5242_ _5238_/Y _5262_/B _5235_/X VGND VGND VPWR VPWR _5243_/C sky130_fd_sc_hd__a21bo_1
XFILLER_69_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7131_/CLK sky130_fd_sc_hd__clkbuf_16
X_5173_ _5263_/A _5263_/B _5173_/C VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__and3_1
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4124_ _6539_/A0 _4124_/A1 _4126_/S VGND VGND VPWR VPWR _4124_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_4
X_4055_ _4055_/A1 _3249_/A _3346_/D _5666_/C VGND VGND VPWR VPWR _4055_/X sky130_fd_sc_hd__o31a_1
XFILLER_37_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7173_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4957_ _4643_/Y _4951_/X _4955_/X _4956_/X VGND VGND VPWR VPWR _4957_/X sky130_fd_sc_hd__o211a_1
XFILLER_51_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3908_ _6543_/A0 hold350/X _3912_/S VGND VGND VPWR VPWR _3908_/X sky130_fd_sc_hd__mux2_1
X_4888_ _4888_/A _5228_/A _4888_/C VGND VGND VPWR VPWR _4890_/A sky130_fd_sc_hd__and3_1
X_3839_ _5331_/C _4139_/C _3344_/X _3428_/X _7012_/Q VGND VGND VPWR VPWR _3839_/X
+ sky130_fd_sc_hd__a32o_1
X_6627_ _7219_/CLK _6627_/D VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6558_ _7270_/CLK _6558_/D fanout579/X VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5509_ _4049_/B hold338/X _5511_/S VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6489_ _6489_/A1 _4166_/B _6488_/X VGND VGND VPWR VPWR _6489_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire410 _3412_/X VGND VGND VPWR VPWR _5440_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_168_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5860_ _5726_/Y _6873_/Q _5859_/X _5849_/X _5759_/A VGND VGND VPWR VPWR _5860_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4811_ _5040_/C _4265_/Y _4348_/X _5131_/A VGND VGND VPWR VPWR _4811_/X sky130_fd_sc_hd__o31a_1
XFILLER_178_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5791_ _5965_/B _5911_/C VGND VGND VPWR VPWR _5791_/X sky130_fd_sc_hd__and2_2
X_4742_ _4786_/B _4760_/B _4742_/C VGND VGND VPWR VPWR _4775_/B sky130_fd_sc_hd__and3_1
XFILLER_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4673_ _4984_/A _4675_/B _4732_/C VGND VGND VPWR VPWR _4673_/X sky130_fd_sc_hd__and3_1
XFILLER_174_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6412_ _7267_/Q _6106_/X _6109_/X _6599_/Q _6411_/X VGND VGND VPWR VPWR _6412_/X
+ sky130_fd_sc_hd__a221o_1
X_3624_ _7040_/Q _5548_/C _5281_/A2 _3623_/X VGND VGND VPWR VPWR _3624_/X sky130_fd_sc_hd__a31o_1
XFILLER_147_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6343_ _6342_/X _6343_/A1 _6343_/S VGND VGND VPWR VPWR _7214_/D sky130_fd_sc_hd__mux2_1
X_3555_ _6837_/Q _5295_/D _3446_/X _4139_/C _5311_/C VGND VGND VPWR VPWR _3555_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6274_ _7124_/Q _5750_/X _6325_/A2 _6884_/Q _6273_/X VGND VGND VPWR VPWR _6285_/A
+ sky130_fd_sc_hd__a221o_1
X_3486_ _6548_/C _5327_/D _6536_/D VGND VGND VPWR VPWR _5323_/S sky130_fd_sc_hd__and3_4
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5225_ _5225_/A _5225_/B _5225_/C _5225_/D VGND VGND VPWR VPWR _5226_/C sky130_fd_sc_hd__and4_1
XFILLER_102_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5156_ _5152_/X _5204_/B _5204_/C VGND VGND VPWR VPWR _5159_/A sky130_fd_sc_hd__and3b_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4107_ _6546_/A0 hold439/X _4108_/S VGND VGND VPWR VPWR _4107_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5087_ _5087_/A _5087_/B VGND VGND VPWR VPWR _5087_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4038_ _3919_/C hold354/X _4040_/S VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5989_ _6607_/Q _6025_/B _6003_/C _5988_/X VGND VGND VPWR VPWR _5989_/X sky130_fd_sc_hd__a31o_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_50 _3548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_61 _3905_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _5708_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_83 _5782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 _5836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput190 _3262_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_153_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold309 hold309/A VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3340_ _6790_/Q _3340_/A1 _6852_/Q VGND VGND VPWR VPWR _3340_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _6986_/Q VGND VGND VPWR VPWR _3271_/Y sky130_fd_sc_hd__inv_2
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4815_/A _4923_/B _5128_/C _5128_/A VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__o211a_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 hold1421/X VGND VGND VPWR VPWR _6521_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6961_ _7073_/CLK _6961_/D fanout585/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5912_ _6916_/Q _6028_/B _5934_/C VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__and3_1
X_6892_ _7160_/CLK _6892_/D fanout592/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_4
X_5843_ _7121_/Q _6059_/S _5911_/C _5784_/X _7025_/Q VGND VGND VPWR VPWR _5843_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5774_ _5814_/C _5934_/C _5782_/C VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__and3_4
X_4725_ _5128_/A _4519_/C _4729_/D _4724_/Y VGND VGND VPWR VPWR _4731_/A sky130_fd_sc_hd__a31oi_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4656_ _4698_/A _4657_/C _4656_/C VGND VGND VPWR VPWR _4750_/B sky130_fd_sc_hd__and3b_1
XFILLER_175_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3607_ _6952_/Q _5273_/D _5440_/C _6560_/Q _3372_/B VGND VGND VPWR VPWR _3607_/X
+ sky130_fd_sc_hd__a32o_1
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _3352_/B sky130_fd_sc_hd__buf_2
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_4
Xhold810 _5653_/X VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 _6544_/X VGND VGND VPWR VPWR _7271_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4587_ _4587_/A _4587_/B VGND VGND VPWR VPWR _4587_/Y sky130_fd_sc_hd__nor2_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR _3325_/B sky130_fd_sc_hd__clkbuf_2
Xhold832 hold832/A VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 _5645_/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap551 _4853_/C VGND VGND VPWR VPWR _4791_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_190_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap562 _4277_/Y VGND VGND VPWR VPWR _4280_/A sky130_fd_sc_hd__buf_6
Xhold854 _6920_/Q VGND VGND VPWR VPWR hold854/X sky130_fd_sc_hd__dlygate4sd3_1
X_3538_ _5620_/A _5512_/B hold27/A VGND VGND VPWR VPWR _3538_/X sky130_fd_sc_hd__and3_1
X_6326_ _6998_/Q _6176_/B _6347_/C _6103_/X _7070_/Q VGND VGND VPWR VPWR _6326_/X
+ sky130_fd_sc_hd__a32o_1
Xhold865 _5690_/X VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _7154_/Q VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold887 _5418_/X VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 _3976_/X VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6257_ _7123_/Q _5750_/X _6129_/C _7155_/Q _6256_/X VGND VGND VPWR VPWR _6264_/A
+ sky130_fd_sc_hd__a221o_1
X_3469_ _4127_/C _5476_/C _3528_/C VGND VGND VPWR VPWR _3469_/X sky130_fd_sc_hd__and3_2
XFILLER_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5208_ _4945_/B _4792_/B _4789_/D _5207_/X VGND VGND VPWR VPWR _5209_/C sky130_fd_sc_hd__a31oi_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6188_ _7112_/Q _6110_/X _6112_/X _7104_/Q _6187_/X VGND VGND VPWR VPWR _6188_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1510 _7218_/Q VGND VGND VPWR VPWR _6467_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 _7197_/Q VGND VGND VPWR VPWR _5886_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1532 _7212_/Q VGND VGND VPWR VPWR _6293_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5139_ _4277_/Y _4398_/X _4403_/X _5048_/X _5138_/X VGND VGND VPWR VPWR _5142_/B
+ sky130_fd_sc_hd__o311a_1
Xhold1543 _7259_/Q VGND VGND VPWR VPWR _7250_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _4606_/B _4586_/B VGND VGND VPWR VPWR _4510_/Y sky130_fd_sc_hd__nand2_2
X_5490_ hold254/X _3924_/B _5493_/S VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold106 _6940_/Q VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _4441_/A _4441_/B _4441_/C VGND VGND VPWR VPWR _4442_/A sky130_fd_sc_hd__nor3_1
Xhold117 _7053_/Q VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold128 _6870_/Q VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold139 _5275_/X VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ _7160_/CLK _7160_/D fanout592/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfstp_2
X_4372_ _4761_/C _4280_/A _4691_/B VGND VGND VPWR VPWR _4372_/Y sky130_fd_sc_hd__o21ai_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _7186_/Q _7190_/Q _7189_/Q _7185_/Q VGND VGND VPWR VPWR _6112_/C sky130_fd_sc_hd__and4bb_2
Xfanout608 fanout611/X VGND VGND VPWR VPWR fanout608/X sky130_fd_sc_hd__buf_6
X_3323_ _6862_/Q input91/X _3327_/A VGND VGND VPWR VPWR _3323_/X sky130_fd_sc_hd__mux2_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7130_/CLK hold15/X fanout600/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout619 _4494_/C VGND VGND VPWR VPWR _4600_/B sky130_fd_sc_hd__buf_6
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6556_/Q _5767_/X _5780_/X _7272_/Q _6041_/X VGND VGND VPWR VPWR _6042_/X
+ sky130_fd_sc_hd__a221o_1
X_3254_ _7122_/Q VGND VGND VPWR VPWR _3254_/Y sky130_fd_sc_hd__inv_2
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6944_ _6967_/CLK _6944_/D fanout586/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6875_ _6875_/CLK _6875_/D fanout598/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfrtp_4
X_5826_ _7064_/Q _5826_/B _6010_/C _6010_/D VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__and4_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5757_ _7177_/Q _7176_/Q _5757_/C _6803_/Q VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__and4b_1
XFILLER_108_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4708_ _4708_/A _4792_/C VGND VGND VPWR VPWR _4711_/B sky130_fd_sc_hd__nand2_1
XFILLER_148_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5688_ hold363/X _3921_/B _5692_/S VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4639_ _4722_/A _4777_/A _4945_/C VGND VGND VPWR VPWR _4641_/B sky130_fd_sc_hd__and3_1
XFILLER_163_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold640 _4149_/X VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 _7081_/Q VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _7245_/Q VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _5524_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6309_ _6901_/Q _6129_/A _6454_/B1 _6957_/Q _6308_/X VGND VGND VPWR VPWR _6314_/B
+ sky130_fd_sc_hd__a221o_1
Xhold684 _7261_/Q VGND VGND VPWR VPWR hold684/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold695 hold695/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
X_7289_ _7289_/A VGND VGND VPWR VPWR _7289_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1340 _7087_/Q VGND VGND VPWR VPWR hold966/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 _6734_/Q VGND VGND VPWR VPWR hold371/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1362 _6887_/Q VGND VGND VPWR VPWR hold1362/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1373 _4104_/X VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 _6732_/Q VGND VGND VPWR VPWR _4102_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1395 _5442_/X VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4990_ _4719_/B _4903_/B _4851_/X _4987_/X _4989_/X VGND VGND VPWR VPWR _4992_/C
+ sky130_fd_sc_hd__a2111oi_1
X_3941_ _6538_/A0 hold446/X _3944_/S VGND VGND VPWR VPWR _3941_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6660_ _7239_/CLK _6660_/D fanout573/X VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfstp_1
X_3872_ _7013_/Q _3428_/X _5639_/B _7133_/Q _3871_/X VGND VGND VPWR VPWR _3873_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5611_ hold13/X _5611_/B VGND VGND VPWR VPWR _5619_/S sky130_fd_sc_hd__nand2_4
X_6591_ _7278_/CLK _6591_/D fanout597/X VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5542_ hold2/X hold186/X hold77/X VGND VGND VPWR VPWR _5542_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5473_ _4049_/B hold502/X _5475_/S VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7212_ _7259_/CLK _7212_/D fanout595/X VGND VGND VPWR VPWR _7212_/Q sky130_fd_sc_hd__dfrtp_1
X_4424_ _4939_/A _4945_/B VGND VGND VPWR VPWR _4752_/A sky130_fd_sc_hd__nand2_1
XFILLER_145_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7143_ _7143_/CLK _7143_/D fanout587/X VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfstp_1
X_4355_ _4356_/A _4848_/A _4427_/D VGND VGND VPWR VPWR _5260_/A sky130_fd_sc_hd__and3_2
Xfanout405 _4460_/C VGND VGND VPWR VPWR _5260_/B sky130_fd_sc_hd__buf_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout427 _5732_/X VGND VGND VPWR VPWR _6136_/A sky130_fd_sc_hd__buf_12
XFILLER_59_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3306_ _6800_/Q _6850_/Q _3300_/Y _3305_/Y VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__a22o_1
X_7074_ _7161_/CLK _7074_/D fanout600/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4286_ _4346_/A _4285_/A _4288_/C VGND VGND VPWR VPWR _4625_/B sky130_fd_sc_hd__o21ai_1
XFILLER_140_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6025_ _6561_/Q _6025_/B _6025_/C VGND VGND VPWR VPWR _6025_/X sky130_fd_sc_hd__and3_1
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _7159_/CLK _6927_/D fanout599/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_120_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6858_ _7099_/CLK _6858_/D fanout598/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfrtp_1
X_5809_ _7055_/Q _7181_/Q _7180_/Q _5814_/C _5808_/X VGND VGND VPWR VPWR _5809_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_167_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6789_ _7053_/CLK _6789_/D fanout601/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold470 hold470/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_145_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold481 _5465_/X VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold492 _6896_/Q VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1170 _3914_/X VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1181 _5330_/X VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 _4174_/X VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_310 _6122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _6954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_332 _7068_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_343 _6781_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_354 _3313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_365 _6086_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 hold83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_387 _3918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_398 _6098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4140_ _4140_/A0 _4152_/B _4144_/S VGND VGND VPWR VPWR _4140_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4071_ hold8/X _3539_/X _3924_/X hold57/X hold619/X VGND VGND VPWR VPWR _4071_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_49_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4973_ _4973_/A _4973_/B _4973_/C VGND VGND VPWR VPWR _4973_/Y sky130_fd_sc_hd__nor3_1
X_6712_ _7123_/CLK hold58/X fanout610/X VGND VGND VPWR VPWR _7302_/A sky130_fd_sc_hd__dfrtp_1
X_3924_ hold65/X _3924_/B VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__and2_4
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6643_ _7270_/CLK _6643_/D fanout579/X VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfrtp_4
X_3855_ _7053_/Q _3548_/X _3852_/X _3854_/X VGND VGND VPWR VPWR _3856_/D sky130_fd_sc_hd__a211o_1
X_3786_ _7019_/Q _3563_/A _5440_/C _3782_/X _3785_/X VGND VGND VPWR VPWR _3810_/B
+ sky130_fd_sc_hd__a311o_1
X_6574_ _7240_/CLK _6574_/D fanout596/X VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5525_ hold381/X _3921_/B _5529_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5456_ hold680/X _4051_/B _5457_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4407_ _4668_/C _4409_/C _4654_/B VGND VGND VPWR VPWR _4987_/A sky130_fd_sc_hd__and3_2
X_5387_ _5387_/A0 _5649_/A0 _5394_/S VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7126_ _7132_/CLK _7126_/D fanout611/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_4
X_4338_ _4208_/Y _4246_/Y _4940_/C _4327_/Y _4509_/B VGND VGND VPWR VPWR _4597_/B
+ sky130_fd_sc_hd__o311a_4
XFILLER_113_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7057_ _7167_/CLK _7057_/D fanout604/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_4
X_4269_ _4689_/B _5036_/B VGND VGND VPWR VPWR _4970_/A sky130_fd_sc_hd__nand2_1
X_6008_ _6764_/Q _5770_/X _5793_/X _6749_/Q _6007_/X VGND VGND VPWR VPWR _6008_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _6636_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_151 _6656_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _7259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _6452_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _6028_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3640_ input45/X _4204_/S _3550_/X _7153_/Q _3639_/X VGND VGND VPWR VPWR _3652_/B
+ sky130_fd_sc_hd__a221o_2
X_3571_ _5630_/C _5476_/C _5311_/C VGND VGND VPWR VPWR _3571_/X sky130_fd_sc_hd__and3_4
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5310_ hold130/X _3922_/C hold40/X VGND VGND VPWR VPWR _5310_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6290_ _6339_/D _6290_/B _6290_/C _6290_/D VGND VGND VPWR VPWR _6290_/Y sky130_fd_sc_hd__nor4_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5241_ _5141_/X _5241_/B _5241_/C _5241_/D VGND VGND VPWR VPWR _5262_/B sky130_fd_sc_hd__and4b_1
XFILLER_69_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5172_ _5089_/X _5102_/Y _5172_/C _5217_/C VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__and4bb_1
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4123_ _6538_/A0 hold440/X _4126_/S VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4054_ hold174/X _4053_/B _4054_/S VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__mux2_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4956_ _4601_/Y _5248_/A3 _4643_/Y _4940_/Y _4635_/Y VGND VGND VPWR VPWR _4956_/X
+ sky130_fd_sc_hd__o32a_1
X_3907_ hold12/X _3907_/B VGND VGND VPWR VPWR _3912_/S sky130_fd_sc_hd__nand2_4
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4887_ _5040_/B _4376_/Y _4715_/Y _4720_/B VGND VGND VPWR VPWR _4888_/C sky130_fd_sc_hd__o31a_1
XFILLER_177_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6626_ _7219_/CLK _6626_/D VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfxtp_1
X_3838_ _7004_/Q _3438_/X _3469_/X input8/X _3837_/X VGND VGND VPWR VPWR _3843_/B
+ sky130_fd_sc_hd__a221o_1
X_6557_ _6761_/CLK _6557_/D _3291_/A VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfrtp_4
X_3769_ _6931_/Q _3542_/B _3902_/A3 _3498_/X _6767_/Q VGND VGND VPWR VPWR _3769_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5508_ _3924_/B hold278/X _5511_/S VGND VGND VPWR VPWR _5508_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6488_ _7259_/Q _6488_/A2 _6487_/X VGND VGND VPWR VPWR _6488_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5439_ _4053_/B hold204/X hold67/X VGND VGND VPWR VPWR _5439_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7163_/CLK hold33/X fanout608/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4810_ _4751_/A _4597_/C _5143_/D _5060_/B _4475_/B VGND VGND VPWR VPWR _5131_/A
+ sky130_fd_sc_hd__o2111ai_2
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _6991_/Q _5934_/C _6025_/C _5970_/B1 _6927_/Q VGND VGND VPWR VPWR _5790_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4737_/Y _4739_/Y _4740_/Y _4623_/Y VGND VGND VPWR VPWR _4808_/B sky130_fd_sc_hd__a31oi_1
XFILLER_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4672_ _4672_/A _4672_/B _4672_/C _4672_/D VGND VGND VPWR VPWR _4678_/C sky130_fd_sc_hd__nand4_1
XFILLER_174_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6411_ _6589_/Q _6138_/A _6110_/C _6107_/X _6813_/Q VGND VGND VPWR VPWR _6411_/X
+ sky130_fd_sc_hd__a32o_1
X_3623_ _6812_/Q _5341_/A _5485_/B _5404_/B _6920_/Q VGND VGND VPWR VPWR _3623_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6342_ _6292_/S _7213_/Q _6340_/Y _6341_/X VGND VGND VPWR VPWR _6342_/X sky130_fd_sc_hd__a22o_1
X_3554_ _6842_/Q _5311_/B _5295_/D VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__and3_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3485_ _3485_/A _3485_/B _3485_/C _3485_/D VGND VGND VPWR VPWR _3508_/C sky130_fd_sc_hd__nor4_2
X_6273_ _7068_/Q _6465_/A2 _6102_/X _6323_/B1 _6964_/Q VGND VGND VPWR VPWR _6273_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5224_ _4751_/A _4970_/B _5007_/A _5007_/C _5008_/X VGND VGND VPWR VPWR _5225_/D
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5155_ _4946_/X _4613_/Y _4599_/Y _5248_/A3 _4663_/Y VGND VGND VPWR VPWR _5204_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4106_ _6539_/A0 hold974/X _4111_/S VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__mux2_1
X_5086_ _5084_/X _5085_/X _4206_/B _5064_/X VGND VGND VPWR VPWR _5087_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4037_ _6538_/A0 hold504/X _4040_/S VGND VGND VPWR VPWR _4037_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _6663_/Q _6028_/B _6028_/C VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__and3_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4939_ _4939_/A _4939_/B VGND VGND VPWR VPWR _4939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_40 _3496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _5593_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _3915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_73 _5750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _5782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _7264_/CLK _6609_/D fanout579/X VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_95 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput180 _3271_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput191 _3261_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_91_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6828_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_44_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7156_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _6994_/Q VGND VGND VPWR VPWR _3270_/Y sky130_fd_sc_hd__inv_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7093_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6960_ _7151_/CLK _6960_/D fanout586/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5911_ _7124_/Q _5965_/B _5911_/C VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__and3_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6891_ _7133_/CLK _6891_/D fanout601/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfrtp_4
X_5842_ _7113_/Q _6025_/B _5842_/C VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__and3_1
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ _7183_/Q _7182_/Q _6010_/C VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__and3b_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4724_ _4479_/Y _4514_/Y _4723_/Y VGND VGND VPWR VPWR _4724_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4655_ _4939_/A _4984_/B _4984_/C _4982_/D VGND VGND VPWR VPWR _4672_/B sky130_fd_sc_hd__nand4_1
XFILLER_147_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
Xhold800 _6657_/Q VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__dlygate4sd3_1
X_3606_ _6689_/Q _5341_/A _5327_/D _3359_/B _6555_/Q VGND VGND VPWR VPWR _3606_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_128_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold811 _6898_/Q VGND VGND VPWR VPWR _3249_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_2
Xinput82 spi_sdoenb VGND VGND VPWR VPWR _3329_/A sky130_fd_sc_hd__buf_2
X_4586_ _4815_/A _4586_/B _4923_/A _4589_/C VGND VGND VPWR VPWR _4587_/A sky130_fd_sc_hd__and4_1
Xhold822 _6606_/Q VGND VGND VPWR VPWR hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_4
Xhold833 _7116_/Q VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 _6860_/Q VGND VGND VPWR VPWR hold844/X sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _6886_/Q _6325_/A2 _6104_/X _7166_/Q _6324_/X VGND VGND VPWR VPWR _6330_/B
+ sky130_fd_sc_hd__a221o_1
Xmax_cap552 _4748_/B VGND VGND VPWR VPWR _4853_/C sky130_fd_sc_hd__clkbuf_2
Xhold855 _5406_/X VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3537_ _6569_/Q _6536_/A _5341_/A _3536_/X _6983_/Q VGND VGND VPWR VPWR _3537_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_1_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold866 _7270_/Q VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold877 _5670_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _7119_/Q VGND VGND VPWR VPWR hold888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 _6777_/Q VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _7171_/Q _6130_/A _6114_/X _6325_/A2 _6883_/Q VGND VGND VPWR VPWR _6256_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_170_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3468_ _7111_/Q _3463_/X _5639_/B _7127_/Q _3467_/X VGND VGND VPWR VPWR _3485_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5207_ _4689_/C _4792_/B _4788_/A _4792_/A VGND VGND VPWR VPWR _5207_/X sky130_fd_sc_hd__o211a_1
X_6187_ _7072_/Q _6425_/B _6139_/X _6137_/X _7096_/Q VGND VGND VPWR VPWR _6187_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1500 _3445_/X VGND VGND VPWR VPWR _5372_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3399_ _6550_/A0 hold731/X _3402_/S VGND VGND VPWR VPWR _3399_/X sky130_fd_sc_hd__mux2_1
Xhold1511 _7209_/Q VGND VGND VPWR VPWR _6242_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _7190_/Q VGND VGND VPWR VPWR _5752_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1533 _7204_/Q VGND VGND VPWR VPWR _6047_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5138_ _4299_/Y _4391_/Y _4490_/Y _4414_/X VGND VGND VPWR VPWR _5138_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1544 _7201_/Q VGND VGND VPWR VPWR _5977_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5069_ _4645_/A _4947_/X _5065_/X _5067_/X _5068_/X VGND VGND VPWR VPWR _5069_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_25_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4440_ _4440_/A _4440_/B _4440_/C _4440_/D VGND VGND VPWR VPWR _4441_/C sky130_fd_sc_hd__nand4_1
Xhold107 _5428_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold118 _5555_/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _5349_/X VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4371_ _4689_/B _4427_/D _4369_/X VGND VGND VPWR VPWR _4371_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_172_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6110_ _6143_/D _6141_/B _6110_/C VGND VGND VPWR VPWR _6110_/X sky130_fd_sc_hd__and3_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3300_/Y _6177_/A _6444_/B _3296_/Y _3322_/B2 VGND VGND VPWR VPWR _6803_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_140_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7111_/CLK _7090_/D fanout600/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout609 fanout611/X VGND VGND VPWR VPWR fanout609/X sky130_fd_sc_hd__buf_6
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _7262_/Q _5777_/X _5813_/X _6566_/Q _6040_/X VGND VGND VPWR VPWR _6041_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ hold52/A VGND VGND VPWR VPWR _3253_/Y sky130_fd_sc_hd__inv_2
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6943_ _7159_/CLK _6943_/D fanout599/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6874_ _7129_/CLK _6874_/D fanout604/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5825_ _7080_/Q _5965_/B _6009_/C VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__and3_1
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ _5756_/A1 _5758_/S _5755_/Y VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__o21a_1
XFILLER_182_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4707_ _4722_/A _4730_/A VGND VGND VPWR VPWR _4707_/Y sky130_fd_sc_hd__nand2_4
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5687_ _5687_/A0 hold2/X _5692_/S VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__mux2_1
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4638_ _4940_/A _4940_/D VGND VGND VPWR VPWR _4638_/Y sky130_fd_sc_hd__nand2_4
XFILLER_118_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold630 hold630/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4569_ _5140_/C _4923_/A _4606_/D _4589_/C VGND VGND VPWR VPWR _4570_/B sky130_fd_sc_hd__and4_1
Xhold641 _7129_/Q VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _5587_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold663 _6526_/X VGND VGND VPWR VPWR _7245_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _6981_/Q VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ hold79/A _6176_/B _6143_/C _6110_/X _7117_/Q VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a32o_1
Xmax_cap382 _4730_/C VGND VGND VPWR VPWR _4738_/A sky130_fd_sc_hd__clkbuf_1
Xhold685 _6532_/X VGND VGND VPWR VPWR _7261_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap393 _6096_/Y VGND VGND VPWR VPWR wire392/A sky130_fd_sc_hd__buf_4
X_7288_ _7288_/A VGND VGND VPWR VPWR _7288_/X sky130_fd_sc_hd__clkbuf_1
Xhold696 _6917_/Q VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6239_ _6239_/A _6239_/B _6239_/C _6339_/D VGND VGND VPWR VPWR _6239_/Y sky130_fd_sc_hd__nor4_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 _7057_/Q VGND VGND VPWR VPWR hold1330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 _6833_/Q VGND VGND VPWR VPWR _5300_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 _4105_/X VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 _5369_/X VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1374 _7008_/Q VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _7039_/Q VGND VGND VPWR VPWR hold1385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 _7096_/Q VGND VGND VPWR VPWR hold783/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3940_ _4152_/B _3940_/A1 _3944_/S VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3871_ _6835_/Q _5325_/C _5311_/C _7005_/Q _3438_/X VGND VGND VPWR VPWR _3871_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5610_ _6511_/A1 hold297/X _5610_/S VGND VGND VPWR VPWR _5610_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6590_ _7275_/CLK _6590_/D fanout596/X VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5541_ _3915_/B hold248/X hold77/X VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5472_ _3925_/C hold424/X _5475_/S VGND VGND VPWR VPWR _5472_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7211_ _7254_/CLK _7211_/D fanout595/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfrtp_1
X_4423_ _4730_/A _4699_/B VGND VGND VPWR VPWR _4423_/Y sky130_fd_sc_hd__nand2_4
X_7142_ _7160_/CLK _7142_/D fanout592/X VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_4
X_4354_ _4860_/C _4860_/B VGND VGND VPWR VPWR _5040_/B sky130_fd_sc_hd__nand2_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout417 _6145_/C VGND VGND VPWR VPWR _6177_/C sky130_fd_sc_hd__buf_12
Xfanout428 _5720_/Y VGND VGND VPWR VPWR _5795_/C sky130_fd_sc_hd__buf_12
X_3305_ _6177_/A _6444_/B VGND VGND VPWR VPWR _3305_/Y sky130_fd_sc_hd__nand2_1
X_7073_ _7073_/CLK hold60/X fanout582/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dfrtp_4
X_4285_ _4285_/A _4637_/A VGND VGND VPWR VPWR _4288_/C sky130_fd_sc_hd__nand2_1
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6024_ _6024_/A1 _5761_/X _6023_/X VGND VGND VPWR VPWR _7203_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6926_ _7053_/CLK _6926_/D fanout603/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6857_ _6875_/CLK _6857_/D fanout596/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5808_ _7047_/Q _5815_/C _5814_/C _6072_/C _7015_/Q VGND VGND VPWR VPWR _5808_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6788_ _7150_/CLK _6788_/D fanout602/X VGND VGND VPWR VPWR _7290_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_167_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5739_ _5737_/Y _5738_/X _5759_/B _6141_/B _5712_/Y VGND VGND VPWR VPWR _7187_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_108_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold460 _3971_/X VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold471 _6963_/Q VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _6891_/Q VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold493 _5379_/X VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1160 _4140_/X VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _7239_/Q VGND VGND VPWR VPWR _6519_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 _7285_/A VGND VGND VPWR VPWR _4089_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 _6098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _7293_/A VGND VGND VPWR VPWR _4195_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_311 _6122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_322 _6768_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _7076_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _6782_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 _3313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_366 _6073_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_377 _4053_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 _5723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_399 _6109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4070_ hold24/X _4070_/A1 hold57/X VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__mux2_1
XFILLER_110_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4972_ _4718_/D _4804_/C _4294_/B _4799_/B VGND VGND VPWR VPWR _4973_/C sky130_fd_sc_hd__o211a_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6711_ _7122_/CLK _6711_/D fanout608/X VGND VGND VPWR VPWR _7301_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_51_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3923_ hold13/X _3913_/B _3921_/X _3914_/S hold880/X VGND VGND VPWR VPWR _3923_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6642_ _7248_/CLK _6642_/D fanout580/X VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3854_ _7165_/Q _3509_/X _3559_/X _6909_/Q _3853_/X VGND VGND VPWR VPWR _3854_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ _7096_/CLK _6573_/D fanout596/X VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfrtp_1
X_3785_ _6772_/Q _5304_/A _5494_/C _6536_/D _3784_/X VGND VGND VPWR VPWR _3785_/X
+ sky130_fd_sc_hd__a41o_1
X_5524_ hold672/X _3918_/B _5529_/S VGND VGND VPWR VPWR _5524_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5455_ hold123/X hold83/X _5457_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4406_ _4359_/Y _4372_/Y _4848_/B VGND VGND VPWR VPWR _4878_/B sky130_fd_sc_hd__a21oi_4
X_5386_ _6524_/B _5449_/B _5548_/D _5422_/D VGND VGND VPWR VPWR _5394_/S sky130_fd_sc_hd__and4_4
XFILLER_160_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7125_ _7171_/CLK _7125_/D fanout609/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_4
X_4337_ _4246_/Y _4301_/Y _4327_/Y VGND VGND VPWR VPWR _4509_/C sky130_fd_sc_hd__o21ai_1
X_7056_ _7131_/CLK _7056_/D fanout606/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_87_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4268_ _4632_/A _4511_/A VGND VGND VPWR VPWR _4940_/C sky130_fd_sc_hd__nor2_8
X_6007_ _6754_/Q _6073_/B2 _5774_/X _6669_/Q _6006_/X VGND VGND VPWR VPWR _6007_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4199_ _4199_/A0 _4198_/X _4205_/S VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6957_/CLK _6909_/D fanout591/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold290 _7118_/Q VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _6987_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 _6636_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_152 _6945_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_163 input23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _6072_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_196 _6425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3570_ _7261_/Q _5512_/B _3457_/X _3496_/X _6992_/Q VGND VGND VPWR VPWR _3570_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5240_ _4398_/X _4403_/X _5239_/X _5047_/X VGND VGND VPWR VPWR _5241_/B sky130_fd_sc_hd__o31a_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5171_ _4620_/B _4786_/B _4923_/A _5033_/A _5033_/B VGND VGND VPWR VPWR _5217_/C
+ sky130_fd_sc_hd__a311oi_1
X_4122_ _4152_/B hold941/X _4126_/S VGND VGND VPWR VPWR _4122_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ hold64/X _4053_/B VGND VGND VPWR VPWR _4053_/X sky130_fd_sc_hd__and2_2
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4955_ _4650_/Y _4658_/Y _4745_/Y _4944_/X _4954_/Y VGND VGND VPWR VPWR _4955_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3906_ _3905_/Y _3906_/A1 _3906_/S VGND VGND VPWR VPWR _6586_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4886_ _4859_/C _4862_/A _4729_/D _4708_/A _4788_/A VGND VGND VPWR VPWR _5007_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6625_ _7219_/CLK _6625_/D VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3837_ _6916_/Q _5422_/D _5281_/A2 _3471_/X input25/X VGND VGND VPWR VPWR _3837_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6556_ _7260_/CLK _6556_/D fanout579/X VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfstp_1
X_3768_ _6747_/Q _5311_/B _5273_/D _3767_/X VGND VGND VPWR VPWR _3768_/X sky130_fd_sc_hd__a31o_1
XFILLER_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5507_ _3428_/X _3922_/X _5511_/S hold894/X VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__a22o_1
XFILLER_180_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6487_ _7257_/Q _6487_/A2 _6487_/B1 _7258_/Q VGND VGND VPWR VPWR _6487_/X sky130_fd_sc_hd__a22o_1
X_3699_ _3346_/D _5341_/A hold56/A _3698_/X VGND VGND VPWR VPWR _3699_/X sky130_fd_sc_hd__a31o_2
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5438_ _4051_/B hold450/X hold67/X VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__mux2_1
Xoutput340 hold589/X VGND VGND VPWR VPWR hold590/A sky130_fd_sc_hd__buf_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5369_ _5369_/A0 _5649_/A0 _5376_/S VGND VGND VPWR VPWR _5369_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ _7108_/CLK _7108_/D fanout607/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7039_ _7159_/CLK _7039_/D fanout599/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _5128_/A _4859_/C _4740_/C _4878_/B VGND VGND VPWR VPWR _4740_/Y sky130_fd_sc_hd__nand4_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ _4666_/Y _4376_/Y _4663_/Y _4667_/Y _4670_/Y VGND VGND VPWR VPWR _4672_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_186_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6410_ _7277_/Q _6444_/C _5750_/C _6098_/X _6750_/Q VGND VGND VPWR VPWR _6410_/X
+ sky130_fd_sc_hd__a32o_1
X_3622_ _6830_/Q _5325_/C _5311_/C _7032_/Q _3547_/X VGND VGND VPWR VPWR _3622_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_128_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6341_ _6878_/Q _6134_/Y _3246_/Y VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__o21a_1
X_3553_ _5304_/A _5575_/C _4158_/D VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__and3_2
XFILLER_127_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6272_ _7092_/Q _6106_/X _6107_/X _7004_/Q _6271_/X VGND VGND VPWR VPWR _6290_/B
+ sky130_fd_sc_hd__a221o_1
X_3484_ input61/X _5334_/B _3913_/B _6592_/Q _3483_/X VGND VGND VPWR VPWR _3485_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5223_ _5220_/X _5266_/B _5217_/X VGND VGND VPWR VPWR _5243_/A sky130_fd_sc_hd__a21bo_1
XFILLER_142_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5154_ _5153_/X _4271_/Y _5248_/A3 _4648_/Y VGND VGND VPWR VPWR _5204_/B sky130_fd_sc_hd__a211o_1
X_4105_ _6538_/A0 hold371/X _4108_/S VGND VGND VPWR VPWR _4105_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5085_ _4804_/A _5036_/C _5128_/C wire442/X VGND VGND VPWR VPWR _5085_/X sky130_fd_sc_hd__a31o_1
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4036_ _6543_/A0 hold837/X _4040_/S VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5987_ _6658_/Q _5794_/X _5983_/X _5985_/X _5986_/X VGND VGND VPWR VPWR _5987_/X
+ sky130_fd_sc_hd__a2111o_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _4945_/B _4712_/B _4747_/Y _4791_/X VGND VGND VPWR VPWR _4938_/X sky130_fd_sc_hd__a31o_1
XANTENNA_30 _3466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4859_/C _5255_/A _4683_/X _4641_/B _4718_/D VGND VGND VPWR VPWR _4872_/C
+ sky130_fd_sc_hd__a32o_1
XANTENNA_41 _3496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _5593_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _3918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6608_ _7248_/CLK _6608_/D fanout580/X VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_74 _5750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _5782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _6129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6539_ _6539_/A0 _6539_/A1 _6541_/S VGND VGND VPWR VPWR _6539_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput181 _3270_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3260_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5910_ _7004_/Q _5795_/D _5795_/C VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__o21a_1
X_6890_ _7143_/CLK _6890_/D fanout589/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ _6961_/Q wire398/X _5934_/C _7049_/Q _5814_/X VGND VGND VPWR VPWR _5841_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5772_ _7183_/Q _7182_/Q VGND VGND VPWR VPWR _5814_/C sky130_fd_sc_hd__and2b_4
X_4723_ _4723_/A _4723_/B _4723_/C VGND VGND VPWR VPWR _4723_/Y sky130_fd_sc_hd__nor3_1
X_4654_ _4848_/B _4654_/B _4691_/B _4662_/B VGND VGND VPWR VPWR _4982_/D sky130_fd_sc_hd__and4_2
XFILLER_135_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
X_3605_ _6856_/Q _5327_/D _3902_/A3 _4121_/B _6749_/Q VGND VGND VPWR VPWR _3605_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_2
Xhold801 _3998_/X VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_1
X_4585_ _4585_/A _4585_/B _4925_/C VGND VGND VPWR VPWR _4587_/B sky130_fd_sc_hd__nand3_1
XFILLER_162_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold812 _7020_/Q VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold823 _3938_/X VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_2
Xinput94 uart_enabled VGND VGND VPWR VPWR _3349_/A sky130_fd_sc_hd__clkbuf_2
X_6324_ _7126_/Q _6176_/B _6425_/B _6143_/X _6950_/Q VGND VGND VPWR VPWR _6324_/X
+ sky130_fd_sc_hd__a32o_1
Xhold834 _5626_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3536_ _5476_/B _5476_/C _5494_/C VGND VGND VPWR VPWR _3536_/X sky130_fd_sc_hd__and3_4
Xhold845 _5338_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap564 _4799_/A VGND VGND VPWR VPWR _4294_/B sky130_fd_sc_hd__clkbuf_2
Xhold856 _7044_/Q VGND VGND VPWR VPWR hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _6543_/X VGND VGND VPWR VPWR _7270_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _6656_/Q VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 _5631_/X VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ _6255_/A _6255_/B _6255_/C _6255_/D VGND VGND VPWR VPWR _6255_/Y sky130_fd_sc_hd__nor4_1
X_3467_ _7275_/Q _5630_/A _3466_/X _4204_/S input43/X VGND VGND VPWR VPWR _3467_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_131_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5206_ _4423_/Y _4633_/Y _4638_/Y _5082_/A VGND VGND VPWR VPWR _5246_/C sky130_fd_sc_hd__o31a_1
XFILLER_131_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6186_ _6920_/Q _6129_/B _6454_/B1 _6952_/Q VGND VGND VPWR VPWR _6186_/X sky130_fd_sc_hd__a22o_1
X_3398_ _6549_/A0 _3398_/A1 _3402_/S VGND VGND VPWR VPWR _3398_/X sky130_fd_sc_hd__mux2_1
Xhold1501 _5372_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 _6832_/Q VGND VGND VPWR VPWR hold116/A sky130_fd_sc_hd__dlygate4sd3_1
X_5137_ _4380_/X _5040_/X _4403_/X _4820_/X _5136_/X VGND VGND VPWR VPWR _5261_/C
+ sky130_fd_sc_hd__o311a_1
Xhold1523 _6984_/Q VGND VGND VPWR VPWR hold342/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _7198_/Q VGND VGND VPWR VPWR _5909_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1545 _5977_/X VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_184_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5068_ _4689_/C _4945_/B _4945_/C _4942_/X VGND VGND VPWR VPWR _5068_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4019_ _4017_/B _3916_/X _4021_/S hold946/X VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold108 _6853_/Q VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold119 _6828_/Q VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ _4689_/B _4761_/C _4209_/Y _4369_/X VGND VGND VPWR VPWR _4848_/B sky130_fd_sc_hd__o31a_2
XFILLER_172_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3321_ _4168_/B _3321_/B VGND VGND VPWR VPWR _7249_/D sky130_fd_sc_hd__nand2b_1
XFILLER_171_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6599_/Q _6025_/B _6028_/B _5789_/X _6780_/Q VGND VGND VPWR VPWR _6040_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _7138_/Q VGND VGND VPWR VPWR _3252_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6942_ _7160_/CLK _6942_/D fanout592/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6873_ _7274_/CLK _6873_/D fanout577/X VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ _6960_/Q _5770_/X _5793_/X _6984_/Q _5823_/X VGND VGND VPWR VPWR _5824_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_139_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5755_ _5759_/A _3307_/B _5758_/S VGND VGND VPWR VPWR _5755_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_90_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7239_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4706_ _4848_/A _4706_/B _4730_/A VGND VGND VPWR VPWR _4792_/C sky130_fd_sc_hd__and3_4
XFILLER_30_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5686_ hold275/X _3915_/B _5692_/S VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4637_ _4637_/A _4747_/A _4747_/B _4747_/C VGND VGND VPWR VPWR _4637_/Y sky130_fd_sc_hd__nor4_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold620 _4071_/X VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold631 _7162_/Q VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _4815_/A _4923_/A _4606_/D _4589_/C VGND VGND VPWR VPWR _4570_/A sky130_fd_sc_hd__and4_1
XFILLER_116_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold642 _5642_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _6693_/Q VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3519_ _6536_/C _6530_/C _4127_/C VGND VGND VPWR VPWR _3927_/B sky130_fd_sc_hd__and3_2
Xhold664 _7242_/Q VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlygate4sd3_1
X_6307_ _6981_/Q _6452_/B1 _6143_/X _6949_/Q _6306_/X VGND VGND VPWR VPWR _6314_/A
+ sky130_fd_sc_hd__a221o_1
Xhold675 _5474_/X VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7287_ _7287_/A VGND VGND VPWR VPWR _7287_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap383 _4984_/B VGND VGND VPWR VPWR _4859_/A sky130_fd_sc_hd__buf_4
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold686 hold686/A VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap394 _5789_/X VGND VGND VPWR VPWR _5970_/B1 sky130_fd_sc_hd__buf_12
X_4499_ _4632_/A _4511_/A _4632_/C VGND VGND VPWR VPWR _4792_/B sky130_fd_sc_hd__nor3_4
Xhold697 _5402_/X VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6238_ _7018_/Q _6177_/X _6235_/X _6237_/X VGND VGND VPWR VPWR _6239_/C sky130_fd_sc_hd__a211o_1
XFILLER_103_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _7168_/Q _6117_/X _6323_/B1 _6960_/Q _6168_/X VGND VGND VPWR VPWR _6169_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _6670_/Q VGND VGND VPWR VPWR hold945/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1331 _5560_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1342 _6742_/Q VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1353 _7024_/Q VGND VGND VPWR VPWR hold802/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 _7151_/Q VGND VGND VPWR VPWR hold1364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 _7267_/Q VGND VGND VPWR VPWR hold1375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1386 _6834_/Q VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1397 _5604_/X VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7174_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7088_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3870_ _6739_/Q _3441_/X _3525_/X _7125_/Q _3869_/X VGND VGND VPWR VPWR _3873_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ _6549_/A0 _5540_/A1 hold77/X VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5471_ _3921_/B hold550/X _5475_/S VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7210_ _7259_/CLK _7210_/D fanout595/X VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfrtp_1
X_4422_ _4698_/A _4657_/C _4656_/C _4647_/C VGND VGND VPWR VPWR _4422_/Y sky130_fd_sc_hd__nor4_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7141_ _7148_/CLK _7141_/D fanout592/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_2
X_4353_ _4632_/A _4511_/A _4633_/B VGND VGND VPWR VPWR _4859_/C sky130_fd_sc_hd__and3_4
Xfanout407 _3457_/X VGND VGND VPWR VPWR _5325_/C sky130_fd_sc_hd__buf_12
Xfanout418 _6347_/C VGND VGND VPWR VPWR _6143_/C sky130_fd_sc_hd__clkbuf_16
X_3304_ _7188_/Q _7189_/Q _7190_/Q _7187_/Q VGND VGND VPWR VPWR _6444_/B sky130_fd_sc_hd__and4bb_4
X_7072_ _7072_/CLK _7072_/D fanout599/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_98_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout429 _5720_/Y VGND VGND VPWR VPWR _5815_/B sky130_fd_sc_hd__buf_6
X_4284_ _4284_/A _4284_/B _4284_/C _4310_/B VGND VGND VPWR VPWR _4667_/C sky130_fd_sc_hd__nand4_4
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6023_ _6442_/S _6023_/A2 _6443_/S _6022_/X VGND VGND VPWR VPWR _6023_/X sky130_fd_sc_hd__a211o_1
XFILLER_67_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6957_/CLK _6925_/D fanout591/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6856_ _7244_/CLK _6856_/D fanout581/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_1
X_5807_ _6895_/Q _5795_/X _5805_/X _5806_/X _5790_/X VGND VGND VPWR VPWR _5807_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3999_ _5304_/A _5476_/B _6536_/B _4158_/D VGND VGND VPWR VPWR _4003_/S sky130_fd_sc_hd__nand4_4
X_6787_ _7053_/CLK _6787_/D fanout601/X VGND VGND VPWR VPWR _7289_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5738_ _7186_/Q _7185_/Q _6141_/B VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5669_ _5674_/S hold923/X _3550_/X _3919_/X VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold450 _6949_/Q VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold461 _6621_/Q VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold472 _5454_/X VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _5373_/X VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _6696_/Q VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1150 _6549_/X VGND VGND VPWR VPWR _7275_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1161 _7111_/Q VGND VGND VPWR VPWR _5621_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1172 _6519_/X VGND VGND VPWR VPWR _7239_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1183 _4089_/X VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 _6129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _4195_/X VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_312 _6129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _6962_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 _7261_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_345 _6779_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_356 _3313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _6176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_378 _6444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_389 _5723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4971_ _4729_/A _4480_/B _4792_/B _4970_/X VGND VGND VPWR VPWR _4973_/B sky130_fd_sc_hd__a31o_1
XFILLER_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6710_ _7117_/CLK _6710_/D fanout608/X VGND VGND VPWR VPWR _7300_/A sky130_fd_sc_hd__dfrtp_1
X_3922_ _5494_/A hold64/X _3922_/C VGND VGND VPWR VPWR _3922_/X sky130_fd_sc_hd__and3_4
XFILLER_189_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3853_ _7037_/Q _3547_/X _5593_/B _7093_/Q VGND VGND VPWR VPWR _3853_/X sky130_fd_sc_hd__a22o_1
X_6641_ _7275_/CLK _6641_/D fanout596/X VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3784_ _6822_/Q _3434_/X _3564_/X _7269_/Q _3783_/X VGND VGND VPWR VPWR _3784_/X
+ sky130_fd_sc_hd__a221o_1
X_6572_ _6650_/CLK _6572_/D fanout596/X VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5523_ hold802/X _3915_/B _5529_/S VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5454_ hold471/X _3925_/C _5457_/S VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4405_ _5042_/A _5042_/B _4519_/C VGND VGND VPWR VPWR _4878_/A sky130_fd_sc_hd__and3_2
X_5385_ hold194/X _4053_/B _5385_/S VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4336_ _4208_/Y _4246_/Y _4940_/C _4327_/Y VGND VGND VPWR VPWR _4336_/X sky130_fd_sc_hd__o31a_1
X_7124_ _7132_/CLK _7124_/D fanout610/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_2
X_7055_ _7087_/CLK _7055_/D fanout589/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4267_ _5036_/B _4632_/C _4729_/A VGND VGND VPWR VPWR _4689_/C sky130_fd_sc_hd__and3_2
X_6006_ _6664_/Q _5934_/C _6028_/B _6003_/X _6005_/X VGND VGND VPWR VPWR _6006_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4198_ hold571/X _3924_/X _4204_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6908_ _6908_/CLK _6908_/D fanout609/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6839_ _7071_/CLK _6839_/D fanout585/X VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold280 _6913_/Q VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold291 _5628_/X VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _6489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _6643_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _6773_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _3351_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _7312_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _6072_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _6446_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5170_ _4786_/B _4620_/C _5089_/A VGND VGND VPWR VPWR _5172_/C sky130_fd_sc_hd__o21ai_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4121_ _6542_/A _4121_/B VGND VGND VPWR VPWR _4126_/S sky130_fd_sc_hd__nand2_4
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4052_ hold136/X hold21/X _4054_/S VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4954_ _4954_/A _4954_/B _4954_/C _4954_/D VGND VGND VPWR VPWR _4954_/Y sky130_fd_sc_hd__nor4_1
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3905_ _3905_/A _3905_/B _3905_/C VGND VGND VPWR VPWR _3905_/Y sky130_fd_sc_hd__nand3_4
XFILLER_177_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4885_ _4862_/A _5128_/B _4729_/D _4717_/A VGND VGND VPWR VPWR _5228_/A sky130_fd_sc_hd__a31oi_1
XFILLER_177_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6624_ _7269_/CLK _6624_/D fanout580/X VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3836_ _7068_/Q _5566_/B _4092_/S _3349_/B _3835_/X VGND VGND VPWR VPWR _3843_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6555_ _7274_/CLK hold99/X fanout577/X VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfrtp_2
X_3767_ _6777_/Q _3542_/B _3457_/X _3548_/X _7051_/Q VGND VGND VPWR VPWR _3767_/X
+ sky130_fd_sc_hd__a32o_1
X_5506_ _3428_/X _3919_/X _5511_/S _5506_/B2 VGND VGND VPWR VPWR _5506_/X sky130_fd_sc_hd__a22o_1
X_3698_ _6636_/Q _3969_/C _4187_/S input38/X _3697_/X VGND VGND VPWR VPWR _3698_/X
+ sky130_fd_sc_hd__a221o_1
X_6486_ _6485_/X _6486_/B _6486_/C VGND VGND VPWR VPWR _6511_/S sky130_fd_sc_hd__nand3b_4
XFILLER_105_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5437_ hold83/X hold149/X hold67/X VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__mux2_1
Xoutput330 hold597/X VGND VGND VPWR VPWR hold598/A sky130_fd_sc_hd__buf_12
Xoutput341 hold617/X VGND VGND VPWR VPWR hold618/A sky130_fd_sc_hd__buf_12
X_5368_ _6524_/B _5476_/C _5575_/C _5422_/D VGND VGND VPWR VPWR _5376_/S sky130_fd_sc_hd__and4_4
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7107_ _7108_/CLK _7107_/D fanout607/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4319_ _4312_/A _4544_/D _4637_/A _4214_/A VGND VGND VPWR VPWR _4319_/X sky130_fd_sc_hd__a211o_1
X_5299_ _3922_/C hold116/X hold73/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7038_ _7156_/CLK _7038_/D fanout602/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire402 _5476_/Y VGND VGND VPWR VPWR _5484_/S sky130_fd_sc_hd__buf_6
XFILLER_128_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout590 fanout593/X VGND VGND VPWR VPWR fanout590/X sky130_fd_sc_hd__buf_8
XFILLER_76_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4670_ _4984_/A _4859_/A _4732_/C _4670_/D VGND VGND VPWR VPWR _4670_/Y sky130_fd_sc_hd__nand4_1
XFILLER_187_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3621_ _6674_/Q _3533_/C _4139_/C _3434_/X _6819_/Q VGND VGND VPWR VPWR _3621_/X
+ sky130_fd_sc_hd__a32o_1
X_3552_ _7151_/Q _3550_/X _5593_/B _7087_/Q _3549_/X VGND VGND VPWR VPWR _3561_/C
+ sky130_fd_sc_hd__a221o_2
X_6340_ _6321_/X _6340_/B _6340_/C VGND VGND VPWR VPWR _6340_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_143_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6271_ _7012_/Q _6444_/C _6328_/A3 _6098_/X _6988_/Q VGND VGND VPWR VPWR _6271_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3483_ _6688_/Q _5341_/A _5327_/D _3482_/X _6768_/Q VGND VGND VPWR VPWR _3483_/X
+ sky130_fd_sc_hd__a32o_2
X_5222_ _4556_/A _5094_/B _5222_/C _5222_/D VGND VGND VPWR VPWR _5266_/B sky130_fd_sc_hd__and4bb_1
X_5153_ _4689_/B _4255_/A _4208_/Y _4496_/Y VGND VGND VPWR VPWR _5153_/X sky130_fd_sc_hd__o31a_2
X_4104_ _4152_/B _4104_/A1 _4108_/S VGND VGND VPWR VPWR _4104_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5084_ _5128_/A _4788_/A _4718_/D _5083_/X VGND VGND VPWR VPWR _5084_/X sky130_fd_sc_hd__a31o_1
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4035_ _6524_/A _6524_/B _6530_/D _5327_/D VGND VGND VPWR VPWR _4040_/S sky130_fd_sc_hd__nand4_4
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5986_ _6587_/Q _5814_/X _5815_/X _6638_/Q _5978_/X VGND VGND VPWR VPWR _5986_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4937_ _4620_/A _5128_/C _5263_/B _5036_/A _5140_/C VGND VGND VPWR VPWR _4976_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_178_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_20 _3428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _3466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4868_ _4853_/C _4945_/C _4756_/C _4683_/X _4878_/A VGND VGND VPWR VPWR _4872_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA_42 _3499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _3918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _7265_/CLK _6607_/D fanout575/X VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_2
X_3819_ _6834_/Q _5325_/C _5311_/C _7148_/Q _3474_/X VGND VGND VPWR VPWR _3819_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA_75 _5764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _5782_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4799_/A _4799_/B _4799_/C VGND VGND VPWR VPWR _4799_/X sky130_fd_sc_hd__and3_1
XANTENNA_97 _6129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6538_ _6538_/A0 hold431/X _6541_/S VGND VGND VPWR VPWR _6538_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6469_ _7253_/Q _7256_/Q VGND VGND VPWR VPWR _6469_/Y sky130_fd_sc_hd__nor2_1
Xoutput171 _3351_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
Xoutput182 _3269_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3259_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5840_ _5861_/A2 _5761_/X _5839_/X _5838_/X VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__o22a_1
XFILLER_62_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5771_ _7183_/Q _7182_/Q _6010_/C _5795_/D VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__and4_4
XFILLER_15_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4722_ _4722_/A _4984_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _4722_/Y sky130_fd_sc_hd__nand4_2
XFILLER_187_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4653_ _5255_/A _4653_/B _4755_/B _4860_/B VGND VGND VPWR VPWR _4672_/C sky130_fd_sc_hd__nand4_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
X_3604_ _6684_/Q _4029_/B _3558_/X _6608_/Q VGND VGND VPWR VPWR _3604_/X sky130_fd_sc_hd__a22o_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_2
Xhold802 hold802/A VGND VGND VPWR VPWR hold802/X sky130_fd_sc_hd__dlygate4sd3_1
X_4584_ _4751_/A _4584_/B _5263_/A _4589_/C VGND VGND VPWR VPWR _4925_/C sky130_fd_sc_hd__nand4_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _7314_/A sky130_fd_sc_hd__clkbuf_2
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR _7308_/A sky130_fd_sc_hd__clkbuf_2
Xhold813 _5518_/X VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold824 _7127_/Q VGND VGND VPWR VPWR hold824/X sky130_fd_sc_hd__dlygate4sd3_1
X_6323_ _6990_/Q _6098_/X _6323_/B1 _6966_/Q _6322_/X VGND VGND VPWR VPWR _6330_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3535_ _6753_/Q _3531_/X _3534_/X _3530_/X _3529_/X VGND VGND VPWR VPWR _3561_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold835 _7068_/Q VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _6938_/Q VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap554 _4600_/Y VGND VGND VPWR VPWR _4620_/C sky130_fd_sc_hd__clkbuf_2
Xhold857 _5545_/X VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold868 _7036_/Q VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 _3997_/X VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ _6987_/Q _6098_/X _6115_/X _7139_/Q _6253_/X VGND VGND VPWR VPWR _6255_/D
+ sky130_fd_sc_hd__a221o_1
X_3466_ _5324_/B _6804_/Q _6805_/Q _6548_/D VGND VGND VPWR VPWR _3466_/X sky130_fd_sc_hd__and4_4
XFILLER_143_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5205_ _5153_/X _4701_/Y _4961_/X _5159_/C _5076_/C VGND VGND VPWR VPWR _5249_/B
+ sky130_fd_sc_hd__o2111a_1
X_6185_ _7160_/Q _6104_/X _6130_/X _6928_/Q _6184_/X VGND VGND VPWR VPWR _6190_/B
+ sky130_fd_sc_hd__a221o_1
X_3397_ _6548_/B _3397_/B VGND VGND VPWR VPWR _3402_/S sky130_fd_sc_hd__nand2_4
Xhold1502 _7205_/Q VGND VGND VPWR VPWR _6090_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _7199_/Q VGND VGND VPWR VPWR _5954_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5136_ _4391_/Y _4490_/Y _4348_/X _4356_/Y _4382_/Y VGND VGND VPWR VPWR _5136_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1524 _7207_/Q VGND VGND VPWR VPWR _6167_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _7206_/Q VGND VGND VPWR VPWR _6091_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1546 _7225_/Q VGND VGND VPWR VPWR _6477_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5067_ _5263_/B _4748_/B _4945_/C _4903_/B VGND VGND VPWR VPWR _5067_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4018_ _4152_/B hold929/X _4021_/S VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5969_ _6974_/Q _5771_/X _5956_/X _5958_/X _5968_/X VGND VGND VPWR VPWR _5969_/Y
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_40_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 _5329_/X VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3320_ _3354_/B _7249_/Q VGND VGND VPWR VPWR _3321_/B sky130_fd_sc_hd__nand2b_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _7146_/Q VGND VGND VPWR VPWR _3251_/Y sky130_fd_sc_hd__inv_2
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6941_ _7143_/CLK _6941_/D fanout588/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfrtp_4
X_6872_ _7099_/CLK _6872_/D fanout598/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5823_ _6976_/Q _6073_/B2 _5774_/X _6904_/Q _5822_/X VGND VGND VPWR VPWR _5823_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5754_ _6803_/Q _6442_/S _6800_/Q _5759_/B _5753_/X VGND VGND VPWR VPWR _5758_/S
+ sky130_fd_sc_hd__o41a_1
XFILLER_175_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4705_ _4705_/A _4705_/B _4705_/C VGND VGND VPWR VPWR _4711_/A sky130_fd_sc_hd__nor3_1
XFILLER_147_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5685_ _5685_/A0 _6549_/A0 _5692_/S VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4636_ _4637_/A _4747_/A VGND VGND VPWR VPWR _4940_/D sky130_fd_sc_hd__nor2_1
Xhold610 _3400_/X VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 hold621/A VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlygate4sd3_1
X_4567_ _4320_/A _4523_/C _4322_/Y _4870_/B VGND VGND VPWR VPWR _4567_/Y sky130_fd_sc_hd__o211ai_4
Xhold632 _5679_/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold643 hold643/A VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 _4043_/Y VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _7061_/Q _6136_/A _6465_/A3 _6145_/X _7013_/Q VGND VGND VPWR VPWR _6306_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3518_ _4127_/C _5422_/D _5575_/D VGND VGND VPWR VPWR _5377_/C sky130_fd_sc_hd__and3_4
Xhold665 _6522_/X VGND VGND VPWR VPWR _7242_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap373 _6134_/Y VGND VGND VPWR VPWR _6466_/A1 sky130_fd_sc_hd__buf_8
X_7286_ _7286_/A VGND VGND VPWR VPWR _7286_/X sky130_fd_sc_hd__clkbuf_2
Xmax_cap384 _6142_/X VGND VGND VPWR VPWR _6454_/B1 sky130_fd_sc_hd__buf_12
Xhold676 hold676/A VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _5060_/A _5060_/B _5143_/D _4718_/D VGND VGND VPWR VPWR _4504_/B sky130_fd_sc_hd__nand4_1
Xhold687 hold687/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
Xmax_cap395 _5781_/X VGND VGND VPWR VPWR _6072_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold698 _7027_/Q VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6237_ _7114_/Q _6110_/X _6137_/X _7098_/Q _6236_/X VGND VGND VPWR VPWR _6237_/X
+ sky130_fd_sc_hd__a221o_1
X_3449_ _3351_/B _4092_/S _3445_/X _6887_/Q _3448_/X VGND VGND VPWR VPWR _3462_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _7032_/Q _6465_/A2 _6465_/A3 _6325_/A2 _6880_/Q VGND VGND VPWR VPWR _6168_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _4002_/X VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _4014_/X VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1332 _6970_/Q VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _4114_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5119_ _4939_/A _4738_/B _4411_/B _4984_/B _4984_/C VGND VGND VPWR VPWR _5120_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_182_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1354 _5523_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6099_ _6967_/Q _6097_/X _6098_/X _6983_/Q VGND VGND VPWR VPWR _6099_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1365 _5667_/X VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1376 _6539_/X VGND VGND VPWR VPWR _7267_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1387 _6806_/Q VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _6578_/Q VGND VGND VPWR VPWR hold786/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5470_ _3918_/B hold318/X _5475_/S VGND VGND VPWR VPWR _5470_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4421_ _4656_/C _4647_/C VGND VGND VPWR VPWR _4699_/B sky130_fd_sc_hd__nor2_2
XFILLER_172_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7140_ _7140_/CLK _7140_/D fanout609/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_1
X_4352_ _4632_/C _4612_/C VGND VGND VPWR VPWR _4633_/B sky130_fd_sc_hd__nor2_8
XFILLER_153_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout408 _5684_/C VGND VGND VPWR VPWR _5281_/A2 sky130_fd_sc_hd__buf_12
X_3303_ _7188_/Q _6141_/B VGND VGND VPWR VPWR _6138_/A sky130_fd_sc_hd__and2b_4
X_7071_ _7071_/CLK _7071_/D fanout585/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfstp_1
Xfanout419 _6092_/Y VGND VGND VPWR VPWR _6347_/C sky130_fd_sc_hd__buf_12
X_4283_ _4235_/A _4282_/Y _4285_/A _4747_/A VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__a2bb2oi_4
X_6022_ _6689_/Q _5726_/Y _6008_/X _6021_/X _5759_/A VGND VGND VPWR VPWR _6022_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ _7148_/CLK _6924_/D fanout591/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _6855_/CLK _6855_/D fanout584/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5806_ _7039_/Q _6072_/B _6028_/B _5793_/X _6983_/Q VGND VGND VPWR VPWR _5806_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6786_ _7006_/CLK _6786_/D fanout601/X VGND VGND VPWR VPWR _7288_/A sky130_fd_sc_hd__dfrtp_1
X_3998_ _3994_/S hold800/X _3502_/X _3925_/X VGND VGND VPWR VPWR _3998_/X sky130_fd_sc_hd__a22o_1
X_5737_ _6141_/B _6136_/A VGND VGND VPWR VPWR _5737_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5668_ _5674_/S hold798/X _3550_/X _3916_/X VGND VGND VPWR VPWR _5668_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4619_ _4620_/A _5128_/C _5263_/B _5036_/A _4859_/C VGND VGND VPWR VPWR _4619_/X
+ sky130_fd_sc_hd__a32o_1
X_5599_ _4049_/B hold367/X hold14/X VGND VGND VPWR VPWR _5599_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold440 _6749_/Q VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold451 _5438_/X VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold462 _3956_/X VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold473 _6907_/Q VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold484 _7113_/Q VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold495 _4047_/X VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7269_ _7269_/CLK _7269_/D fanout580/X VGND VGND VPWR VPWR _7269_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_49_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1140 _6842_/Q VGND VGND VPWR VPWR _5312_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1151 _6753_/Q VGND VGND VPWR VPWR _4128_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _5621_/X VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1173 _6574_/Q VGND VGND VPWR VPWR _3398_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _6993_/Q VGND VGND VPWR VPWR _5488_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1195 _6851_/Q VGND VGND VPWR VPWR _5326_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_302 _6109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_313 _6129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 _6756_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 _7083_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _6776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_357 _6739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_368 _6425_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 _6444_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4970_ _4970_/A _4970_/B _5089_/C _4970_/D VGND VGND VPWR VPWR _4970_/X sky130_fd_sc_hd__and4_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3921_ hold65/X _3921_/B VGND VGND VPWR VPWR _3921_/X sky130_fd_sc_hd__and2_4
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6640_ _7263_/CLK _6640_/D fanout577/X VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfstp_2
X_3852_ _7101_/Q _3510_/X _3515_/X _7029_/Q VGND VGND VPWR VPWR _3852_/X sky130_fd_sc_hd__a22o_1
X_6571_ _7275_/CLK _6571_/D fanout596/X VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfstp_1
X_3783_ _6573_/Q _6548_/A _5341_/A _3525_/X _7123_/Q VGND VGND VPWR VPWR _3783_/X
+ sky130_fd_sc_hd__a32o_2
X_5522_ _5522_/A0 _6549_/A0 _5529_/S VGND VGND VPWR VPWR _5522_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5453_ hold232/X _3922_/C _5457_/S VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4404_ _4427_/C _4429_/D _4388_/Y _4383_/A _4380_/X VGND VGND VPWR VPWR _4444_/C
+ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_42_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7168_/CLK sky130_fd_sc_hd__clkbuf_16
X_5384_ hold702/X _4051_/B _5385_/S VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7123_ _7123_/CLK _7123_/D fanout607/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_4
X_4335_ _4356_/A _4848_/A _4295_/A VGND VGND VPWR VPWR _4484_/C sky130_fd_sc_hd__a21oi_1
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7054_ _7163_/CLK _7054_/D fanout610/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4266_ _5040_/C _4244_/Y _4265_/Y _7257_/Q VGND VGND VPWR VPWR _4266_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_140_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6005_ _6684_/Q _5768_/X _5794_/X _6659_/Q VGND VGND VPWR VPWR _6005_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_57_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7035_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4197_ _4197_/A0 _4196_/X _4205_/S VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _7015_/CLK _6907_/D fanout588/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6838_ _7073_/CLK _6838_/D fanout585/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6769_ _7007_/CLK _6769_/D fanout590/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold270 _7064_/Q VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _5398_/X VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold292/A VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_110 _6136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_121 _6492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _6621_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _6577_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _6773_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _3353_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_176 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 _6072_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _6446_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4120_ _3925_/C hold448/X _4120_/S VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4051_ hold65/X _4051_/B VGND VGND VPWR VPWR _4051_/X sky130_fd_sc_hd__and2_4
XFILLER_37_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4953_ _4923_/B _4945_/C _4659_/B _4945_/X VGND VGND VPWR VPWR _4954_/C sky130_fd_sc_hd__a31o_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3904_ _3904_/A _3904_/B _3904_/C _3904_/D VGND VGND VPWR VPWR _3905_/C sky130_fd_sc_hd__nor4_4
X_4884_ _4884_/A _4884_/B _5002_/A VGND VGND VPWR VPWR _4888_/A sky130_fd_sc_hd__nor3_1
X_6623_ _7260_/CLK _6623_/D fanout579/X VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfrtp_4
X_3835_ _6940_/Q hold39/A _3533_/C _3452_/X _6964_/Q VGND VGND VPWR VPWR _3835_/X
+ sky130_fd_sc_hd__a32o_1
X_6554_ _6751_/CLK _6554_/D _3291_/A VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3766_ _3766_/A _3766_/B _3766_/C _3766_/D VGND VGND VPWR VPWR _3811_/A sky130_fd_sc_hd__nor4_1
XFILLER_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5505_ _6550_/A0 hold292/X _5511_/S VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6485_ _7258_/Q _6482_/Y _6483_/Y _7257_/Q _4165_/Y VGND VGND VPWR VPWR _6485_/X
+ sky130_fd_sc_hd__a221o_1
X_3697_ _6890_/Q _5440_/C _5422_/D _3553_/X _6681_/Q VGND VGND VPWR VPWR _3697_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5436_ _3925_/C hold394/X hold67/X VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__mux2_1
Xoutput320 hold579/X VGND VGND VPWR VPWR hold580/A sky130_fd_sc_hd__buf_12
XFILLER_145_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput331 hold649/X VGND VGND VPWR VPWR hold650/A sky130_fd_sc_hd__buf_12
Xoutput342 hold621/X VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__buf_12
X_5367_ _6511_/A1 hold305/X _5367_/S VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7106_ _7114_/CLK _7106_/D fanout605/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4318_ _4318_/A _4318_/B _4760_/C VGND VGND VPWR VPWR _4620_/A sky130_fd_sc_hd__and3_4
X_5298_ _3919_/C hold277/X hold73/X VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7037_ _7037_/CLK _7037_/D fanout591/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4249_ _4209_/Y _4246_/Y _4662_/B VGND VGND VPWR VPWR _4249_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire447 _3427_/Y VGND VGND VPWR VPWR wire447/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout580 fanout581/X VGND VGND VPWR VPWR fanout580/X sky130_fd_sc_hd__buf_8
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout591 fanout592/X VGND VGND VPWR VPWR fanout591/X sky130_fd_sc_hd__buf_8
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3620_ _7240_/Q _6548_/A _3457_/X _3615_/X _3619_/X VGND VGND VPWR VPWR _3631_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_128_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3551_ _6536_/A _6548_/D hold28/A VGND VGND VPWR VPWR _5593_/B sky130_fd_sc_hd__and3_4
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6270_ _7036_/Q _6138_/B _6108_/X _6109_/X _7044_/Q VGND VGND VPWR VPWR _6270_/X
+ sky130_fd_sc_hd__a32o_1
X_3482_ _6524_/A _5273_/D _6536_/D VGND VGND VPWR VPWR _3482_/X sky130_fd_sc_hd__and3_2
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5221_ _4522_/Y _4613_/Y _4663_/Y _4903_/Y _5020_/D VGND VGND VPWR VPWR _5222_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_142_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5152_ _4945_/C _5151_/Y _4945_/X _5068_/X VGND VGND VPWR VPWR _5152_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4103_ _6524_/A _6536_/B _6530_/D _5279_/D VGND VGND VPWR VPWR _4108_/S sky130_fd_sc_hd__nand4_4
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5083_ _4970_/D _5089_/C _4970_/B _5082_/Y VGND VGND VPWR VPWR _5083_/X sky130_fd_sc_hd__a31o_1
XFILLER_110_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4034_ _6535_/A0 _4034_/A1 _4034_/S VGND VGND VPWR VPWR _4034_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5985_ _6668_/Q _6028_/C _6003_/C _5984_/X VGND VGND VPWR VPWR _5985_/X sky130_fd_sc_hd__a31o_1
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4936_ _5060_/A _4615_/C _4484_/D _4615_/X VGND VGND VPWR VPWR _4976_/B sky130_fd_sc_hd__a31o_1
XANTENNA_10 _3370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _3428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _5120_/A _4867_/B _4867_/C VGND VGND VPWR VPWR _4872_/A sky130_fd_sc_hd__nand3_1
XANTENNA_32 _3466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_43 _3499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _6945_/CLK _6606_/D fanout583/X VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_54 _3609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3818_ _7317_/A _5334_/B _3544_/X _6948_/Q _3817_/X VGND VGND VPWR VPWR _3825_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _5260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _5842_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4632_/A _4209_/Y _4293_/Y _4797_/X VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__o31a_1
XANTENNA_87 _6025_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 _6103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6537_ _4152_/B _6537_/A1 _6541_/S VGND VGND VPWR VPWR _6537_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3749_ _6605_/Q _5666_/C _4139_/C _4152_/C _6776_/Q VGND VGND VPWR VPWR _3749_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6468_ _6468_/A1 _5761_/X _6467_/X VGND VGND VPWR VPWR _7219_/D sky130_fd_sc_hd__o21a_1
XFILLER_161_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5419_ _6505_/A1 hold718/X _5421_/S VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__mux2_1
X_6399_ _7272_/Q _6138_/B _5750_/C _6113_/X _6635_/Q VGND VGND VPWR VPWR _6399_/X
+ sky130_fd_sc_hd__a32o_1
Xoutput172 _7281_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
XFILLER_121_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput183 _3268_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3258_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_99_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _7181_/Q _7180_/Q _6010_/D _5795_/D VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__and4_4
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4859_/A _4984_/C _4721_/C VGND VGND VPWR VPWR _4723_/B sky130_fd_sc_hd__and3_1
XFILLER_147_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4652_ _5255_/A _4653_/B _4860_/B VGND VGND VPWR VPWR _4708_/A sky130_fd_sc_hd__and3_2
XFILLER_30_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3603_ _6565_/Q _3368_/X _5512_/B _3470_/X _7245_/Q VGND VGND VPWR VPWR _3603_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__buf_2
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4583_ _4584_/B _4597_/C _4923_/A _4589_/C VGND VGND VPWR VPWR _4585_/B sky130_fd_sc_hd__nand4_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _3350_/B sky130_fd_sc_hd__clkbuf_4
Xhold803 _6996_/Q VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _7315_/A sky130_fd_sc_hd__clkbuf_2
X_6322_ _7006_/Q _6138_/B _6328_/A3 _6145_/X _7014_/Q VGND VGND VPWR VPWR _6322_/X
+ sky130_fd_sc_hd__a32o_1
Xhold814 _6933_/Q VGND VGND VPWR VPWR hold814/X sky130_fd_sc_hd__dlygate4sd3_1
X_3534_ _6919_/Q _3540_/B _5422_/D _5359_/B _6879_/Q VGND VGND VPWR VPWR _3534_/X
+ sky130_fd_sc_hd__a32o_1
Xhold825 _5640_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR _7310_/A sky130_fd_sc_hd__clkbuf_2
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__clkbuf_2
Xhold836 _5572_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _5426_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap555 _4746_/A VGND VGND VPWR VPWR _4761_/A sky130_fd_sc_hd__clkbuf_2
Xhold858 _6775_/Q VGND VGND VPWR VPWR hold858/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap566 _4742_/C VGND VGND VPWR VPWR _4760_/C sky130_fd_sc_hd__buf_2
X_6253_ _7035_/Q _6465_/A2 _6465_/A3 _6122_/X _6891_/Q VGND VGND VPWR VPWR _6253_/X
+ sky130_fd_sc_hd__a32o_1
Xhold869 _5536_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3465_ _5620_/A _6548_/C _5684_/B VGND VGND VPWR VPWR _4204_/S sky130_fd_sc_hd__and3_4
XFILLER_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5204_ _5204_/A _5204_/B _5204_/C VGND VGND VPWR VPWR _5210_/A sky130_fd_sc_hd__and3_1
X_6184_ _6896_/Q _6129_/A _6097_/X _6968_/Q VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3396_ _3987_/A _6548_/D _5684_/B VGND VGND VPWR VPWR _3397_/B sky130_fd_sc_hd__and3_4
Xhold1503 _6069_/X VGND VGND VPWR VPWR _7205_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5135_ _5060_/C _4460_/C _5260_/C _5134_/X VGND VGND VPWR VPWR _5238_/A sky130_fd_sc_hd__a31o_1
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1514 _7220_/Q VGND VGND VPWR VPWR _6471_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 _7214_/Q VGND VGND VPWR VPWR _6343_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1536 _7254_/Q VGND VGND VPWR VPWR _3945_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _6803_/Q VGND VGND VPWR VPWR _3322_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_5066_ _5263_/B _4853_/C _4945_/C _4659_/B VGND VGND VPWR VPWR _5066_/X sky130_fd_sc_hd__o211a_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4017_ _6542_/A _4017_/B VGND VGND VPWR VPWR _4021_/S sky130_fd_sc_hd__nand2_4
XFILLER_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5968_ _6950_/Q _5779_/X _5782_/X _6942_/Q _5957_/X VGND VGND VPWR VPWR _5968_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4919_ _4919_/A _4919_/B VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__nand2_1
XFILLER_166_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5899_ _7043_/Q _5965_/B _5959_/B _5970_/B1 _6931_/Q VGND VGND VPWR VPWR _5899_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6940_ _7077_/CLK _6940_/D fanout587/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _6976_/CLK _6871_/D fanout590/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5822_ _6880_/Q _5768_/X _5794_/X _6920_/Q _5820_/X VGND VGND VPWR VPWR _5822_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5753_ _5757_/C _5703_/Y _6803_/Q VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__a21bo_1
XFILLER_147_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4704_ _4939_/A _4704_/B _4862_/A VGND VGND VPWR VPWR _4705_/B sky130_fd_sc_hd__and3_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5684_ _6548_/B _5684_/B _5684_/C VGND VGND VPWR VPWR _5692_/S sky130_fd_sc_hd__and3_4
XFILLER_187_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4635_ _4722_/A _4777_/A VGND VGND VPWR VPWR _4635_/Y sky130_fd_sc_hd__nand2_2
XFILLER_175_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 _4064_/X VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 _7263_/Q VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ _4761_/C _4320_/A _4301_/Y _4322_/Y _4870_/B VGND VGND VPWR VPWR _4574_/C
+ sky130_fd_sc_hd__o311a_1
Xhold622 hold622/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
Xhold633 hold633/A VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6305_/A _6305_/B _6305_/C _6305_/D VGND VGND VPWR VPWR _6305_/Y sky130_fd_sc_hd__nor4_1
Xhold644 hold644/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3517_ _7023_/Q _3515_/X _6542_/B _7270_/Q _3514_/X VGND VGND VPWR VPWR _3523_/B
+ sky130_fd_sc_hd__a221o_1
Xhold655 _4044_/X VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7285_ _7285_/A VGND VGND VPWR VPWR _7285_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold666 hold666/A VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap374 _6339_/D VGND VGND VPWR VPWR _6440_/D sky130_fd_sc_hd__buf_12
X_4497_ _5060_/A _4505_/B VGND VGND VPWR VPWR _4497_/Y sky130_fd_sc_hd__nand2_1
Xmax_cap385 _6141_/X VGND VGND VPWR VPWR _6452_/B1 sky130_fd_sc_hd__buf_12
Xhold677 hold677/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xhold688 _6623_/Q VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap396 _5777_/X VGND VGND VPWR VPWR _5971_/A2 sky130_fd_sc_hd__buf_12
X_6236_ _7138_/Q _6177_/C _6114_/X _6135_/X _6938_/Q VGND VGND VPWR VPWR _6236_/X
+ sky130_fd_sc_hd__a32o_1
Xhold699 _5526_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3448_ _7265_/Q hold17/A _4139_/C _3447_/X _6658_/Q VGND VGND VPWR VPWR _3448_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6167_ _6166_/X _5759_/A _5759_/B _6443_/S _6167_/B2 VGND VGND VPWR VPWR _7207_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _5476_/B _6536_/B _6536_/C _6530_/C VGND VGND VPWR VPWR _3384_/S sky130_fd_sc_hd__nand4_4
Xhold1300 _7238_/Q VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _7279_/Q VGND VGND VPWR VPWR hold799/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1322 _7155_/Q VGND VGND VPWR VPWR hold832/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5118_ _4408_/X _4722_/Y _4681_/C _5257_/C _4867_/C VGND VGND VPWR VPWR _5121_/D
+ sky130_fd_sc_hd__o2111a_1
Xhold1333 _5462_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6098_ _6143_/D _7187_/Q _6177_/A _6143_/C VGND VGND VPWR VPWR _6098_/X sky130_fd_sc_hd__and4_4
Xhold1344 _7040_/Q VGND VGND VPWR VPWR hold248/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1355 _7072_/Q VGND VGND VPWR VPWR hold671/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 _6741_/Q VGND VGND VPWR VPWR hold1366/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1377 _6836_/Q VGND VGND VPWR VPWR _5303_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ _4414_/X _5040_/X _5241_/D _5047_/X _5048_/X VGND VGND VPWR VPWR _5049_/Y
+ sky130_fd_sc_hd__o2111ai_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1388 _3356_/X VGND VGND VPWR VPWR hold1388/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _3402_/X VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4420_ _5060_/C _5260_/A _5140_/B _5143_/A _4860_/C VGND VGND VPWR VPWR _4441_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_129_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4351_ _4632_/C _5089_/C VGND VGND VPWR VPWR _4860_/C sky130_fd_sc_hd__nor2_8
XFILLER_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3302_ _7189_/Q _7190_/Q VGND VGND VPWR VPWR _6117_/A sky130_fd_sc_hd__and2b_2
X_7070_ _7132_/CLK _7070_/D fanout611/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4282_ _4310_/B _4984_/A _4282_/C _4760_/B VGND VGND VPWR VPWR _4282_/Y sky130_fd_sc_hd__nand4_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6021_ _6744_/Q _5788_/X _6009_/X _6012_/X _6020_/X VGND VGND VPWR VPWR _6021_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6923_ _7152_/CLK _6923_/D fanout587/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6854_ _7089_/CLK _6854_/D fanout596/X VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5805_ _7087_/Q _6072_/B wire398/X _5768_/X _6879_/Q VGND VGND VPWR VPWR _5805_/X
+ sky130_fd_sc_hd__a32o_1
X_6785_ _7006_/CLK _6785_/D fanout601/X VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtp_1
X_3997_ _3994_/S hold878/X _3502_/X _3922_/X VGND VGND VPWR VPWR _3997_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5736_ _6800_/Q _5759_/B _7186_/Q _5735_/Y VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__o31a_1
XFILLER_176_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5667_ _5667_/A0 _5667_/A1 _5674_/S VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__mux2_1
X_4618_ _4860_/B _4333_/Y _4512_/Y _4518_/X _4617_/Y VGND VGND VPWR VPWR _4618_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_163_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5598_ hold5/X _5598_/A1 hold14/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__mux2_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold430 hold430/A VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold441 _4123_/X VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4632_/B _4612_/C _4600_/B _4549_/D VGND VGND VPWR VPWR _4923_/B sky130_fd_sc_hd__and4bb_4
Xhold452 _6941_/Q VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _6989_/Q VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 _5391_/X VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7268_ _7268_/CLK _7268_/D fanout572/X VGND VGND VPWR VPWR _7268_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold485 _5623_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _7300_/A VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlygate4sd3_1
X_6219_ _7074_/Q _6425_/B _6425_/C _6129_/C _7154_/Q VGND VGND VPWR VPWR _6219_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7199_ _7251_/CLK _7199_/D fanout595/X VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1130 _5677_/X VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 _5312_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1152 _4128_/X VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1163 hold1358/X VGND VGND VPWR VPWR _5676_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1174 _3398_/X VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _5488_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1196 _5326_/X VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 _6109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 _6130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 _6995_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_336 _7085_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_347 _6789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 _6740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 _5815_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3920_ hold8/X _3913_/B _3918_/X _3914_/S hold656/X VGND VGND VPWR VPWR _3920_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_44_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3851_ input69/X _4092_/S _3445_/X _6893_/Q _3850_/X VGND VGND VPWR VPWR _3856_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ _6875_/CLK _6570_/D fanout596/X VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3782_ _6833_/Q _5325_/C _5311_/C _6987_/Q _3536_/X VGND VGND VPWR VPWR _3782_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_158_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5521_ _6548_/B _5548_/C _6548_/D hold28/X VGND VGND VPWR VPWR _5529_/S sky130_fd_sc_hd__and4_4
XFILLER_157_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5452_ hold316/X _3919_/C _5457_/S VGND VGND VPWR VPWR _5452_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4403_ _4247_/Y _4248_/X _4427_/C _4429_/D VGND VGND VPWR VPWR _4403_/X sky130_fd_sc_hd__a2bb2o_4
X_5383_ hold415/X _4049_/B _5385_/S VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__mux2_1
X_7122_ _7122_/CLK _7122_/D fanout607/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4334_ _5040_/C _4293_/Y _4299_/Y _4333_/Y VGND VGND VPWR VPWR _4487_/B sky130_fd_sc_hd__o22a_1
XFILLER_141_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7053_ _7053_/CLK _7053_/D fanout603/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfrtp_2
X_4265_ _5060_/B _5143_/D VGND VGND VPWR VPWR _4265_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6004_ _6028_/C _6072_/C _6679_/Q _5776_/X _6769_/Q VGND VGND VPWR VPWR _6004_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4196_ hold561/X _3921_/X _4204_/S VGND VGND VPWR VPWR _4196_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _7077_/CLK _6906_/D fanout587/X VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6837_ _7067_/CLK _6837_/D fanout582/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6768_ _6768_/CLK _6768_/D fanout576/X VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5719_ _7182_/Q _5712_/Y _5718_/X _5759_/B VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__a22o_1
X_6699_ _7053_/CLK _6699_/D fanout601/X VGND VGND VPWR VPWR _6699_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold260 _7043_/Q VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _5568_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _6876_/Q VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _6985_/Q VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_100 _6106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _6501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _6609_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _6593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 _7175_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_177 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _6003_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _6446_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4050_ hold320/X _4049_/B _4054_/S VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4952_ _4777_/B _4674_/C _4674_/D _4945_/C _4716_/A VGND VGND VPWR VPWR _4954_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_45_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3903_ _7142_/Q _3503_/X _3528_/X input19/X _3902_/X VGND VGND VPWR VPWR _3904_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4883_ _4862_/A _4718_/D _4792_/C _4465_/B VGND VGND VPWR VPWR _5002_/A sky130_fd_sc_hd__a31o_1
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6622_ _7268_/CLK _6622_/D fanout572/X VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfstp_2
X_3834_ _3834_/A _3834_/B _3834_/C _3834_/D VGND VGND VPWR VPWR _3834_/Y sky130_fd_sc_hd__nor4_1
XFILLER_137_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6553_ _3924_/B hold799/X _6553_/S VGND VGND VPWR VPWR _6553_/X sky130_fd_sc_hd__mux2_1
X_3765_ _6558_/Q _3359_/B _3463_/X _7115_/Q _3756_/X VGND VGND VPWR VPWR _3766_/D
+ sky130_fd_sc_hd__a221o_1
X_5504_ _5667_/A0 _5504_/A1 _5511_/S VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__mux2_1
X_6484_ _6514_/B _6514_/C _7259_/Q VGND VGND VPWR VPWR _6486_/B sky130_fd_sc_hd__a21bo_1
X_3696_ _6661_/Q _4158_/D _3446_/X _3492_/X _6666_/Q VGND VGND VPWR VPWR _3696_/X
+ sky130_fd_sc_hd__a32o_1
Xpad_flashh_clk_buff_inst input83/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_146_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5435_ _3921_/B hold603/X hold67/X VGND VGND VPWR VPWR _5435_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput310 _7315_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput321 hold581/X VGND VGND VPWR VPWR hold582/A sky130_fd_sc_hd__buf_12
Xoutput332 hold676/X VGND VGND VPWR VPWR hold677/A sky130_fd_sc_hd__buf_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 hold686/X VGND VGND VPWR VPWR hold687/A sky130_fd_sc_hd__buf_12
X_5366_ _5359_/B _4073_/X _5367_/S hold781/X VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4317_ _4313_/A _4346_/A _4670_/D _4313_/Y VGND VGND VPWR VPWR _4317_/Y sky130_fd_sc_hd__o211ai_1
X_7105_ _7129_/CLK _7105_/D fanout598/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5297_ _3916_/C hold303/X hold73/X VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7036_ _7171_/CLK _7036_/D fanout609/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_4
X_4248_ _4209_/Y _4246_/Y _4662_/B VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4179_ hold494/X _3921_/X _4187_/S VGND VGND VPWR VPWR _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout570 input99/X VGND VGND VPWR VPWR _4754_/B sky130_fd_sc_hd__clkbuf_8
Xfanout581 input75/X VGND VGND VPWR VPWR fanout581/X sky130_fd_sc_hd__buf_6
Xfanout592 fanout593/X VGND VGND VPWR VPWR fanout592/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_56_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7119_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3550_ _4127_/C _5666_/C _5575_/D VGND VGND VPWR VPWR _3550_/X sky130_fd_sc_hd__and3_4
XFILLER_155_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3481_ _6524_/A _6530_/D _5327_/D VGND VGND VPWR VPWR _3481_/X sky130_fd_sc_hd__and3_1
XFILLER_143_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5220_ _5220_/A _5220_/B _5220_/C _5220_/D VGND VGND VPWR VPWR _5220_/X sky130_fd_sc_hd__and4_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5151_ _4496_/Y _4658_/Y _4752_/B _4752_/D VGND VGND VPWR VPWR _5151_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4102_ _4053_/B _4102_/A1 _4102_/S VGND VGND VPWR VPWR _4102_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5082_ _5082_/A _5082_/B _5209_/A VGND VGND VPWR VPWR _5082_/Y sky130_fd_sc_hd__nand3_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4033_ hold24/X hold230/X _4034_/S VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5984_ _6748_/Q _5842_/C _6028_/C _6753_/Q _6073_/B2 VGND VGND VPWR VPWR _5984_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_80_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4935_ _5089_/A _4620_/C _4933_/Y _5033_/B VGND VGND VPWR VPWR _4976_/A sky130_fd_sc_hd__a211o_1
Xclkbuf_3_7_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 hold38/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _3438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4866_ _4377_/X _4411_/B _4496_/Y _4645_/Y VGND VGND VPWR VPWR _4867_/C sky130_fd_sc_hd__o2bb2a_1
XANTENNA_33 _5350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6605_ _6835_/CLK _6605_/D fanout582/X VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_55 _3657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3817_ _6932_/Q _3542_/B _5629_/C _5611_/B _7108_/Q VGND VGND VPWR VPWR _3817_/X
+ sky130_fd_sc_hd__a32o_1
X_4797_ _4549_/D _4208_/Y _4479_/Y _4796_/X _4795_/Y VGND VGND VPWR VPWR _4797_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA_66 _4358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_77 _5842_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_88 _5788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6536_/A _6536_/B _6536_/C _6536_/D VGND VGND VPWR VPWR _6541_/S sky130_fd_sc_hd__nand4_4
X_3748_ input6/X _3469_/X _5377_/C _6898_/Q _3747_/X VGND VGND VPWR VPWR _3751_/C
+ sky130_fd_sc_hd__a221o_2
XANTENNA_99 _6106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3679_ _7267_/Q _3564_/X _3674_/X _3676_/X _3678_/X VGND VGND VPWR VPWR _3679_/X
+ sky130_fd_sc_hd__a2111o_1
X_6467_ _6442_/S _6467_/A2 _6443_/S _6466_/X VGND VGND VPWR VPWR _6467_/X sky130_fd_sc_hd__a211o_1
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5418_ _5413_/B _3925_/X _5421_/S hold886/X VGND VGND VPWR VPWR _5418_/X sky130_fd_sc_hd__a22o_1
X_6398_ _6760_/Q _6097_/X _6462_/B1 _6655_/Q _6397_/X VGND VGND VPWR VPWR _6405_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput173 _3352_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
X_5349_ hold128/X _4053_/B _5349_/S VGND VGND VPWR VPWR _5349_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput184 _3267_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput195 _3257_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_102_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7019_ _7108_/CLK _7019_/D fanout606/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4720_/A _4720_/B _4720_/C _4720_/D VGND VGND VPWR VPWR _4723_/C sky130_fd_sc_hd__nand4_1
XFILLER_42_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4651_ _4804_/C _4945_/C _4755_/B VGND VGND VPWR VPWR _4678_/A sky130_fd_sc_hd__and3_1
XFILLER_175_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ _6764_/Q _3498_/X _3593_/X _3594_/X _3601_/X VGND VGND VPWR VPWR _3631_/A
+ sky130_fd_sc_hd__a2111o_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4582_ _4582_/A _4582_/B _4582_/C VGND VGND VPWR VPWR _4585_/A sky130_fd_sc_hd__nor3_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3533_ _5476_/B _5548_/D _3533_/C VGND VGND VPWR VPWR _5404_/B sky130_fd_sc_hd__and3_4
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_16
X_6321_ _7158_/Q _6129_/C _6118_/X _7062_/Q _6320_/X VGND VGND VPWR VPWR _6321_/X
+ sky130_fd_sc_hd__a221o_1
Xhold804 _5491_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 _5420_/X VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _7311_/A sky130_fd_sc_hd__clkbuf_4
Xhold826 _7052_/Q VGND VGND VPWR VPWR hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_2
Xhold837 _6688_/Q VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold848 _7028_/Q VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap556 _4600_/Y VGND VGND VPWR VPWR _4746_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6252_ _6907_/Q _6129_/D _6130_/X _6931_/Q _6251_/X VGND VGND VPWR VPWR _6255_/C
+ sky130_fd_sc_hd__a221o_1
Xhold859 _4155_/X VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3464_ _5630_/A _5630_/C _5675_/D VGND VGND VPWR VPWR _5639_/B sky130_fd_sc_hd__and3_4
XFILLER_115_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5203_ _4494_/C _4940_/C _4682_/B _4757_/X _5065_/X VGND VGND VPWR VPWR _5204_/A
+ sky130_fd_sc_hd__a311oi_1
X_6183_ _7024_/Q _6136_/X _6452_/B1 _6976_/Q _6182_/X VGND VGND VPWR VPWR _6190_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3395_ hold54/X hold16/X hold75/X hold65/A VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__and4b_2
XFILLER_97_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5134_ _5055_/D _5260_/B _5133_/X _4837_/X VGND VGND VPWR VPWR _5134_/X sky130_fd_sc_hd__a31o_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1504 _7194_/Q VGND VGND VPWR VPWR _5817_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1515 _7253_/Q VGND VGND VPWR VPWR _4168_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _7192_/Q VGND VGND VPWR VPWR _5756_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1537 _7258_/Q VGND VGND VPWR VPWR _7251_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5065_ _4712_/B _4754_/X _4755_/B _4939_/B VGND VGND VPWR VPWR _5065_/X sky130_fd_sc_hd__o211a_1
XFILLER_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1548 _6805_/Q VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__dlygate4sd3_1
X_4016_ hold962/X _6535_/A0 _4016_/S VGND VGND VPWR VPWR _4016_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5967_ _7054_/Q _5814_/X _5815_/X _7022_/Q _5966_/X VGND VGND VPWR VPWR _5967_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4918_ _4746_/A _5263_/C _4939_/B _4576_/B VGND VGND VPWR VPWR _4918_/X sky130_fd_sc_hd__a31o_1
X_5898_ _7067_/Q _5965_/B _5723_/X _5887_/X _5897_/X VGND VGND VPWR VPWR _5898_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_178_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4849_ _4849_/A _4987_/A VGND VGND VPWR VPWR _4849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6519_ _4152_/B _6519_/A1 _6523_/S VGND VGND VPWR VPWR _6519_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6870_ _7143_/CLK _6870_/D fanout587/X VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfrtp_1
X_5821_ _5934_/C _6072_/C _6888_/Q _5776_/X _6952_/Q VGND VGND VPWR VPWR _5821_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_179_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5752_ _5752_/A1 _5712_/Y _5751_/X _5752_/B2 VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4703_ _5255_/A _4791_/B _4923_/C VGND VGND VPWR VPWR _4705_/A sky130_fd_sc_hd__and3_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5683_ _5692_/A1 _5683_/A1 _5683_/S VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4634_ _4698_/A _4722_/A _4870_/B VGND VGND VPWR VPWR _4640_/A sky130_fd_sc_hd__and3_2
XFILLER_135_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold601 hold601/A VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _4565_/A _4565_/B _4565_/C _4565_/D VGND VGND VPWR VPWR _4570_/C sky130_fd_sc_hd__nand4_1
Xhold612 _6534_/X VGND VGND VPWR VPWR _7263_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _6593_/Q VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 hold634/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
X_6304_ _6933_/Q _6130_/X _6135_/X _6941_/Q _6303_/X VGND VGND VPWR VPWR _6305_/D
+ sky130_fd_sc_hd__a221o_1
X_3516_ _6524_/A _6536_/A _4127_/C VGND VGND VPWR VPWR _6542_/B sky130_fd_sc_hd__and3_4
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold645 _6706_/Q VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlygate4sd3_1
X_7284_ _7284_/A VGND VGND VPWR VPWR _7284_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold656 _6594_/Q VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlygate4sd3_1
X_4496_ _4689_/B _5036_/B _4860_/B _4632_/C VGND VGND VPWR VPWR _4496_/Y sky130_fd_sc_hd__nand4_4
Xhold667 _6646_/Q VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _6610_/Q VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap386 _6135_/X VGND VGND VPWR VPWR _6462_/B1 sky130_fd_sc_hd__buf_12
X_3447_ _5304_/A _5476_/B _4158_/D VGND VGND VPWR VPWR _3447_/X sky130_fd_sc_hd__and3_4
Xhold689 _3958_/X VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6235_ _7050_/Q _6130_/A _6110_/C _6097_/X _6970_/Q VGND VGND VPWR VPWR _6235_/X
+ sky130_fd_sc_hd__a32o_1
Xmax_cap397 _5773_/X VGND VGND VPWR VPWR _6003_/C sky130_fd_sc_hd__buf_12
XFILLER_103_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ wire347/X wire368/X _6871_/Q _6466_/A1 VGND VGND VPWR VPWR _6166_/X sky130_fd_sc_hd__o2bb2a_1
X_3378_ hold54/X hold16/X hold75/X _5324_/B VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__and4bb_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 _6852_/Q VGND VGND VPWR VPWR hold512/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1312 _6553_/X VGND VGND VPWR VPWR _7279_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 _5671_/X VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5117_ _4984_/A _4862_/A _4732_/C _4991_/X _5112_/X VGND VGND VPWR VPWR _5121_/C
+ sky130_fd_sc_hd__a311oi_1
XFILLER_69_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1334 _7251_/Q VGND VGND VPWR VPWR _7257_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6097_ _6143_/D _6141_/B _6138_/B _6143_/C VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__and4_4
Xhold1345 _6827_/Q VGND VGND VPWR VPWR hold954/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1356 _5577_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 _4113_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5048_ _5040_/C _5040_/B _5040_/A _4415_/X VGND VGND VPWR VPWR _5048_/X sky130_fd_sc_hd__a31o_1
Xhold1378 _6824_/Q VGND VGND VPWR VPWR hold372/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1389 _5556_/S VGND VGND VPWR VPWR _5550_/S sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6999_ _7130_/CLK _6999_/D fanout600/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4350_ _4984_/A _4788_/A _5044_/A VGND VGND VPWR VPWR _4465_/A sky130_fd_sc_hd__and3_1
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3301_ _7185_/Q _7186_/Q VGND VGND VPWR VPWR _6177_/A sky130_fd_sc_hd__and2b_4
XFILLER_98_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4281_ _4284_/C _4310_/B _4984_/A _4282_/C VGND VGND VPWR VPWR _4285_/A sky130_fd_sc_hd__nand4_4
XFILLER_98_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6020_ _6555_/Q _6025_/B _5842_/C _6016_/X _6019_/X VGND VGND VPWR VPWR _6020_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6922_ _7152_/CLK _6922_/D fanout587/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6853_ _7268_/CLK _6853_/D fanout572/X VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5804_ _6943_/Q _5779_/X _5783_/X _7007_/Q _5803_/X VGND VGND VPWR VPWR _5804_/X
+ sky130_fd_sc_hd__a221o_1
X_6784_ _7157_/CLK _6784_/D fanout592/X VGND VGND VPWR VPWR _7287_/A sky130_fd_sc_hd__dfrtp_1
X_3996_ _3994_/S hold773/X _3502_/X _3919_/X VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5735_ _5732_/X _6138_/B _5759_/B VGND VGND VPWR VPWR _5735_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5666_ _6524_/B _6548_/D _5666_/C hold28/X VGND VGND VPWR VPWR _5674_/S sky130_fd_sc_hd__nand4_4
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4617_ _4617_/A _4617_/B VGND VGND VPWR VPWR _4617_/Y sky130_fd_sc_hd__nand2_1
X_5597_ _3921_/B hold769/X hold14/X VGND VGND VPWR VPWR _5597_/X sky130_fd_sc_hd__mux2_1
Xhold420 _6684_/Q VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _7266_/Q VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _5090_/A _5090_/B _4615_/C _4786_/B VGND VGND VPWR VPWR _4554_/C sky130_fd_sc_hd__nand4_1
XFILLER_190_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold442 _6759_/Q VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold453 _5429_/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _5483_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold475 hold475/A VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _6754_/Q VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlygate4sd3_1
X_7267_ _7267_/CLK _7267_/D fanout572/X VGND VGND VPWR VPWR _7267_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_143_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4479_ _4792_/A _4788_/A VGND VGND VPWR VPWR _4479_/Y sky130_fd_sc_hd__nand2_1
Xhold497 _4068_/X VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6218_ _6217_/X _6242_/A2 _6343_/S VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__mux2_1
X_7198_ _7251_/CLK _7198_/D fanout595/X VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _6537_/X VGND VGND VPWR VPWR _7265_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ _7015_/Q _6177_/C _6110_/C _6143_/X _6943_/Q VGND VGND VPWR VPWR _6149_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1131 _6607_/Q VGND VGND VPWR VPWR _3940_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _7296_/A VGND VGND VPWR VPWR _4201_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 _6811_/Q VGND VGND VPWR VPWR _5274_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1164 hold1400/X VGND VGND VPWR VPWR _5459_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 hold1360/X VGND VGND VPWR VPWR _5522_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 hold1446/X VGND VGND VPWR VPWR _5504_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 _6718_/Q VGND VGND VPWR VPWR _4081_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_304 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_315 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _6995_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 _7105_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 _6845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_359 _6440_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3850_ _7061_/Q _3563_/A _3902_/A3 _5359_/B _6885_/Q VGND VGND VPWR VPWR _3850_/X
+ sky130_fd_sc_hd__a32o_1
X_3781_ _7075_/Q _3488_/X _3777_/X _3780_/X VGND VGND VPWR VPWR _3810_/A sky130_fd_sc_hd__a211o_2
X_5520_ _5692_/A1 hold911/X _5520_/S VGND VGND VPWR VPWR _5520_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5451_ hold387/X _3916_/C _5457_/S VGND VGND VPWR VPWR _5451_/X sky130_fd_sc_hd__mux2_1
X_4402_ _4427_/C _4429_/D _4383_/A VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__a21oi_4
X_5382_ hold352/X _3925_/C _5385_/S VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7121_ _7131_/CLK hold30/X fanout606/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_4
X_4333_ _4333_/A VGND VGND VPWR VPWR _4333_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4264_ _4429_/A _5143_/D _4429_/D VGND VGND VPWR VPWR _4505_/B sky130_fd_sc_hd__and3_2
X_7052_ _7122_/CLK _7052_/D fanout610/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_115_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6003_ _6608_/Q _6072_/B _6003_/C VGND VGND VPWR VPWR _6003_/X sky130_fd_sc_hd__and3_1
XFILLER_86_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4195_ _4195_/A0 _4194_/X _4205_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6905_ _7071_/CLK _6905_/D fanout585/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ _7067_/CLK _6836_/D fanout582/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6767_ _6780_/CLK _6767_/D fanout575/X VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3979_ hold207/X hold24/X _3980_/S VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__mux2_1
X_5718_ _7182_/Q _5782_/C VGND VGND VPWR VPWR _5718_/X sky130_fd_sc_hd__xor2_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6698_ _7053_/CLK _6698_/D fanout601/X VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5649_ _5649_/A0 hold780/X _5656_/S VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold250 _5553_/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold261 _5544_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold272 _7306_/A VGND VGND VPWR VPWR hold272/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold283 _5356_/X VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _5479_/X VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _6141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_123 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _7059_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _7206_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_178 input164/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _6003_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4951_ _4753_/A _4512_/Y _5248_/A3 _4650_/Y VGND VGND VPWR VPWR _4951_/X sky130_fd_sc_hd__o31a_1
XFILLER_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3902_ _7062_/Q _3563_/A _3902_/A3 _3504_/X input33/X VGND VGND VPWR VPWR _3902_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4882_ _4704_/B _4375_/X _5128_/B _4705_/A VGND VGND VPWR VPWR _4884_/B sky130_fd_sc_hd__a31o_1
X_6621_ _7273_/CLK _6621_/D fanout579/X VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfrtp_4
X_3833_ input40/X _4187_/S _3503_/X _7140_/Q _3832_/X VGND VGND VPWR VPWR _3834_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6552_ hold24/X hold196/X _6553_/S VGND VGND VPWR VPWR _6552_/X sky130_fd_sc_hd__mux2_1
X_3764_ hold91/A _3438_/X _5611_/B _7107_/Q _3763_/X VGND VGND VPWR VPWR _3766_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5503_ hold66/X _5503_/B VGND VGND VPWR VPWR _5511_/S sky130_fd_sc_hd__nand2_8
X_6483_ _6514_/C _6483_/B VGND VGND VPWR VPWR _6483_/Y sky130_fd_sc_hd__nand2_1
X_3695_ _6781_/Q _5311_/B _3533_/C _3502_/X _6656_/Q VGND VGND VPWR VPWR _3695_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_145_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput300 _6841_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_5434_ hold2/X _5434_/A1 hold67/X VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__mux2_1
XFILLER_173_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput311 _7316_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
Xoutput322 hold469/X VGND VGND VPWR VPWR hold470/A sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput333 hold635/X VGND VGND VPWR VPWR hold636/A sky130_fd_sc_hd__buf_12
Xoutput344 hold526/X VGND VGND VPWR VPWR hold527/A sky130_fd_sc_hd__buf_12
X_5365_ _6505_/A1 hold852/X _5367_/S VGND VGND VPWR VPWR _5365_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_3_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_113_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7104_ _7167_/CLK _7104_/D fanout604/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfstp_1
X_4316_ _4313_/A _4346_/A _4670_/D _4313_/Y VGND VGND VPWR VPWR _5090_/B sky130_fd_sc_hd__o211a_4
X_5296_ _5649_/A0 _5296_/A1 hold73/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7035_ _7035_/CLK _7035_/D fanout591/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4247_ _4427_/D _4320_/A VGND VGND VPWR VPWR _4247_/Y sky130_fd_sc_hd__nor2_2
XFILLER_68_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4178_ _4178_/A0 _4177_/X _4188_/S VGND VGND VPWR VPWR _4178_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6819_ _7265_/CLK _6819_/D fanout575/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire438 _4792_/A VGND VGND VPWR VPWR _4804_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout560 _4422_/Y VGND VGND VPWR VPWR _4945_/B sky130_fd_sc_hd__buf_4
Xfanout571 fanout581/X VGND VGND VPWR VPWR _3291_/A sky130_fd_sc_hd__buf_8
Xfanout582 fanout584/X VGND VGND VPWR VPWR fanout582/X sky130_fd_sc_hd__buf_8
XFILLER_120_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout593 input75/X VGND VGND VPWR VPWR fanout593/X sky130_fd_sc_hd__buf_6
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3480_ _6548_/C _6548_/D _5684_/B VGND VGND VPWR VPWR _3913_/B sky130_fd_sc_hd__and3_4
XFILLER_170_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _5235_/D _5148_/Y _5130_/X _5107_/X VGND VGND VPWR VPWR _5150_/X sky130_fd_sc_hd__a211o_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4101_ _5494_/A _3571_/X _4051_/X _4102_/S _4101_/B2 VGND VGND VPWR VPWR _4101_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5081_ _4788_/A _4950_/X _5080_/X VGND VGND VPWR VPWR _5209_/A sky130_fd_sc_hd__a21oi_1
X_4032_ _6539_/A0 _4032_/A1 _4034_/S VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5983_ _7270_/Q _5780_/X _5980_/X _5981_/X _5982_/X VGND VGND VPWR VPWR _5983_/X
+ sky130_fd_sc_hd__a2111o_1
X_4934_ _4939_/A _4620_/A _4595_/A _4607_/A VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__a31o_1
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4865_ _4864_/Y _4852_/X _4983_/B _4865_/D VGND VGND VPWR VPWR _4867_/B sky130_fd_sc_hd__and4bb_1
XANTENNA_12 hold38/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _3438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _6945_/CLK _6604_/D fanout583/X VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_34 _5350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3816_ _7036_/Q _3547_/X _5593_/B _7092_/Q _3815_/X VGND VGND VPWR VPWR _3825_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_45 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _3710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _4271_/Y _4293_/Y _4479_/Y _4633_/Y VGND VGND VPWR VPWR _4796_/X sky130_fd_sc_hd__o22a_1
XFILLER_177_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_67 _4849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _5773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6535_ _6535_/A0 _6535_/A1 _6535_/S VGND VGND VPWR VPWR _6535_/X sky130_fd_sc_hd__mux2_1
XANTENNA_89 _5788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3747_ _6914_/Q _5422_/D _5281_/A2 _3528_/X input14/X VGND VGND VPWR VPWR _3747_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_180_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6466_ _6466_/A1 _6692_/Q _6465_/X _6458_/X _5759_/A VGND VGND VPWR VPWR _6466_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3678_ _7081_/Q _3413_/X _3565_/X _6650_/Q _3677_/X VGND VGND VPWR VPWR _3678_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_161_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5417_ _3921_/B hold567/X _5421_/S VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6397_ _7241_/Q _6177_/C _6114_/X _6130_/X _6780_/Q VGND VGND VPWR VPWR _6397_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput174 _3353_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
X_5348_ hold530/X _4051_/B _5349_/S VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__mux2_1
Xoutput185 _3266_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3256_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5279_ _5476_/B _6536_/B _5575_/D _5279_/D VGND VGND VPWR VPWR _5280_/S sky130_fd_sc_hd__nand4_2
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7018_ _7117_/CLK _7018_/D fanout605/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4650_ _4804_/C _4945_/C VGND VGND VPWR VPWR _4650_/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3601_ _6621_/Q _3954_/B _3597_/X _3598_/X _3600_/X VGND VGND VPWR VPWR _3601_/X
+ sky130_fd_sc_hd__a2111o_1
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4581_ _5140_/C _4581_/B _4589_/C VGND VGND VPWR VPWR _4582_/B sky130_fd_sc_hd__and3_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
X_6320_ _6894_/Q _6122_/X _6129_/D _6910_/Q _6319_/X VGND VGND VPWR VPWR _6320_/X
+ sky130_fd_sc_hd__a221o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7316_/A sky130_fd_sc_hd__buf_2
X_3532_ _5575_/C _5422_/D _5575_/D VGND VGND VPWR VPWR _5359_/B sky130_fd_sc_hd__and3_4
XFILLER_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold805 _7108_/Q VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 qspi_enabled VGND VGND VPWR VPWR _3327_/A sky130_fd_sc_hd__buf_6
Xhold816 _7100_/Q VGND VGND VPWR VPWR hold816/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7312_/A sky130_fd_sc_hd__clkbuf_2
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold827 _5554_/X VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 _4036_/X VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap546 _4747_/Y VGND VGND VPWR VPWR _4789_/D sky130_fd_sc_hd__clkbuf_2
Xhold849 _5527_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _7043_/Q _6444_/C _6108_/X _6104_/X _7163_/Q VGND VGND VPWR VPWR _6251_/X
+ sky130_fd_sc_hd__a32o_1
X_3463_ _5620_/A _5630_/A _5675_/D VGND VGND VPWR VPWR _3463_/X sky130_fd_sc_hd__and3_4
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5202_ _5235_/D _5188_/Y _5198_/X _4981_/X _5180_/Y VGND VGND VPWR VPWR _5202_/X
+ sky130_fd_sc_hd__a221o_1
X_6182_ _7088_/Q _6136_/A _6102_/X _6109_/X _7040_/Q VGND VGND VPWR VPWR _6182_/X
+ sky130_fd_sc_hd__a32o_1
X_3394_ hold42/X hold37/X _5324_/B VGND VGND VPWR VPWR _5449_/B sky130_fd_sc_hd__and3b_4
X_5133_ _4729_/A _5044_/A _4557_/B _4878_/A VGND VGND VPWR VPWR _5133_/X sky130_fd_sc_hd__a31o_1
XFILLER_97_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1505 _7202_/Q VGND VGND VPWR VPWR _6023_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1516 _7196_/Q VGND VGND VPWR VPWR _5862_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1527 _6629_/Q VGND VGND VPWR VPWR _3965_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1538 _7257_/Q VGND VGND VPWR VPWR _7254_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5064_ _5089_/C _4789_/B _4734_/X _4805_/X VGND VGND VPWR VPWR _5064_/X sky130_fd_sc_hd__a31o_1
Xhold1549 _7253_/Q VGND VGND VPWR VPWR _6470_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_4015_ hold587/X _6546_/A0 _4016_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5966_ _7014_/Q _5783_/X _5791_/X _7126_/Q _5965_/X VGND VGND VPWR VPWR _5966_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4917_ _4490_/Y _4537_/X _4567_/Y _4629_/Y _4745_/Y VGND VGND VPWR VPWR _4919_/B
+ sky130_fd_sc_hd__o32a_1
X_5897_ _7051_/Q _5814_/X _5815_/X _7019_/Q _5896_/X VGND VGND VPWR VPWR _5897_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4848_ _4848_/A _4848_/B _4987_/A VGND VGND VPWR VPWR _4857_/C sky130_fd_sc_hd__and3_1
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4779_ _4779_/A _4779_/B _4779_/C VGND VGND VPWR VPWR _4779_/Y sky130_fd_sc_hd__nor3_1
XFILLER_148_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6518_ _6536_/A _6536_/B _6536_/C _6530_/D VGND VGND VPWR VPWR _6523_/S sky130_fd_sc_hd__nand4_4
XFILLER_4_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6449_ _6747_/Q _6446_/B _6347_/C _6129_/A _6677_/Q VGND VGND VPWR VPWR _6449_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_122_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6908_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_csclk _7277_/CLK VGND VGND VPWR VPWR _7065_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5820_ _7032_/Q _6072_/B _6003_/C _5819_/X VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__a31o_1
XFILLER_62_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5751_ _5741_/Y _7190_/Q _6117_/A _5750_/X VGND VGND VPWR VPWR _5751_/X sky130_fd_sc_hd__a211o_1
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4702_ _4650_/Y _4699_/Y _4700_/Y _4697_/Y VGND VGND VPWR VPWR _4705_/C sky130_fd_sc_hd__o211ai_1
XFILLER_148_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5682_ hold13/X _3509_/X _4051_/X _5683_/S hold739/X VGND VGND VPWR VPWR _5682_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_30_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4633_ _4940_/C _4633_/B VGND VGND VPWR VPWR _4633_/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4564_ _4321_/Y _4322_/Y _4509_/A _4527_/X _5040_/C VGND VGND VPWR VPWR _4565_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold602 hold602/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
XFILLER_128_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold613 _6702_/Q VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6303_ _7037_/Q _6465_/A2 _6465_/A3 _6115_/X _7141_/Q VGND VGND VPWR VPWR _6303_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold624 _3917_/X VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _5548_/C _6548_/D hold28/A VGND VGND VPWR VPWR _3515_/X sky130_fd_sc_hd__and3_4
Xhold635 hold635/A VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlygate4sd3_1
X_7283_ _7283_/A VGND VGND VPWR VPWR _7283_/X sky130_fd_sc_hd__clkbuf_1
Xhold646 _4063_/X VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _4632_/C _4940_/C _4860_/B VGND VGND VPWR VPWR _4718_/D sky130_fd_sc_hd__and3_4
Xhold657 _3920_/X VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 _3985_/X VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold679 _3943_/X VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6930_/Q _6130_/X _6452_/B1 _6978_/Q _6233_/X VGND VGND VPWR VPWR _6239_/B
+ sky130_fd_sc_hd__a221o_1
Xmax_cap387 _6126_/X VGND VGND VPWR VPWR _6323_/B1 sky130_fd_sc_hd__buf_8
XFILLER_170_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3446_ _6805_/Q _5620_/A hold65/A _6804_/Q VGND VGND VPWR VPWR _3446_/X sky130_fd_sc_hd__and4b_4
XFILLER_131_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6165_/A _6165_/B _6165_/C _6440_/D VGND VGND VPWR VPWR _6165_/Y sky130_fd_sc_hd__nor4_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _6535_/A0 _3377_/A1 _3377_/S VGND VGND VPWR VPWR _3377_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _5328_/X VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5116_ _4862_/A _4854_/X _5111_/X _5115_/X VGND VGND VPWR VPWR _5258_/A sky130_fd_sc_hd__a211oi_2
XFILLER_57_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1313 _7031_/Q VGND VGND VPWR VPWR hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 _6911_/Q VGND VGND VPWR VPWR hold1324/X sky130_fd_sc_hd__dlygate4sd3_1
X_6096_ _6143_/D _6141_/B _6134_/C VGND VGND VPWR VPWR _6096_/Y sky130_fd_sc_hd__nor3_4
Xhold1335 _6770_/Q VGND VGND VPWR VPWR hold417/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 _5293_/X VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1357 _6830_/Q VGND VGND VPWR VPWR hold303/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 _6622_/Q VGND VGND VPWR VPWR hold1368/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5047_ _5040_/C _5040_/B _4358_/X _4403_/X VGND VGND VPWR VPWR _5047_/X sky130_fd_sc_hd__a211o_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1379 _5290_/X VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6998_ _7132_/CLK _6998_/D fanout611/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfrtp_2
X_5949_ _7093_/Q _6072_/B wire398/X _5795_/X _6901_/Q VGND VGND VPWR VPWR _5949_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ _5759_/A _3300_/B _3307_/B VGND VGND VPWR VPWR _3300_/Y sky130_fd_sc_hd__nor3_1
XFILLER_125_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4280_ _4280_/A _4280_/B VGND VGND VPWR VPWR _4284_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6921_ _7073_/CLK _6921_/D fanout582/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6852_ _7089_/CLK _6852_/D fanout580/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_4
X_5803_ _7095_/Q _5780_/X _5784_/X _7023_/Q VGND VGND VPWR VPWR _5803_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6783_ _7237_/CLK _6783_/D _6472_/A VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfrtp_1
X_3995_ _3994_/S hold907/X _3502_/X _3916_/X VGND VGND VPWR VPWR _3995_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5734_ _7186_/Q _7185_/Q VGND VGND VPWR VPWR _6117_/C sky130_fd_sc_hd__and2b_4
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5665_ _5692_/A1 _5665_/A1 _5665_/S VGND VGND VPWR VPWR _5665_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4616_ _4815_/A _4620_/A _4615_/C _4615_/X _5216_/B VGND VGND VPWR VPWR _4617_/B
+ sky130_fd_sc_hd__a311oi_1
X_5596_ _3918_/B hold522/X hold14/X VGND VGND VPWR VPWR _5596_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold410 _5481_/X VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _4031_/X VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _5090_/A _5090_/B _5128_/B _4620_/B VGND VGND VPWR VPWR _4554_/B sky130_fd_sc_hd__nand4_1
Xhold432 _6538_/X VGND VGND VPWR VPWR _7266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _4135_/X VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold454 _6558_/Q VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7266_ _7269_/CLK _7266_/D fanout576/X VGND VGND VPWR VPWR _7266_/Q sky130_fd_sc_hd__dfrtp_4
Xhold465 _6728_/Q VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold476 _6781_/Q VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4730_/A _4799_/B _4674_/C VGND VGND VPWR VPWR _4480_/B sky130_fd_sc_hd__and3_2
Xhold487 _4129_/X VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 hold498/A VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6217_ _6292_/S _6217_/A2 _6215_/Y _6216_/X VGND VGND VPWR VPWR _6217_/X sky130_fd_sc_hd__a22o_1
X_3429_ input93/X _3902_/A3 _3721_/A3 _3428_/X _7007_/Q VGND VGND VPWR VPWR _3437_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_58_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7197_ _7251_/CLK _7197_/D fanout595/X VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _7031_/Q _6138_/X _6144_/X _7079_/Q _6147_/X VGND VGND VPWR VPWR _6148_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1110 _5332_/X VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _6935_/Q VGND VGND VPWR VPWR _5423_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1132 _3940_/X VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 _4201_/X VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 _5274_/X VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6079_ _6611_/Q _5782_/C _5814_/C _6009_/C _6652_/Q VGND VGND VPWR VPWR _6079_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1165 hold1349/X VGND VGND VPWR VPWR _5603_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 _7297_/A VGND VGND VPWR VPWR _4203_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 _7283_/A VGND VGND VPWR VPWR _4085_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 _6113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1198 _4081_/X VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 _6175_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_327 _6995_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 _7276_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 _6805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3780_ _6692_/Q _3386_/X _5327_/D _3779_/X VGND VGND VPWR VPWR _3780_/X sky130_fd_sc_hd__a31o_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5450_ _5450_/A0 _5667_/A0 _5457_/S VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4401_ _4848_/A _4356_/A _4392_/Y _4295_/A _4348_/X VGND VGND VPWR VPWR _4450_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_172_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5381_ _3249_/Y _5385_/S _3922_/X _5377_/C VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_160_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7120_ _7120_/CLK _7120_/D fanout607/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4332_ _4615_/C _4517_/B _5090_/B VGND VGND VPWR VPWR _4333_/A sky130_fd_sc_hd__and3_4
XFILLER_153_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7051_ _7131_/CLK _7051_/D fanout606/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_141_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4263_ _4209_/Y _4246_/Y _4848_/A _4356_/A VGND VGND VPWR VPWR _4263_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6002_ _6812_/Q _6028_/C _5782_/C _5795_/C VGND VGND VPWR VPWR _6002_/X sky130_fd_sc_hd__o211a_1
XFILLER_140_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4194_ hold569/X _3918_/X _4204_/S VGND VGND VPWR VPWR _4194_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6904_ _7171_/CLK _6904_/D fanout610/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6835_ _6835_/CLK _6835_/D fanout582/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfstp_2
X_6766_ _7241_/CLK _6766_/D fanout575/X VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3978_ hold304/X _3918_/B _3980_/S VGND VGND VPWR VPWR _3978_/X sky130_fd_sc_hd__mux2_1
X_5717_ _7181_/Q _7180_/Q _5716_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__a21o_1
XFILLER_109_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6697_ _7053_/CLK _6697_/D fanout601/X VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ _6548_/B _5684_/B _5657_/D hold27/X VGND VGND VPWR VPWR _5656_/S sky130_fd_sc_hd__nand4_4
XFILLER_191_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5579_ hold559/X _3921_/B hold18/X VGND VGND VPWR VPWR _5579_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold240 _7307_/A VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _7060_/Q VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold262 _6998_/Q VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _4075_/X VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _6846_/Q VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _6865_/Q VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ _7256_/CLK _7249_/D _6472_/A VGND VGND VPWR VPWR _7249_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _6144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_124 _6767_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _6565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _7219_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _3313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4950_ _4940_/C _4789_/B _4645_/A _4777_/C VGND VGND VPWR VPWR _4950_/X sky130_fd_sc_hd__a31o_2
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3901_ input42/X _4187_/S _3474_/X _7150_/Q _3900_/X VGND VGND VPWR VPWR _3904_/C
+ sky130_fd_sc_hd__a221o_1
X_4881_ _4881_/A _4881_/B VGND VGND VPWR VPWR _4884_/A sky130_fd_sc_hd__nand2_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6620_ _7267_/CLK _6620_/D _3291_/A VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_4
X_3832_ input31/X _3466_/X _5311_/C _6972_/Q _5458_/B VGND VGND VPWR VPWR _3832_/X
+ sky130_fd_sc_hd__a32o_2
X_6551_ _3918_/B hold959/X _6553_/S VGND VGND VPWR VPWR _6551_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3763_ _6687_/Q _4029_/B _5350_/B _6875_/Q VGND VGND VPWR VPWR _3763_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5502_ _5502_/A0 _5692_/A1 _5502_/S VGND VGND VPWR VPWR _5502_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6482_ _6514_/C _6482_/B VGND VGND VPWR VPWR _6482_/Y sky130_fd_sc_hd__nand2_1
X_3694_ _3693_/Y _3694_/A1 _3906_/S VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5433_ _3916_/C hold375/X hold67/X VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput301 _6842_/Q VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
Xoutput312 _7317_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput323 hold557/X VGND VGND VPWR VPWR hold558/A sky130_fd_sc_hd__buf_12
XFILLER_133_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5364_ _5359_/B _3925_/X _5367_/S hold984/X VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__a22o_1
Xoutput334 hold754/X VGND VGND VPWR VPWR hold755/A sky130_fd_sc_hd__buf_12
Xoutput345 hold585/X VGND VGND VPWR VPWR hold586/A sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7103_ _7167_/CLK _7103_/D fanout604/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfstp_4
X_4315_ _4284_/A _4308_/Y _4314_/X VGND VGND VPWR VPWR _4544_/A sky130_fd_sc_hd__o21ai_4
X_5295_ _6524_/B _6548_/C _6530_/D _5295_/D VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__nand4_4
XFILLER_141_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7034_ _7114_/CLK _7034_/D fanout604/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_4
X_4246_ _4656_/C _4647_/C VGND VGND VPWR VPWR _4246_/Y sky130_fd_sc_hd__nand2_8
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4177_ hold301/X _3918_/X _4187_/S VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6818_ _6827_/CLK _6818_/D fanout573/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire406 _4170_/C VGND VGND VPWR VPWR wire406/X sky130_fd_sc_hd__clkbuf_2
X_6749_ _6768_/CLK _6749_/D fanout576/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout572 fanout581/X VGND VGND VPWR VPWR fanout572/X sky130_fd_sc_hd__buf_6
Xfanout583 fanout584/X VGND VGND VPWR VPWR fanout583/X sky130_fd_sc_hd__buf_8
Xfanout594 fanout595/X VGND VGND VPWR VPWR fanout594/X sky130_fd_sc_hd__buf_6
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4100_ hold83/X hold94/X _4102_/S VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__mux2_1
XFILLER_110_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5080_ _4939_/A _5128_/C _4789_/D _4788_/X VGND VGND VPWR VPWR _5080_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4031_ _6538_/A0 hold420/X _4034_/S VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5982_ _6554_/Q _6025_/B _5842_/C _5784_/X _6620_/Q VGND VGND VPWR VPWR _5982_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4933_ _4929_/X _4933_/B _4933_/C VGND VGND VPWR VPWR _4933_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4864_ _4856_/X _4864_/B _4864_/C VGND VGND VPWR VPWR _4864_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_178_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_13 _3407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6835_/CLK _6603_/D fanout582/X VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_2
X_3815_ _7100_/Q _6548_/A _6548_/D _5675_/D _3814_/X VGND VGND VPWR VPWR _3815_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA_24 _3438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_35 _5350_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_46 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4795_ _4860_/B _5082_/A _4793_/X _4790_/Y VGND VGND VPWR VPWR _4795_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_177_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_57 _3758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _6540_/A0 hold611/X _6535_/S VGND VGND VPWR VPWR _6534_/X sky130_fd_sc_hd__mux2_1
XANTENNA_68 _4827_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3746_ _7146_/Q _3474_/X _3742_/X _3743_/X _3745_/X VGND VGND VPWR VPWR _3751_/B
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_79 _5773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6465_ _6611_/Q _6465_/A2 _6465_/A3 _6461_/X _6464_/X VGND VGND VPWR VPWR _6465_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_146_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3677_ _7129_/Q _6548_/A hold39/A _3558_/X _6609_/Q VGND VGND VPWR VPWR _3677_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5416_ _5413_/B _3919_/X _5421_/S hold771/X VGND VGND VPWR VPWR _5416_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6396_ _6604_/Q _6105_/X _6451_/B1 _6665_/Q _6395_/X VGND VGND VPWR VPWR _6396_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5347_ hold102/X hold83/X _5349_/S VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput175 _3338_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 _3348_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3282_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5278_ _6535_/A0 _5278_/A1 _5278_/S VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7017_ _7017_/CLK _7017_/D fanout598/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_4
X_4229_ _4229_/A _4229_/B _4229_/C _4229_/D VGND VGND VPWR VPWR _4230_/B sky130_fd_sc_hd__nand4_4
XFILLER_75_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout380 _5044_/A VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__buf_4
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3600_ _6853_/Q _5311_/B _5327_/D _3599_/X VGND VGND VPWR VPWR _3600_/X sky130_fd_sc_hd__a31o_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
X_4580_ _4815_/A _4584_/B _4923_/A _4589_/C VGND VGND VPWR VPWR _4582_/A sky130_fd_sc_hd__and4_1
XFILLER_190_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3531_ _6536_/C _4127_/C _5273_/D VGND VGND VPWR VPWR _3531_/X sky130_fd_sc_hd__and3_2
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7317_/A sky130_fd_sc_hd__buf_2
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold806 _5617_/X VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 _5608_/X VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _7145_/Q VGND VGND VPWR VPWR hold828/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _7313_/A sky130_fd_sc_hd__clkbuf_4
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__clkbuf_1
Xhold839 _6925_/Q VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlygate4sd3_1
X_6250_ _7067_/Q _6103_/X _6143_/X _6947_/Q _6249_/X VGND VGND VPWR VPWR _6255_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap547 _5173_/C VGND VGND VPWR VPWR _4756_/C sky130_fd_sc_hd__clkbuf_2
X_3462_ _3462_/A _3462_/B _3462_/C _3462_/D VGND VGND VPWR VPWR _3508_/B sky130_fd_sc_hd__nor4_1
XFILLER_143_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5201_ _5128_/A _4815_/A _5128_/C _4729_/X _5128_/X VGND VGND VPWR VPWR _5226_/B
+ sky130_fd_sc_hd__a311oi_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6181_ _6181_/A _6181_/B _6181_/C _6181_/D VGND VGND VPWR VPWR _6181_/Y sky130_fd_sc_hd__nor4_1
X_3393_ _3924_/B hold752/X _3393_/S VGND VGND VPWR VPWR _3393_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5132_ _5128_/B _5140_/C _5143_/A VGND VGND VPWR VPWR _5132_/Y sky130_fd_sc_hd__o21ai_2
Xhold1506 _7203_/Q VGND VGND VPWR VPWR _6024_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 _7200_/Q VGND VGND VPWR VPWR _5955_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5063_ _5149_/C _5061_/X _5062_/X _4266_/Y VGND VGND VPWR VPWR _5087_/A sky130_fd_sc_hd__a31o_1
XFILLER_96_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1528 _7211_/Q VGND VGND VPWR VPWR _6268_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _7175_/Q VGND VGND VPWR VPWR _5695_/A3 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4014_ hold945/X _6539_/A0 _4016_/S VGND VGND VPWR VPWR _4014_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5965_ _7070_/Q _5965_/B _6010_/C _6010_/D VGND VGND VPWR VPWR _5965_/X sky130_fd_sc_hd__and4_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4916_ _4898_/X _4916_/B _5264_/D VGND VGND VPWR VPWR _4919_/A sky130_fd_sc_hd__and3b_1
X_5896_ _7011_/Q _5826_/B _5815_/B _5783_/C _5895_/X VGND VGND VPWR VPWR _5896_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4847_ _4633_/Y _4638_/Y _4648_/Y _4444_/B VGND VGND VPWR VPWR _5120_/A sky130_fd_sc_hd__o31a_1
X_4778_ _5263_/B _4939_/B _4778_/C VGND VGND VPWR VPWR _4779_/B sky130_fd_sc_hd__and3_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3729_ _7018_/Q _3499_/X _3718_/X _3721_/X _3728_/X VGND VGND VPWR VPWR _3729_/X
+ sky130_fd_sc_hd__a2111o_1
X_6517_ _4166_/B _6469_/Y _6513_/X _6516_/X VGND VGND VPWR VPWR _7238_/D sky130_fd_sc_hd__a31o_1
XFILLER_107_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6448_ _7248_/Q _6103_/X _6126_/X _6767_/Q _6446_/X VGND VGND VPWR VPWR _6448_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6379_ _6679_/Q _6122_/X _6126_/X _6764_/Q _6378_/X VGND VGND VPWR VPWR _6380_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5750_ _7186_/Q _7185_/Q _5750_/C VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__and3_4
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4701_ _4939_/B _4923_/C VGND VGND VPWR VPWR _4701_/Y sky130_fd_sc_hd__nand2_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _4049_/B hold286/X _5683_/S VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4632_ _4632_/A _4632_/B _4632_/C _4729_/A VGND VGND VPWR VPWR _4799_/C sky130_fd_sc_hd__nor4_2
XFILLER_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4563_ _4321_/Y _4322_/Y _4509_/A _4490_/Y _4527_/X VGND VGND VPWR VPWR _4565_/B
+ sky130_fd_sc_hd__a2111o_1
Xhold603 _6946_/Q VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _6564_/Q _5311_/B _6530_/C _3513_/X _6668_/Q VGND VGND VPWR VPWR _3514_/X
+ sky130_fd_sc_hd__a32o_1
X_6302_ _7149_/Q _6113_/X _6323_/B1 _6965_/Q _6301_/X VGND VGND VPWR VPWR _6305_/C
+ sky130_fd_sc_hd__a221o_1
Xhold614 _4059_/X VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7282_ _7282_/A VGND VGND VPWR VPWR _7282_/X sky130_fd_sc_hd__clkbuf_1
Xhold625 _6871_/Q VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold636 hold636/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
X_4494_ _4689_/B _5036_/B _4494_/C VGND VGND VPWR VPWR _4653_/B sky130_fd_sc_hd__and3_1
Xhold647 _6814_/Q VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _6986_/Q VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _6994_/Q _6176_/B _6143_/C _6122_/X _6890_/Q VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3445_ _5476_/C _5575_/C _3533_/C VGND VGND VPWR VPWR _3445_/X sky130_fd_sc_hd__and3_4
Xhold669 _6909_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap388 _6120_/X VGND VGND VPWR VPWR _6451_/B1 sky130_fd_sc_hd__buf_12
XFILLER_171_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap399 _5764_/X VGND VGND VPWR VPWR _6086_/B1 sky130_fd_sc_hd__buf_8
XFILLER_143_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _7127_/Q _6116_/X _6452_/B1 _6975_/Q _6163_/X VGND VGND VPWR VPWR _6165_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _6546_/A0 hold506/X _3377_/S VGND VGND VPWR VPWR _3376_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5115_ _4375_/X _4712_/B _4903_/B _4987_/X VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__a31o_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _6640_/Q VGND VGND VPWR VPWR hold304/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _5531_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6095_ _7185_/Q _7190_/Q _7189_/Q _7186_/Q VGND VGND VPWR VPWR _6110_/C sky130_fd_sc_hd__and4bb_4
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 _5396_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1336 _7152_/Q VGND VGND VPWR VPWR hold798/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1347 _6680_/Q VGND VGND VPWR VPWR hold978/A sky130_fd_sc_hd__dlygate4sd3_1
X_5046_ _4358_/X _4403_/X _5040_/A _5142_/D VGND VGND VPWR VPWR _5241_/D sky130_fd_sc_hd__o31a_1
Xhold1358 _7159_/Q VGND VGND VPWR VPWR hold1358/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 _6636_/Q VGND VGND VPWR VPWR hold475/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6997_ _7140_/CLK hold80/X fanout609/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__dfrtp_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5948_ _7109_/Q _5764_/X _5784_/X _7029_/Q _5947_/X VGND VGND VPWR VPWR _5948_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5879_ _7042_/Q _5826_/B _5959_/B _5971_/A2 _7074_/Q VGND VGND VPWR VPWR _5879_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_138_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6920_ _7015_/CLK _6920_/D fanout588/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_35_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6851_ _7143_/CLK _6851_/D fanout587/X VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5802_ _6951_/Q _5776_/X _5786_/X _5798_/X _5801_/X VGND VGND VPWR VPWR _5802_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_90_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6782_ _6828_/CLK _6782_/D fanout583/X VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_4
X_3994_ _4152_/B _3994_/A1 _3994_/S VGND VGND VPWR VPWR _3994_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5733_ _7186_/Q _7185_/Q VGND VGND VPWR VPWR _5733_/Y sky130_fd_sc_hd__nor2_1
X_5664_ hold13/X _3474_/X _4051_/X _5665_/S hold722/X VGND VGND VPWR VPWR _5664_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_54_csclk _7277_/CLK VGND VGND VPWR VPWR _7159_/CLK sky130_fd_sc_hd__clkbuf_16
X_4615_ _4600_/B _4620_/A _4615_/C _4755_/D VGND VGND VPWR VPWR _4615_/X sky130_fd_sc_hd__and4b_1
X_5595_ _3916_/C hold521/X hold14/X VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold400 _4160_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold411 _6764_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4620_/B _5263_/A VGND VGND VPWR VPWR _4546_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold422 _6589_/Q VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _6598_/Q VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _6591_/Q VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _3366_/X VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _4098_/X VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7265_ _7265_/CLK _7265_/D fanout575/X VGND VGND VPWR VPWR _7265_/Q sky130_fd_sc_hd__dfrtp_2
X_4477_ _5042_/A _4505_/B _5042_/B _4751_/A VGND VGND VPWR VPWR _4482_/B sky130_fd_sc_hd__nand4_1
Xhold477 _4162_/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold488 _6661_/Q VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7152_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold499 hold499/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
X_6216_ _6873_/Q _6466_/A1 _5759_/A VGND VGND VPWR VPWR _6216_/X sky130_fd_sc_hd__o21a_1
X_3428_ _5548_/C _5657_/D hold27/X VGND VGND VPWR VPWR _3428_/X sky130_fd_sc_hd__and3_4
X_7196_ _7251_/CLK _7196_/D fanout594/X VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6147_ _6919_/Q _6129_/B _6129_/C _7151_/Q _6140_/X VGND VGND VPWR VPWR _6147_/X
+ sky130_fd_sc_hd__a221o_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1100 _4099_/X VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3359_ _6542_/A _3359_/B VGND VGND VPWR VPWR _3366_/S sky130_fd_sc_hd__nand2_4
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 hold1432/X VGND VGND VPWR VPWR _5612_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _5423_/X VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 _6837_/Q VGND VGND VPWR VPWR _5305_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 _6668_/Q VGND VGND VPWR VPWR _4012_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ _6772_/Q _5776_/X _6074_/X _6075_/X _6077_/X VGND VGND VPWR VPWR _6078_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold1155 _7294_/A VGND VGND VPWR VPWR _4197_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _6991_/Q VGND VGND VPWR VPWR _5486_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5029_ _5100_/B _5029_/B _5220_/B VGND VGND VPWR VPWR _5034_/A sky130_fd_sc_hd__and3_1
Xhold1177 _4203_/X VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 _4085_/X VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 _6114_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1199 _7289_/A VGND VGND VPWR VPWR _4180_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 _6177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_328 _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_339 _6606_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4400_ _5060_/C _5143_/A _5260_/B _4738_/B VGND VGND VPWR VPWR _4450_/C sky130_fd_sc_hd__nand4_1
X_5380_ hold310/X _3919_/C _5385_/S VGND VGND VPWR VPWR _5380_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4331_ _4509_/A _4584_/B _4509_/D VGND VGND VPWR VPWR _4615_/C sky130_fd_sc_hd__and3_1
XFILLER_141_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7050_ _7114_/CLK _7050_/D fanout604/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_4
X_4262_ _5036_/B _4208_/Y _4246_/Y _4356_/A _4848_/A VGND VGND VPWR VPWR _4262_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_140_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6001_ _6023_/A2 _5761_/X _6000_/X _5999_/X VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__o22a_1
XFILLER_101_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4193_ _4193_/A0 _4192_/X _4205_/S VGND VGND VPWR VPWR _4193_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6903_ _7071_/CLK _6903_/D fanout585/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfstp_2
X_6834_ _7067_/CLK _6834_/D fanout582/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfstp_2
X_6765_ _7267_/CLK _6765_/D _3291_/A VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3977_ hold765/X _6550_/A0 _3980_/S VGND VGND VPWR VPWR _3977_/X sky130_fd_sc_hd__mux2_1
X_5716_ _6800_/Q _5759_/B _7181_/Q _5715_/Y VGND VGND VPWR VPWR _5716_/X sky130_fd_sc_hd__o31a_1
X_6696_ _7053_/CLK _6696_/D fanout601/X VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _5692_/A1 hold964/X hold9/X VGND VGND VPWR VPWR _5647_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5578_ hold59/X hold2/X hold18/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__mux2_1
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold230 _6686_/Q VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold241 _5337_/X VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7317_ _7317_/A VGND VGND VPWR VPWR _7317_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold252 _5563_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4321_/Y _4322_/Y _4509_/A VGND VGND VPWR VPWR _4529_/X sky130_fd_sc_hd__a21o_1
Xhold263 _5493_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold274 hold274/A VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _5319_/X VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _5344_/X VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7248_ _7248_/CLK _7248_/D fanout580/X VGND VGND VPWR VPWR _7248_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7179_ _7218_/CLK _7179_/D fanout577/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _6115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 _6144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _6970_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_136 _7067_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_147 _6906_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _7211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _7316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3900_ _7006_/Q hold39/A _3407_/X _3433_/X _6942_/Q VGND VGND VPWR VPWR _3900_/X
+ sky130_fd_sc_hd__a32o_1
X_4880_ _4377_/X _4878_/B _4878_/C _4708_/A _4923_/C VGND VGND VPWR VPWR _4881_/B
+ sky130_fd_sc_hd__a32oi_4
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3831_ _6892_/Q _3445_/X _3496_/X _6996_/Q _3830_/X VGND VGND VPWR VPWR _3834_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3762_ _6844_/Q _5323_/S _3571_/X _6729_/Q _3761_/X VGND VGND VPWR VPWR _3766_/B
+ sky130_fd_sc_hd__a221o_1
X_6550_ _6550_/A0 hold746/X _6553_/S VGND VGND VPWR VPWR _6550_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ hold741/X _4051_/B _5502_/S VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__mux2_1
X_3693_ _3693_/A _3693_/B VGND VGND VPWR VPWR _3693_/Y sky130_fd_sc_hd__nand2_2
XFILLER_145_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6481_ _6514_/C _6481_/A2 _7255_/Q VGND VGND VPWR VPWR _6486_/C sky130_fd_sc_hd__a21bo_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5432_ _5667_/A0 _5432_/A1 hold67/X VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput302 _3349_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput313 hold1035/X VGND VGND VPWR VPWR hold1036/A sky130_fd_sc_hd__buf_12
Xoutput324 hold629/X VGND VGND VPWR VPWR hold630/A sky130_fd_sc_hd__buf_12
X_5363_ _3921_/B hold356/X _5367_/S VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__mux2_1
Xoutput335 hold706/X VGND VGND VPWR VPWR hold707/A sky130_fd_sc_hd__buf_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ _7162_/CLK _7102_/D fanout605/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_1
X_4314_ _4310_/B _4310_/C _4310_/D _4637_/A VGND VGND VPWR VPWR _4314_/X sky130_fd_sc_hd__a31o_1
X_5294_ hold119/X hold83/X _5294_/S VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7033_ _7129_/CLK _7033_/D fanout598/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_4
X_4245_ _4656_/C _4647_/C VGND VGND VPWR VPWR _4722_/A sky130_fd_sc_hd__and2_4
XFILLER_68_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4176_ _4176_/A0 _4175_/X _4188_/S VGND VGND VPWR VPWR _4176_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7239_/CLK _6817_/D fanout574/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6748_ _7265_/CLK _6748_/D fanout574/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6679_ _7244_/CLK _6679_/D fanout584/X VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout540 _6802_/Q VGND VGND VPWR VPWR _5759_/B sky130_fd_sc_hd__buf_6
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout573 fanout581/X VGND VGND VPWR VPWR fanout573/X sky130_fd_sc_hd__buf_6
Xmgmt_gpio_14_buff_inst _3340_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
Xfanout584 fanout589/X VGND VGND VPWR VPWR fanout584/X sky130_fd_sc_hd__clkbuf_16
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout595 fanout597/X VGND VGND VPWR VPWR fanout595/X sky130_fd_sc_hd__buf_6
XFILLER_59_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4030_ _3370_/B _4030_/A1 _4034_/S VGND VGND VPWR VPWR _4030_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5981_ _6778_/Q _5789_/X _5813_/X _6564_/Q VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4932_ _4510_/Y _4514_/Y _4522_/Y _5102_/B VGND VGND VPWR VPWR _4933_/C sky130_fd_sc_hd__o31a_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4863_ _4669_/X _4675_/Y _4859_/Y _4862_/Y VGND VGND VPWR VPWR _4864_/C sky130_fd_sc_hd__o211a_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6602_ _6945_/CLK _6602_/D fanout573/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_14 _3407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ hold93/A _5341_/A _5311_/C _3536_/X _6988_/Q VGND VGND VPWR VPWR _3814_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_25 _3446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 _3485_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4632_/B _4970_/D _4480_/B _4792_/X VGND VGND VPWR VPWR _5082_/A sky130_fd_sc_hd__a31oi_2
XANTENNA_47 _5377_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _3869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6533_ _6539_/A0 _6533_/A1 _6535_/S VGND VGND VPWR VPWR _6533_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_69 _5260_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ input29/X _3504_/X _3550_/X _7154_/Q _3744_/X VGND VGND VPWR VPWR _3745_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6464_ _6752_/Q _6098_/X _6447_/X _6463_/X _6440_/D VGND VGND VPWR VPWR _6464_/X
+ sky130_fd_sc_hd__a2111o_1
X_3676_ _6645_/Q _3407_/X _5325_/C _3675_/X VGND VGND VPWR VPWR _3676_/X sky130_fd_sc_hd__a31o_1
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5415_ _5413_/B _3916_/X _5421_/S hold794/X VGND VGND VPWR VPWR _5415_/X sky130_fd_sc_hd__a22o_1
X_6395_ _6685_/Q _6101_/X _6118_/X _6566_/Q _6394_/X VGND VGND VPWR VPWR _6395_/X
+ sky130_fd_sc_hd__a221o_1
X_5346_ hold69/X hold5/X _5349_/S VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__mux2_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput176 _3275_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3265_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3255_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_153_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5277_ _6540_/A0 hold647/X _5278_/S VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__mux2_1
X_7016_ _7108_/CLK _7016_/D fanout606/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfstp_1
X_4228_ _4228_/A _4228_/B _4228_/C _4228_/D VGND VGND VPWR VPWR _4230_/A sky130_fd_sc_hd__nand4_4
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4159_ _4162_/S hold988/X _3370_/X _4158_/D VGND VGND VPWR VPWR _4159_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout381 _4738_/A VGND VGND VPWR VPWR _5128_/A sky130_fd_sc_hd__buf_4
XFILLER_143_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_2
X_3530_ _6741_/Q _5327_/D _5575_/C _5575_/D VGND VGND VPWR VPWR _3530_/X sky130_fd_sc_hd__and4_1
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_2
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _3346_/D sky130_fd_sc_hd__buf_4
Xhold807 _7141_/Q VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_2
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold818 _7124_/Q VGND VGND VPWR VPWR hold818/X sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ _6673_/Q _4017_/B _4029_/B _6683_/Q _3458_/X VGND VGND VPWR VPWR _3462_/D
+ sky130_fd_sc_hd__a221o_1
Xhold829 _5660_/X VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5200_ _4732_/X _5200_/B _5200_/C _5200_/D VGND VGND VPWR VPWR _5226_/A sky130_fd_sc_hd__and4b_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3392_ hold24/X hold220/X _3393_/S VGND VGND VPWR VPWR _3392_/X sky130_fd_sc_hd__mux2_1
X_6180_ _7016_/Q _6177_/X _6176_/X _6175_/X _6179_/X VGND VGND VPWR VPWR _6181_/D
+ sky130_fd_sc_hd__a2111o_1
X_5131_ _5131_/A _5131_/B VGND VGND VPWR VPWR _5146_/B sky130_fd_sc_hd__and2_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1507 _6612_/Q VGND VGND VPWR VPWR _3946_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5062_ _4244_/Y _4423_/Y _4550_/Y _4497_/Y _4496_/Y VGND VGND VPWR VPWR _5062_/X
+ sky130_fd_sc_hd__o32a_1
Xhold1518 _6807_/Q VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _7213_/Q VGND VGND VPWR VPWR _6318_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ hold467/X _6538_/A0 _4016_/S VGND VGND VPWR VPWR _4013_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5964_ _7086_/Q _5965_/B _6009_/C _5788_/X _6998_/Q VGND VGND VPWR VPWR _5964_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4915_ _5040_/C _4535_/Y _4567_/Y _4629_/Y _4552_/Y VGND VGND VPWR VPWR _5264_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5895_ _7083_/Q _5965_/B _6009_/C _5788_/X _6995_/Q VGND VGND VPWR VPWR _5895_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4846_ _4843_/Y _5149_/C _5149_/D _4266_/Y VGND VGND VPWR VPWR _4846_/X sky130_fd_sc_hd__a31o_1
XFILLER_178_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4777_ _4777_/A _4777_/B _4777_/C VGND VGND VPWR VPWR _4779_/A sky130_fd_sc_hd__and3_1
XFILLER_193_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6516_ _7257_/Q _6514_/C _6483_/B _6515_/X VGND VGND VPWR VPWR _6516_/X sky130_fd_sc_hd__a31o_1
X_3728_ _6557_/Q _3359_/B _3723_/X _3725_/X _3727_/X VGND VGND VPWR VPWR _3728_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6447_ _6647_/Q _6444_/C wire392/A _6445_/X VGND VGND VPWR VPWR _6447_/X sky130_fd_sc_hd__a31o_1
X_3659_ _6675_/Q _4158_/D _4139_/C _3954_/B _6622_/Q VGND VGND VPWR VPWR _3659_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6378_ _6644_/Q _6444_/C wire392/A _6137_/X _7271_/Q VGND VGND VPWR VPWR _6378_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5329_ hold89/X hold108/X _5330_/S VGND VGND VPWR VPWR _5329_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4700_ _4708_/A _4923_/C VGND VGND VPWR VPWR _4700_/Y sky130_fd_sc_hd__nand2_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ hold13/X _3509_/X _3924_/X _5683_/S hold563/X VGND VGND VPWR VPWR _5680_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _4718_/D _4687_/B VGND VGND VPWR VPWR _4688_/C sky130_fd_sc_hd__nand2_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4562_ _4562_/A _4562_/B _4562_/C _4562_/D VGND VGND VPWR VPWR _4565_/A sky130_fd_sc_hd__nor4_1
XFILLER_162_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6301_ _7125_/Q _6176_/B _6446_/C _6129_/D _6909_/Q VGND VGND VPWR VPWR _6301_/X
+ sky130_fd_sc_hd__a32o_1
Xhold604 _5435_/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 _7268_/Q VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _6524_/A _4127_/C _4158_/D VGND VGND VPWR VPWR _3513_/X sky130_fd_sc_hd__and3_4
X_7281_ _7281_/A VGND VGND VPWR VPWR _7281_/X sky130_fd_sc_hd__clkbuf_2
Xhold626 _5351_/X VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4493_ _4493_/A _4843_/A _4493_/C VGND VGND VPWR VPWR _4504_/A sky130_fd_sc_hd__nor3_1
Xhold637 hold637/A VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _5277_/X VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold659 _5480_/X VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6232_ _6986_/Q _6098_/X _6112_/X _7106_/Q _6231_/X VGND VGND VPWR VPWR _6239_/A
+ sky130_fd_sc_hd__a221o_1
X_3444_ _5304_/A _6530_/D _5666_/C VGND VGND VPWR VPWR _4092_/S sky130_fd_sc_hd__and3_4
Xmax_cap389 _6105_/X VGND VGND VPWR VPWR _6129_/C sky130_fd_sc_hd__buf_12
X_3375_ _3919_/C hold334/X _3377_/S VGND VGND VPWR VPWR _3375_/X sky130_fd_sc_hd__mux2_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _7055_/Q _6136_/A _6465_/A3 _6145_/X _7007_/Q VGND VGND VPWR VPWR _6163_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5255_/A _4683_/X _5110_/X _4872_/B VGND VGND VPWR VPWR _5257_/C sky130_fd_sc_hd__a31oi_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1304 _3978_/X VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6094_ _6136_/A _6347_/C _6177_/C VGND VGND VPWR VPWR _6129_/A sky130_fd_sc_hd__and3_4
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 _6895_/Q VGND VGND VPWR VPWR hold724/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _6736_/Q VGND VGND VPWR VPWR hold439/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 _5668_/X VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1348 _4026_/X VGND VGND VPWR VPWR _6680_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5045_ _4376_/Y _4391_/Y _4423_/Y _5044_/Y _4827_/C VGND VGND VPWR VPWR _5142_/D
+ sky130_fd_sc_hd__o311a_1
Xhold1359 _5676_/X VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6996_ _7171_/CLK _6996_/D fanout611/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5947_ _7117_/Q _5826_/B _5842_/C _5946_/X VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__a31o_1
XFILLER_179_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5878_ _6930_/Q _5970_/B1 _5815_/X _7018_/Q _5877_/X VGND VGND VPWR VPWR _5878_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4829_ _4829_/A _4829_/B _4829_/C _4829_/D VGND VGND VPWR VPWR _4829_/X sky130_fd_sc_hd__and4_1
XFILLER_193_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6850_ _7263_/CLK _6850_/D fanout578/X VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5801_ _7071_/Q _5971_/A2 _5782_/X _6935_/Q _5800_/X VGND VGND VPWR VPWR _5801_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6781_ _6781_/CLK _6781_/D fanout575/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtp_4
X_3993_ _5304_/A _6536_/B _5630_/C _4158_/D VGND VGND VPWR VPWR _3994_/S sky130_fd_sc_hd__nand4_4
XFILLER_22_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5732_ _7186_/Q _7185_/Q VGND VGND VPWR VPWR _5732_/X sky130_fd_sc_hd__and2_2
XFILLER_50_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5663_ hold83/X hold192/X _5665_/S VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4614_ _4620_/A _4595_/A _5263_/B _4333_/A _4939_/A VGND VGND VPWR VPWR _5216_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_163_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5594_ _5667_/A0 hold966/X hold14/X VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold401 hold401/A VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4545_ _4540_/Y _4541_/Y _4544_/Y VGND VGND VPWR VPWR _4554_/A sky130_fd_sc_hd__o21a_1
Xhold412 _4141_/X VGND VGND VPWR VPWR _6764_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold423 _3910_/X VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _3929_/X VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold445 _3912_/X VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7264_ _7264_/CLK _7264_/D fanout580/X VGND VGND VPWR VPWR _7264_/Q sky130_fd_sc_hd__dfrtp_4
Xhold456 _6826_/Q VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4476_/A _4476_/B _4476_/C VGND VGND VPWR VPWR _4482_/A sky130_fd_sc_hd__nor3_1
XFILLER_131_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold467 _6669_/Q VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _6679_/Q VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _4003_/X VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6196_/X _6215_/B _6215_/C VGND VGND VPWR VPWR _6215_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3427_ hold54/X hold16/X hold75/X _5324_/B VGND VGND VPWR VPWR _3427_/Y sky130_fd_sc_hd__o31ai_4
X_7195_ _7219_/CLK _7195_/D fanout595/X VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6146_ _7087_/Q _6136_/A _6106_/C _6129_/A _6895_/Q VGND VGND VPWR VPWR _6146_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _6524_/A _5476_/B _6536_/A VGND VGND VPWR VPWR _3359_/B sky130_fd_sc_hd__and3_4
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1101 _6862_/Q VGND VGND VPWR VPWR _5340_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1112 hold1330/X VGND VGND VPWR VPWR _5560_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 hold1447/X VGND VGND VPWR VPWR _5513_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _5305_/X VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6077_ _7264_/Q _5777_/X _5779_/X _6777_/Q _6076_/X VGND VGND VPWR VPWR _6077_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1145 _4012_/X VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3289_ _4656_/C VGND VGND VPWR VPWR _4691_/B sky130_fd_sc_hd__inv_4
Xhold1156 _4197_/X VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _5486_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1178 _7292_/A VGND VGND VPWR VPWR _4193_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5028_ _4473_/Y _4514_/Y _4601_/Y _4525_/Y VGND VGND VPWR VPWR _5220_/B sky130_fd_sc_hd__a31o_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _7167_/Q VGND VGND VPWR VPWR _5685_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _6114_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_318 _6177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 _7017_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6979_ _7063_/CLK _6979_/D fanout590/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold990 _7017_/Q VGND VGND VPWR VPWR hold990/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4330_ _4320_/B _4940_/C _4691_/B _4523_/A VGND VGND VPWR VPWR _4584_/B sky130_fd_sc_hd__o211a_2
XFILLER_181_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4261_ _4632_/B _4600_/B _4612_/C _4647_/C _4848_/A VGND VGND VPWR VPWR _4295_/A
+ sky130_fd_sc_hd__a41oi_4
X_6000_ _6442_/S _7201_/Q _6443_/S VGND VGND VPWR VPWR _6000_/X sky130_fd_sc_hd__a21o_1
X_4192_ hold613/X _3915_/X _4204_/S VGND VGND VPWR VPWR _4192_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6902_ _7006_/CLK _6902_/D fanout601/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6833_ _6835_/CLK hold74/X fanout583/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6764_ _7241_/CLK _6764_/D fanout576/X VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_2
X_3976_ hold897/X _6543_/A0 _3980_/S VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5715_ _7181_/Q _7180_/Q _5759_/B VGND VGND VPWR VPWR _5715_/Y sky130_fd_sc_hd__o21ai_1
X_6695_ _7006_/CLK _6695_/D fanout601/X VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5646_ hold21/X hold182/X hold9/X VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ hold671/X _6550_/A0 hold18/X VGND VGND VPWR VPWR _5577_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold220 _6572_/Q VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_7316_ _7316_/A VGND VGND VPWR VPWR _7316_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold231 _4033_/X VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4528_ _4280_/B _4301_/Y _4320_/Y _4657_/C _4509_/D VGND VGND VPWR VPWR _4561_/B
+ sky130_fd_sc_hd__o221a_4
Xhold242 _6877_/Q VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold264 _6878_/Q VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7247_ _7263_/CLK _7247_/D fanout578/X VGND VGND VPWR VPWR _7247_/Q sky130_fd_sc_hd__dfrtp_4
Xhold275 _7168_/Q VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4459_ _4459_/A _4459_/B _4459_/C VGND VGND VPWR VPWR _4461_/C sky130_fd_sc_hd__nand3_1
Xhold286 _7164_/Q VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _7102_/Q VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7178_ _7218_/CLK _7178_/D fanout594/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _6129_/A _6129_/B _6129_/C _6129_/D VGND VGND VPWR VPWR _6132_/B sky130_fd_sc_hd__nor4_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _6115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _6147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _6970_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 _7067_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _6922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _7193_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7031_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _6980_/Q _5485_/B _5684_/C _3525_/X _7124_/Q VGND VGND VPWR VPWR _3830_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7077_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3761_ _6883_/Q _5359_/B _3544_/X _6947_/Q VGND VGND VPWR VPWR _3761_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5500_ hold113/X hold83/X _5502_/S VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6480_ _3905_/Y _6480_/A1 _6480_/S VGND VGND VPWR VPWR _7228_/D sky130_fd_sc_hd__mux2_1
X_3692_ _3692_/A _3692_/B _3692_/C _3692_/D VGND VGND VPWR VPWR _3692_/Y sky130_fd_sc_hd__nor4_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5431_ hold66/A _5494_/C _5575_/C _5575_/D VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__nand4_4
Xoutput303 _3307_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput314 hold637/X VGND VGND VPWR VPWR hold638/A sky130_fd_sc_hd__buf_12
X_5362_ _5359_/B _3919_/X _5367_/S _5362_/B2 VGND VGND VPWR VPWR _5362_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput325 hold633/X VGND VGND VPWR VPWR hold634/A sky130_fd_sc_hd__buf_12
Xoutput336 hold593/X VGND VGND VPWR VPWR hold594/A sky130_fd_sc_hd__buf_12
X_7101_ _7161_/CLK _7101_/D fanout599/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfrtp_1
X_4313_ _4313_/A _4637_/A VGND VGND VPWR VPWR _4313_/Y sky130_fd_sc_hd__nand2_1
X_5293_ hold954/X _6535_/A0 _5294_/S VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7032_ _7088_/CLK _7032_/D fanout590/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4244_ _4760_/C _4488_/B VGND VGND VPWR VPWR _4244_/Y sky130_fd_sc_hd__nand2_2
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4175_ hold360/X _3915_/X _4187_/S VGND VGND VPWR VPWR _4175_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6816_ _6827_/CLK _6816_/D fanout575/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6747_ _7269_/CLK _6747_/D fanout576/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3959_ _3925_/C hold402/X _3959_/S VGND VGND VPWR VPWR _3959_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6678_ _6827_/CLK _6678_/D fanout573/X VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5629_ hold8/X _6548_/A _5629_/C VGND VGND VPWR VPWR _5637_/S sky130_fd_sc_hd__and3_2
XFILLER_152_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout530 hold89/X VGND VGND VPWR VPWR _6550_/A0 sky130_fd_sc_hd__clkbuf_16
Xfanout541 _6292_/S VGND VGND VPWR VPWR _6442_/S sky130_fd_sc_hd__buf_6
XFILLER_76_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout563 _4675_/A VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__buf_6
Xfanout574 fanout575/X VGND VGND VPWR VPWR fanout574/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout585 fanout589/X VGND VGND VPWR VPWR fanout585/X sky130_fd_sc_hd__buf_8
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout596 fanout597/X VGND VGND VPWR VPWR fanout596/X sky130_fd_sc_hd__buf_8
XFILLER_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5980_ _6597_/Q _6025_/B _6028_/B _5777_/X _7260_/Q VGND VGND VPWR VPWR _5980_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_64_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4931_ _4786_/B _4600_/Y _4603_/B VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4862_ _4862_/A _4862_/B VGND VGND VPWR VPWR _4862_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6601_ _6751_/CLK _6601_/D fanout572/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfrtp_4
X_3813_ _3965_/A0 _3813_/A1 _3906_/S VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 _3412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _5611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4799_/B _4712_/B _4792_/C _4791_/X VGND VGND VPWR VPWR _4793_/X sky130_fd_sc_hd__a31o_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _6550_/A0 hold684/X _6535_/S VGND VGND VPWR VPWR _6532_/X sky130_fd_sc_hd__mux2_1
X_3744_ _6938_/Q hold39/A _5422_/D _3559_/X _6906_/Q VGND VGND VPWR VPWR _3744_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_59 _3875_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6463_ _7243_/Q _6115_/X _6119_/X _6591_/Q _6462_/X VGND VGND VPWR VPWR _6463_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3675_ _7017_/Q _5512_/B _3412_/X _3562_/X _6640_/Q VGND VGND VPWR VPWR _3675_/X
+ sky130_fd_sc_hd__a32o_1
X_5414_ _6549_/A0 _5414_/A1 _5421_/S VGND VGND VPWR VPWR _5414_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6394_ _6576_/Q _6444_/B _6465_/A2 _6454_/B1 _6770_/Q VGND VGND VPWR VPWR _6394_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_126_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5345_ hold121/X _3922_/C _5349_/S VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput177 _3274_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3264_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
XFILLER_142_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput199 _3254_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
X_5276_ _6539_/A0 _5276_/A1 _5278_/S VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7015_ _7015_/CLK _7015_/D fanout588/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfstp_2
X_4227_ _4227_/A _4227_/B _4227_/C _4227_/D VGND VGND VPWR VPWR _4235_/A sky130_fd_sc_hd__nand4_4
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ _6542_/A _5476_/B _6536_/C _4158_/D VGND VGND VPWR VPWR _4162_/S sky130_fd_sc_hd__nand4_4
XFILLER_110_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4089_ _4089_/A0 _4088_/X _4093_/S VGND VGND VPWR VPWR _4089_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_1
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _3349_/B sky130_fd_sc_hd__buf_2
Xhold808 _5655_/X VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput79 spi_enabled VGND VGND VPWR VPWR _3350_/A sky130_fd_sc_hd__buf_6
XFILLER_116_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold819 _5636_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3460_ _6536_/C _6530_/D _5327_/D VGND VGND VPWR VPWR _4029_/B sky130_fd_sc_hd__and3_4
XFILLER_115_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3391_ _3918_/B hold435/X _3393_/S VGND VGND VPWR VPWR _3391_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5130_ _5129_/X _4729_/X _5127_/Y _4981_/X VGND VGND VPWR VPWR _5130_/X sky130_fd_sc_hd__o31a_1
XFILLER_123_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1508 _7256_/Q VGND VGND VPWR VPWR _7253_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5061_ _5061_/A _5235_/C _5061_/C _5234_/A VGND VGND VPWR VPWR _5061_/X sky130_fd_sc_hd__and4_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1519 _7210_/Q VGND VGND VPWR VPWR _6243_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4012_ _4012_/A0 _3370_/B _4016_/S VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5963_ _6886_/Q _5768_/X _5794_/X _6926_/Q _5962_/X VGND VGND VPWR VPWR _5963_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4914_ _4899_/X _4914_/B _5174_/D _5265_/A VGND VGND VPWR VPWR _4916_/B sky130_fd_sc_hd__and4b_1
XFILLER_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5894_ _6963_/Q _5770_/X _5793_/X _6987_/Q _5893_/X VGND VGND VPWR VPWR _5894_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_33_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4845_ _4859_/C _4597_/C _5143_/D _5060_/B _5060_/A VGND VGND VPWR VPWR _5149_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4776_ _4776_/A _4776_/B _4776_/C VGND VGND VPWR VPWR _4779_/C sky130_fd_sc_hd__nand3_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6515_ _7258_/Q _6514_/C _6482_/B _6514_/X VGND VGND VPWR VPWR _6515_/X sky130_fd_sc_hd__a31o_1
X_3727_ _7114_/Q _3463_/X _5359_/B _6882_/Q _3726_/X VGND VGND VPWR VPWR _3727_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6446_ _6563_/Q _6446_/B _6446_/C VGND VGND VPWR VPWR _6446_/X sky130_fd_sc_hd__and3_1
X_3658_ _6775_/Q _3533_/C _5325_/C _3536_/X _6985_/Q VGND VGND VPWR VPWR _3658_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6377_ _6575_/Q _6104_/X _6130_/X _6779_/Q _6376_/X VGND VGND VPWR VPWR _6380_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3589_ _6888_/Q _5440_/C _3533_/C _3474_/X _7144_/Q VGND VGND VPWR VPWR _3589_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5328_ _3918_/B hold512/X _5330_/S VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5259_ _5128_/B _5140_/C _5060_/C _5143_/A _5260_/B VGND VGND VPWR VPWR _5259_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4630_ _4984_/B _4984_/C _5263_/C VGND VGND VPWR VPWR _4687_/B sky130_fd_sc_hd__and3_1
XFILLER_187_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4561_ _4751_/A _4561_/B _4581_/B VGND VGND VPWR VPWR _4562_/C sky130_fd_sc_hd__and3_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6300_ _6917_/Q _6451_/B1 _6136_/X _7029_/Q _6299_/X VGND VGND VPWR VPWR _6305_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3512_ _6554_/Q _3359_/B _3397_/B _6574_/Q _3511_/X VGND VGND VPWR VPWR _3523_/A
+ sky130_fd_sc_hd__a221o_1
Xhold605 _7247_/Q VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _6540_/X VGND VGND VPWR VPWR _7268_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _5060_/A _5060_/B _5055_/D _4557_/B VGND VGND VPWR VPWR _4843_/B sky130_fd_sc_hd__and4_1
XFILLER_171_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold627 _7105_/Q VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold649 hold649/A VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _7010_/Q _6444_/C _6096_/Y _6325_/A2 _6882_/Q VGND VGND VPWR VPWR _6231_/X
+ sky130_fd_sc_hd__a32o_1
X_3443_ _6733_/Q _3441_/X _3442_/X _6638_/Q _3440_/X VGND VGND VPWR VPWR _3462_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6911_/Q _6451_/B1 _6122_/X _6887_/Q _6161_/X VGND VGND VPWR VPWR _6165_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ hold89/X hold134/X _3377_/S VGND VGND VPWR VPWR _3374_/X sky130_fd_sc_hd__mux2_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _4675_/A _4862_/A _4732_/C _4989_/X _5112_/X VGND VGND VPWR VPWR _5231_/B
+ sky130_fd_sc_hd__a311oi_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6143_/D _7187_/Q VGND VGND VPWR VPWR _6145_/C sky130_fd_sc_hd__nor2_4
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 _7128_/Q VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _6912_/Q VGND VGND VPWR VPWR hold398/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 _4107_/X VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B VGND VGND VPWR VPWR _5044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1338 _7080_/Q VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 _7095_/Q VGND VGND VPWR VPWR hold1349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6995_ _7108_/CLK _6995_/D fanout606/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5946_ _7077_/Q _5971_/A2 _5813_/X _7061_/Q _5945_/X VGND VGND VPWR VPWR _5946_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5877_ _7090_/Q _5826_/B wire398/X _5788_/X _6994_/Q VGND VGND VPWR VPWR _5877_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4828_ _4738_/B _4597_/C _5140_/B _5055_/D _5143_/A VGND VGND VPWR VPWR _4829_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4759_ _4749_/X _4752_/Y _4758_/Y VGND VGND VPWR VPWR _4765_/A sky130_fd_sc_hd__a21oi_1
XFILLER_181_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6429_ _6646_/Q _6177_/C _6112_/C _6462_/B1 _6656_/Q VGND VGND VPWR VPWR _6429_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__buf_12
XFILLER_82_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5800_ _6903_/Q _5934_/C _6003_/C _5799_/X VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6780_ _6780_/CLK _6780_/D fanout575/X VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfstp_2
X_3992_ _3924_/B hold575/X _3992_/S VGND VGND VPWR VPWR _3992_/X sky130_fd_sc_hd__mux2_1
X_5731_ _5752_/B2 _7185_/Q _5730_/Y VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__a21oi_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5662_ hold13/X _3474_/X _3924_/X _5665_/S hold777/X VGND VGND VPWR VPWR _5662_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4613_ _4789_/B _4755_/D VGND VGND VPWR VPWR _4613_/Y sky130_fd_sc_hd__nand2_4
XFILLER_191_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5593_ hold13/X _5593_/B VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__nand2_8
XFILLER_190_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4544_ _4544_/A _4544_/B _4544_/C _4544_/D VGND VGND VPWR VPWR _4544_/Y sky130_fd_sc_hd__nand4_1
Xhold402 _6624_/Q VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _6856_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold424 _6979_/Q VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7263_ _7263_/CLK _7263_/D fanout578/X VGND VGND VPWR VPWR _7263_/Q sky130_fd_sc_hd__dfrtp_4
Xhold435 _6571_/Q VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _6608_/Q VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4505_/B _4475_/B _4597_/C VGND VGND VPWR VPWR _4476_/B sky130_fd_sc_hd__and3_1
Xhold457 _5292_/X VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold468 _4013_/X VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6214_ _6214_/A _6214_/B _6440_/D _6214_/D VGND VGND VPWR VPWR _6214_/Y sky130_fd_sc_hd__nor4_1
Xhold479 _4025_/X VGND VGND VPWR VPWR _6679_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ hold54/X hold16/X hold75/X VGND VGND VPWR VPWR _3757_/D sky130_fd_sc_hd__nor3_4
X_7194_ _7219_/CLK _7194_/D fanout578/X VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6145_ _6444_/C _6425_/B _6145_/C VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__and3_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3357_ hold16/X hold75/X _5324_/B hold54/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__and4b_4
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _5340_/X VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _6653_/Q VGND VGND VPWR VPWR _3994_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _6903_/Q VGND VGND VPWR VPWR _5387_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_6076_ _6563_/Q _6072_/B _6025_/C _5767_/X _6558_/Q VGND VGND VPWR VPWR _6076_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1135 _6959_/Q VGND VGND VPWR VPWR _5450_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3288_ _4657_/C VGND VGND VPWR VPWR _4870_/B sky130_fd_sc_hd__clkinv_8
Xhold1146 _6816_/Q VGND VGND VPWR VPWR _5280_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1157 _6620_/Q VGND VGND VPWR VPWR _3955_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5027_ _5027_/A _5027_/B _5177_/B VGND VGND VPWR VPWR _5029_/B sky130_fd_sc_hd__nor3_1
Xhold1168 hold1393/X VGND VGND VPWR VPWR _5477_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1179 _4193_/X VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 _6115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_319 _6184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6978_ _7165_/CLK _6978_/D fanout601/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfrtp_4
X_5929_ _6010_/C _5910_/X _5921_/X _5925_/X _5928_/X VGND VGND VPWR VPWR _5929_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold980 _7286_/A VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold991 _5515_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4260_ _4632_/B _4600_/B _4612_/C _4647_/C VGND VGND VPWR VPWR _4356_/A sky130_fd_sc_hd__a31o_4
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4191_ _4191_/A0 _4190_/X _4205_/S VGND VGND VPWR VPWR _4191_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6901_ _6957_/CLK _6901_/D fanout591/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6832_ _6855_/CLK _6832_/D fanout583/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_63_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6763_ _6827_/CLK _6763_/D fanout573/X VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfrtp_2
X_3975_ _6524_/A _6524_/B _6530_/C _6536_/D VGND VGND VPWR VPWR _3980_/S sky130_fd_sc_hd__and4_4
X_5714_ _7181_/Q _7180_/Q VGND VGND VPWR VPWR _5714_/Y sky130_fd_sc_hd__nor2_2
XFILLER_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6694_ _7157_/CLK _6694_/D fanout592/X VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5645_ _6505_/A1 hold842/X hold9/X VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5576_ _5576_/A0 _5649_/A0 hold18/X VGND VGND VPWR VPWR _5576_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold210 _5484_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7315_ _7315_/A VGND VGND VPWR VPWR _7315_/X sky130_fd_sc_hd__buf_2
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold221 _3392_/X VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _4523_/C _4523_/A _4336_/X _4522_/Y VGND VGND VPWR VPWR _4527_/X sky130_fd_sc_hd__a211o_2
XFILLER_2_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold232 _6962_/Q VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _5357_/X VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _6995_/Q VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _5358_/X VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7246_ _7273_/CLK _7246_/D fanout579/X VGND VGND VPWR VPWR _7246_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_131_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4458_ _4860_/C _4457_/X _4396_/X _4456_/Y VGND VGND VPWR VPWR _4459_/A sky130_fd_sc_hd__a211oi_1
Xhold276 _5686_/X VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold287 _5681_/X VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold298 _5610_/X VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ hold16/X hold75/X _5324_/B hold54/X VGND VGND VPWR VPWR _3409_/X sky130_fd_sc_hd__and4bb_2
X_7177_ _7218_/CLK _7177_/D fanout577/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4389_ _5143_/A _5260_/B _4738_/B _5143_/D VGND VGND VPWR VPWR _4459_/C sky130_fd_sc_hd__nand4_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _6130_/A _6138_/B _6143_/C VGND VGND VPWR VPWR _6129_/D sky130_fd_sc_hd__and3_4
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6059_ _6771_/Q _6651_/Q _6059_/S VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__mux2_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _6130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_116 _6181_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 hold61/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _7067_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _6779_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ _6762_/Q _4133_/B _4017_/B _6677_/Q _3759_/X VGND VGND VPWR VPWR _3766_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3691_ _6945_/Q _3544_/X _3686_/X _3688_/X _3690_/X VGND VGND VPWR VPWR _3692_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5430_ _4053_/B hold214/X _5430_/S VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput304 _3344_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
X_5361_ _5359_/B _3916_/X _5367_/S hold921/X VGND VGND VPWR VPWR _5361_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput315 hold519/X VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__buf_12
Xoutput326 hold700/X VGND VGND VPWR VPWR hold701/A sky130_fd_sc_hd__buf_12
XFILLER_126_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput337 hold725/X VGND VGND VPWR VPWR hold726/A sky130_fd_sc_hd__buf_12
X_7100_ _7117_/CLK _7100_/D fanout605/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_2
X_4312_ _4312_/A _4544_/D VGND VGND VPWR VPWR _4517_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5292_ hold456/X _6546_/A0 _5294_/S VGND VGND VPWR VPWR _5292_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7031_ _7031_/CLK _7031_/D fanout599/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4243_ _4243_/A _4243_/B _4760_/C VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__and3_4
XFILLER_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4174_ _4174_/A0 _4173_/X _4188_/S VGND VGND VPWR VPWR _4174_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6815_ _7275_/CLK _6815_/D fanout596/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6746_ _7278_/CLK _6746_/D fanout595/X VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfrtp_4
X_3958_ _6540_/A0 hold688/X _3959_/S VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6677_ _6843_/CLK _6677_/D fanout584/X VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfrtp_1
X_3889_ _3889_/A _3889_/B _3889_/C _3889_/D VGND VGND VPWR VPWR _3889_/Y sky130_fd_sc_hd__nor4_1
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5628_ _6511_/A1 hold290/X _5628_/S VGND VGND VPWR VPWR _5628_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5559_ _3915_/B hold309/X _5565_/S VGND VGND VPWR VPWR _5559_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7229_ _3340_/A1 _7229_/D fanout613/X VGND VGND VPWR VPWR _7229_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout520 _3922_/C VGND VGND VPWR VPWR _6540_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout531 hold89/X VGND VGND VPWR VPWR _3915_/B sky130_fd_sc_hd__buf_4
Xfanout542 _6801_/Q VGND VGND VPWR VPWR _6292_/S sky130_fd_sc_hd__buf_8
XFILLER_59_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout575 fanout581/X VGND VGND VPWR VPWR fanout575/X sky130_fd_sc_hd__buf_8
XFILLER_76_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout586 fanout589/X VGND VGND VPWR VPWR fanout586/X sky130_fd_sc_hd__buf_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout597 fanout598/X VGND VGND VPWR VPWR fanout597/X sky130_fd_sc_hd__buf_6
XFILLER_100_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4930_ _4595_/A _4774_/B _4596_/B VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4861_ _4860_/X _4654_/B _4409_/C _4668_/C _4674_/X VGND VGND VPWR VPWR _4862_/B
+ sky130_fd_sc_hd__a41o_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6600_ _7264_/CLK _6600_/D fanout579/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfrtp_4
X_3812_ _6682_/Q _3553_/X _3758_/X _3811_/Y VGND VGND VPWR VPWR _3812_/X sky130_fd_sc_hd__a211o_2
XANTENNA_16 _3414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4792_ _4792_/A _4792_/B _4792_/C VGND VGND VPWR VPWR _4792_/X sky130_fd_sc_hd__and3_1
XFILLER_177_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_27 _5611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6531_ _6543_/A0 hold890/X _6535_/S VGND VGND VPWR VPWR _6531_/X sky130_fd_sc_hd__mux2_1
X_3743_ _6841_/Q _5666_/C hold39/A _3503_/X _7138_/Q VGND VGND VPWR VPWR _3743_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_49 _3544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6462_ _6642_/Q _6177_/C _6110_/C _6462_/B1 _6657_/Q VGND VGND VPWR VPWR _6462_/X
+ sky130_fd_sc_hd__a32o_1
X_3674_ _7246_/Q _6530_/C _5341_/A _3673_/X VGND VGND VPWR VPWR _3674_/X sky130_fd_sc_hd__a31o_1
X_5413_ hold13/X _5413_/B VGND VGND VPWR VPWR _5421_/S sky130_fd_sc_hd__nand2_8
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6393_ _6392_/X _6393_/A1 _6443_/S VGND VGND VPWR VPWR _7216_/D sky130_fd_sc_hd__mux2_1
X_5344_ hold295/X _3919_/C _5349_/S VGND VGND VPWR VPWR _5344_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput178 _3273_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3263_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ hold89/X hold138/X _5278_/S VGND VGND VPWR VPWR _5275_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4226_ _4227_/A _4227_/B _4227_/C _4227_/D VGND VGND VPWR VPWR _4284_/C sky130_fd_sc_hd__and4_4
X_7014_ _7173_/CLK _7014_/D fanout602/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4157_ _4152_/C _3925_/X _4156_/S hold899/X VGND VGND VPWR VPWR _4157_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4088_ hold102/X _4049_/X _4092_/S VGND VGND VPWR VPWR _4088_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6729_ _6835_/CLK _6729_/D fanout583/X VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_52_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7161_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_67_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7143_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _3351_/B sky130_fd_sc_hd__buf_2
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_4
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold809 _7139_/Q VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_108_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3390_ _6550_/A0 hold763/X _3393_/S VGND VGND VPWR VPWR _3390_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5060_ _5060_/A _5060_/B _5060_/C _5140_/C VGND VGND VPWR VPWR _5235_/C sky130_fd_sc_hd__nand4_1
XFILLER_69_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 _7281_/A VGND VGND VPWR VPWR _5314_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4011_ _6524_/A _6536_/B _4127_/C _4158_/D VGND VGND VPWR VPWR _4016_/S sky130_fd_sc_hd__and4_2
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5962_ _6966_/Q _5770_/X _5793_/X _6990_/Q _5961_/X VGND VGND VPWR VPWR _5962_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4913_ _5040_/C _4527_/X _4529_/X _4552_/Y _4635_/Y VGND VGND VPWR VPWR _5265_/A
+ sky130_fd_sc_hd__o32a_1
X_5893_ _6979_/Q _6073_/B2 _5774_/X _6907_/Q _5892_/X VGND VGND VPWR VPWR _5893_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4844_ _4319_/X _4423_/Y _4490_/Y _4497_/Y _4388_/Y VGND VGND VPWR VPWR _5149_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ _4778_/C _4775_/B VGND VGND VPWR VPWR _4776_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6514_ _7259_/Q _6514_/B _6514_/C VGND VGND VPWR VPWR _6514_/X sky130_fd_sc_hd__and3_1
X_3726_ _7278_/Q _6536_/A _3466_/X _3954_/B _6623_/Q VGND VGND VPWR VPWR _3726_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6445_ _7269_/Q _6136_/A _6106_/C _6107_/X _6815_/Q VGND VGND VPWR VPWR _6445_/X
+ sky130_fd_sc_hd__a32o_1
X_3657_ _7025_/Q _3563_/X _3654_/X _3655_/X _3656_/X VGND VGND VPWR VPWR _3657_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_106_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3588_ _6824_/Q _3497_/X _3571_/X _6726_/Q _3574_/X VGND VGND VPWR VPWR _3588_/X
+ sky130_fd_sc_hd__a221o_1
X_6376_ _6598_/Q _6444_/C _6465_/A3 _6116_/X _6570_/Q VGND VGND VPWR VPWR _6376_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5327_ _5476_/B _6536_/B _6536_/C _5327_/D VGND VGND VPWR VPWR _5330_/S sky130_fd_sc_hd__nand4_4
XFILLER_88_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5258_ _5258_/A _5258_/B _5258_/C _5258_/D VGND VGND VPWR VPWR _5258_/X sky130_fd_sc_hd__and4_1
X_4209_ _4511_/A _4632_/C _4729_/A VGND VGND VPWR VPWR _4209_/Y sky130_fd_sc_hd__nand3_4
X_5189_ _4244_/Y _4423_/Y _4550_/Y _4497_/Y _4299_/Y VGND VGND VPWR VPWR _5189_/Y
+ sky130_fd_sc_hd__o32ai_1
XFILLER_56_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4560_ _4560_/A _4560_/B _4560_/C VGND VGND VPWR VPWR _4562_/D sky130_fd_sc_hd__nand3_1
XFILLER_190_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3511_ _7159_/Q _3509_/X _3510_/X _7095_/Q VGND VGND VPWR VPWR _3511_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold606 _6528_/X VGND VGND VPWR VPWR _7247_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _5060_/A _5060_/B _5055_/D _5140_/C _4488_/X VGND VGND VPWR VPWR _4493_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_7_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold617 hold617/A VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _5614_/X VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3442_ _6524_/A _6530_/C _6536_/D VGND VGND VPWR VPWR _3442_/X sky130_fd_sc_hd__and3_1
Xhold639 _6771_/Q VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6230_/A _6230_/B _6230_/C _6230_/D VGND VGND VPWR VPWR _6230_/Y sky130_fd_sc_hd__nor4_1
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3373_ _3373_/A1 _3377_/S _3370_/X _6536_/A VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__a22o_1
X_6161_ _6879_/Q _6325_/A2 _6454_/B1 _6951_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5255_/A _4738_/B _4857_/C _4850_/X VGND VGND VPWR VPWR _5112_/X sky130_fd_sc_hd__a31o_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _7189_/Q _7190_/Q VGND VGND VPWR VPWR _6092_/Y sky130_fd_sc_hd__nor2_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1306 _5641_/X VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 _5397_/X VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5043_ _5143_/A _5143_/C _5260_/A _5060_/B VGND VGND VPWR VPWR _5058_/C sky130_fd_sc_hd__nand4_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1328 _6820_/Q VGND VGND VPWR VPWR hold971/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 _5586_/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wbbd_sck _7237_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6994_ _7145_/CLK _6994_/D fanout602/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5945_ _7045_/Q _5826_/B _5959_/B _5970_/B1 _6933_/Q VGND VGND VPWR VPWR _5945_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5876_ _6882_/Q _5768_/X _5783_/X _7010_/Q _5875_/X VGND VGND VPWR VPWR _5876_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4827_ _4827_/A _4827_/B _4827_/C _4827_/D VGND VGND VPWR VPWR _4829_/C sky130_fd_sc_hd__and4_1
XFILLER_178_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4758_ _4648_/Y _4745_/Y _4755_/Y _4756_/Y VGND VGND VPWR VPWR _4758_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3709_ _6954_/Q _3424_/X _3482_/X _6771_/Q _3708_/X VGND VGND VPWR VPWR _3717_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4689_ _4689_/A _4689_/B _4689_/C VGND VGND VPWR VPWR _4689_/X sky130_fd_sc_hd__and3_1
XFILLER_107_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6428_ _6600_/Q _6109_/X _6115_/X _7242_/Q _6427_/X VGND VGND VPWR VPWR _6431_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6359_ _6620_/Q _6136_/X _6177_/X _6638_/Q VGND VGND VPWR VPWR _6359_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_82_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3991_ hold24/X hold202/X _3992_/S VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5730_ _6800_/Q _5759_/B _7185_/Q VGND VGND VPWR VPWR _5730_/Y sky130_fd_sc_hd__nor3_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5661_ hold13/X _3474_/X _3921_/X _5665_/S hold748/X VGND VGND VPWR VPWR _5661_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4612_ _4511_/A _4600_/B _4612_/C _4632_/A VGND VGND VPWR VPWR _5263_/B sky130_fd_sc_hd__and4bb_4
X_5592_ _5692_/A1 hold913/X hold44/X VGND VGND VPWR VPWR _5592_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4543_ _4600_/B _4848_/A _4801_/A _4674_/D VGND VGND VPWR VPWR _4544_/C sky130_fd_sc_hd__and4b_1
XFILLER_190_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold403 _3959_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _5333_/X VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _5472_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7262_ _7273_/CLK _7262_/D fanout579/X VGND VGND VPWR VPWR _7262_/Q sky130_fd_sc_hd__dfstp_1
Xhold436 _3391_/X VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _4633_/B _4689_/B _4511_/A VGND VGND VPWR VPWR _4474_/X sky130_fd_sc_hd__and3_2
Xhold447 _3941_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold458 hold458/A VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold469 hold469/A VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6213_ _7017_/Q _6177_/X _6210_/X _6212_/X VGND VGND VPWR VPWR _6214_/D sky130_fd_sc_hd__a211o_1
X_3425_ _6811_/Q _5341_/A _5494_/C _3424_/X _6951_/Q VGND VGND VPWR VPWR _3437_/B
+ sky130_fd_sc_hd__a32o_1
X_7193_ _7237_/CLK _7193_/D fanout578/X VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ hold37/X hold42/X _5324_/B VGND VGND VPWR VPWR _3356_/X sky130_fd_sc_hd__and3b_1
X_6144_ _7187_/Q _6177_/A _6425_/B _7188_/Q VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__and4b_4
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _7120_/Q VGND VGND VPWR VPWR _5632_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _3994_/X VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6767_/Q wire398/X _6028_/C _7274_/Q _5780_/X VGND VGND VPWR VPWR _6075_/X
+ sky130_fd_sc_hd__a32o_1
X_3287_ _4698_/A VGND VGND VPWR VPWR _4662_/B sky130_fd_sc_hd__inv_6
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _5387_/X VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 _5450_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1147 _5280_/X VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 _3955_/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5026_ _4581_/B _4589_/C _5012_/X _4922_/C VGND VGND VPWR VPWR _5177_/B sky130_fd_sc_hd__a31o_1
XFILLER_85_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1169 _6592_/Q VGND VGND VPWR VPWR _3914_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_309 _6118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7031_/CLK _6977_/D fanout599/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5928_ _6972_/Q _5771_/X _5914_/X _5927_/X VGND VGND VPWR VPWR _5928_/X sky130_fd_sc_hd__a211o_2
XFILLER_139_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5859_ _5851_/X _6072_/B _5856_/X _5854_/X _5858_/X VGND VGND VPWR VPWR _5859_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_119_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold970 _5287_/X VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 _4093_/X VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold992 _7299_/A VGND VGND VPWR VPWR hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4190_ hold892/X _6549_/A0 _4204_/S VGND VGND VPWR VPWR _4190_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6900_ _7133_/CLK _6900_/D fanout601/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_2
X_6831_ _6855_/CLK _6831_/D fanout583/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6762_ _6768_/CLK _6762_/D fanout576/X VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_4
X_3974_ hold144/X hold5/X _3974_/S VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__mux2_1
X_5713_ _5759_/B _5712_/Y _7180_/Q VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__mux2_1
X_6693_ _7148_/CLK _6693_/D fanout591/X VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5644_ hold5/X _5644_/A1 hold9/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__mux2_1
XFILLER_148_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5575_ hold17/X hold66/A _5575_/C _5575_/D VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__and4_4
Xhold200 _6590_/Q VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__dlygate4sd3_1
X_7314_ _7314_/A VGND VGND VPWR VPWR _7314_/X sky130_fd_sc_hd__buf_2
Xhold211 hold211/A VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4526_ _5090_/A _5090_/B _4586_/B VGND VGND VPWR VPWR _4589_/B sky130_fd_sc_hd__and3_1
Xhold222 _7033_/Q VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _5453_/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _7019_/Q VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold255 _5490_/X VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7245_ _7245_/CLK _7245_/D fanout597/X VGND VGND VPWR VPWR _7245_/Q sky130_fd_sc_hd__dfrtp_2
Xhold266 _7083_/Q VGND VGND VPWR VPWR hold266/X sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _5055_/D _5143_/A _5260_/B VGND VGND VPWR VPWR _4457_/X sky130_fd_sc_hd__and3_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold277 hold277/A VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold288 _6937_/Q VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold299 _6904_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ _6524_/A _4127_/C _5273_/D VGND VGND VPWR VPWR _4133_/B sky130_fd_sc_hd__and3_4
X_7176_ _7218_/CLK _7176_/D fanout577/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4388_ _4729_/A _4860_/C VGND VGND VPWR VPWR _4388_/Y sky130_fd_sc_hd__nand2_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6127_ _6444_/B _6444_/C _6113_/X _6125_/X _6323_/B1 VGND VGND VPWR VPWR _6127_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _6791_/Q user_clock _6853_/Q VGND VGND VPWR VPWR _3339_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6058_ _6646_/Q _5783_/X _5789_/X _6781_/Q _6057_/X VGND VGND VPWR VPWR _6058_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _5008_/X _5009_/B _5009_/C VGND VGND VPWR VPWR _5009_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_38_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _6134_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 _6246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _6750_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _6635_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3690_ _6953_/Q _3424_/X _3438_/X _7001_/Q _3689_/X VGND VGND VPWR VPWR _3690_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5360_ _5667_/A0 hold972/X _5367_/S VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__mux2_1
Xoutput305 _3345_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput316 hold498/X VGND VGND VPWR VPWR hold499/A sky130_fd_sc_hd__buf_12
XFILLER_160_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput327 hold595/X VGND VGND VPWR VPWR hold596/A sky130_fd_sc_hd__buf_12
Xoutput338 hold694/X VGND VGND VPWR VPWR hold695/A sky130_fd_sc_hd__buf_12
X_4311_ _4318_/A _4318_/B VGND VGND VPWR VPWR _5090_/A sky130_fd_sc_hd__nand2_4
X_5291_ hold950/X _6539_/A0 _5294_/S VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7030_ _7117_/CLK _7030_/D fanout608/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_2
X_4242_ _4734_/B _4416_/B VGND VGND VPWR VPWR _4284_/A sky130_fd_sc_hd__nand2b_4
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4173_ hold653/X _5667_/A0 _4187_/S VGND VGND VPWR VPWR _4173_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6814_ _7263_/CLK _6814_/D fanout578/X VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfrtp_2
X_6745_ _7271_/CLK _6745_/D fanout597/X VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfstp_2
X_3957_ _6539_/A0 _3957_/A1 _3959_/S VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6676_ _6676_/CLK _6676_/D fanout578/X VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfstp_2
X_3888_ _7030_/Q _3515_/X _3884_/X _3885_/X _3887_/X VGND VGND VPWR VPWR _3889_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5627_ hold21/X _5627_/A1 _5628_/S VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__mux2_1
XFILLER_191_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5558_ _5649_/A0 _5558_/A1 _5565_/S VGND VGND VPWR VPWR _5558_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4509_ _4509_/A _4509_/B _4509_/C _4509_/D VGND VGND VPWR VPWR _4620_/B sky130_fd_sc_hd__and4_4
XFILLER_104_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5489_ hold660/X _3921_/B _5493_/S VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7228_ _7254_/CLK _7228_/D VGND VGND VPWR VPWR _7228_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout510 hold21/X VGND VGND VPWR VPWR _4051_/B sky130_fd_sc_hd__buf_6
XFILLER_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout521 hold50/X VGND VGND VPWR VPWR _3922_/C sky130_fd_sc_hd__buf_6
Xfanout532 hold98/X VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__buf_8
XFILLER_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout543 hold65/X VGND VGND VPWR VPWR _5324_/B sky130_fd_sc_hd__buf_6
XFILLER_76_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7159_ _7159_/CLK _7159_/D fanout599/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfstp_1
Xfanout565 _4716_/A VGND VGND VPWR VPWR _4939_/A sky130_fd_sc_hd__buf_8
Xfanout576 fanout581/X VGND VGND VPWR VPWR fanout576/X sky130_fd_sc_hd__buf_8
XFILLER_19_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout587 fanout588/X VGND VGND VPWR VPWR fanout587/X sky130_fd_sc_hd__buf_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout598 input75/X VGND VGND VPWR VPWR fanout598/X sky130_fd_sc_hd__buf_6
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4860_ _4987_/B _4860_/B _4860_/C VGND VGND VPWR VPWR _4860_/X sky130_fd_sc_hd__and3_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ _3811_/A _3811_/B _3811_/C VGND VGND VPWR VPWR _3811_/Y sky130_fd_sc_hd__nand3_2
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4791_ _4945_/B _4791_/B _4945_/C VGND VGND VPWR VPWR _4791_/X sky130_fd_sc_hd__and3_1
XANTENNA_17 _3424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _5611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_39 _3496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6542_/A _6536_/C _6530_/C _6530_/D VGND VGND VPWR VPWR _6535_/S sky130_fd_sc_hd__nand4_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3742_ input46/X _3368_/X _5684_/B _3539_/X input55/X VGND VGND VPWR VPWR _3742_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6461_ _6568_/Q _6118_/X _6137_/X _7274_/Q _6460_/X VGND VGND VPWR VPWR _6461_/X
+ sky130_fd_sc_hd__a221o_1
X_3673_ _7241_/Q _6536_/A _5325_/C _5566_/B _7065_/Q VGND VGND VPWR VPWR _3673_/X
+ sky130_fd_sc_hd__a32o_1
X_5412_ _4053_/B hold188/X _5412_/S VGND VGND VPWR VPWR _5412_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6392_ _6391_/Y _6390_/X _6392_/B1 _6442_/S VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_161_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5343_ hold346/X _3916_/C _5349_/S VGND VGND VPWR VPWR _5343_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput179 _3272_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
X_5274_ _3370_/B _5274_/A1 _5278_/S VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7013_ _7119_/CLK _7013_/D fanout592/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4225_ _4307_/A _4307_/B _4225_/C VGND VGND VPWR VPWR _4416_/A sky130_fd_sc_hd__nand3_2
X_4156_ _6546_/A0 hold517/X _4156_/S VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4087_ _4087_/A0 _4086_/X _4093_/S VGND VGND VPWR VPWR _4087_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4989_ _4859_/C _4862_/A _4859_/D _4673_/X _4988_/X VGND VGND VPWR VPWR _4989_/X
+ sky130_fd_sc_hd__a311o_1
X_6728_ _7239_/CLK _6728_/D fanout576/X VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6659_ _6843_/CLK _6659_/D fanout584/X VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4010_ hold952/X _6535_/A0 _4010_/S VGND VGND VPWR VPWR _4010_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5961_ _6982_/Q _6073_/B2 _5774_/X _6910_/Q _5960_/X VGND VGND VPWR VPWR _5961_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4912_ _4903_/A _5173_/C _4562_/C VGND VGND VPWR VPWR _5174_/D sky130_fd_sc_hd__a21oi_1
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5892_ _6883_/Q _5768_/X _5794_/X _6923_/Q _5890_/X VGND VGND VPWR VPWR _5892_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4843_ _4843_/A _4843_/B _4843_/C _4843_/D VGND VGND VPWR VPWR _4843_/Y sky130_fd_sc_hd__nor4_1
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4774_ _5263_/C _4774_/B VGND VGND VPWR VPWR _4776_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6513_ _7238_/Q _7255_/Q _6486_/C VGND VGND VPWR VPWR _6513_/X sky130_fd_sc_hd__o21a_1
X_3725_ _7263_/Q _5512_/B _3457_/X _3724_/X VGND VGND VPWR VPWR _3725_/X sky130_fd_sc_hd__a31o_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6444_ _6596_/Q _6444_/B _6444_/C VGND VGND VPWR VPWR _6444_/X sky130_fd_sc_hd__and3_1
XFILLER_119_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3656_ _6571_/Q _6548_/A _5341_/A _3463_/X _7113_/Q VGND VGND VPWR VPWR _3656_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_106_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6375_ _6674_/Q _6129_/A _6101_/X _6684_/Q _6374_/X VGND VGND VPWR VPWR _6380_/B
+ sky130_fd_sc_hd__a221o_1
X_3587_ input12/X _3528_/X _3584_/X _3585_/X _3586_/X VGND VGND VPWR VPWR _3587_/X
+ sky130_fd_sc_hd__a2111o_2
X_5326_ _5326_/A0 _5649_/A0 _5326_/S VGND VGND VPWR VPWR _5326_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5257_ _5257_/A _5257_/B _5257_/C _5257_/D VGND VGND VPWR VPWR _5258_/D sky130_fd_sc_hd__and4_1
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4208_ _4632_/C _4612_/C VGND VGND VPWR VPWR _4208_/Y sky130_fd_sc_hd__nand2_8
XFILLER_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5188_ _4293_/Y _4514_/Y _5187_/X VGND VGND VPWR VPWR _5188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4139_ _6542_/A _5273_/D _4139_/C VGND VGND VPWR VPWR _4144_/S sky130_fd_sc_hd__and3_2
XFILLER_113_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3510_ _6548_/A _6548_/D _5675_/D VGND VGND VPWR VPWR _3510_/X sky130_fd_sc_hd__and3_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4490_ _4801_/A _4789_/B VGND VGND VPWR VPWR _4490_/Y sky130_fd_sc_hd__nand2_4
Xhold607 _7077_/Q VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 hold618/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
Xhold629 hold629/A VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _5304_/A _5311_/C _5630_/C VGND VGND VPWR VPWR _3441_/X sky130_fd_sc_hd__and3_2
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6160_ _7119_/Q _5750_/X _6115_/X _7135_/Q _6159_/X VGND VGND VPWR VPWR _6165_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3372_ _6542_/A _3372_/B VGND VGND VPWR VPWR _3377_/S sky130_fd_sc_hd__nand2_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5111_ _4939_/A _4738_/B _5128_/B _4982_/D _4862_/A VGND VGND VPWR VPWR _5111_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6091_/A1 _5761_/X _6090_/X _6089_/X VGND VGND VPWR VPWR _7206_/D sky130_fd_sc_hd__o22a_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1307 _7229_/Q VGND VGND VPWR VPWR hold211/A sky130_fd_sc_hd__dlygate4sd3_1
X_5042_ _5042_/A _5042_/B _5143_/C VGND VGND VPWR VPWR _5260_/C sky130_fd_sc_hd__and3_1
Xhold1318 _7121_/Q VGND VGND VPWR VPWR _5633_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 _5285_/X VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6993_ _7159_/CLK _6993_/D fanout599/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7145_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5944_ _7069_/Q _5826_/B _6010_/C _6010_/D _5943_/X VGND VGND VPWR VPWR _5944_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_53_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5875_ _6970_/Q _5771_/X _5795_/X _6898_/Q VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4826_ _4505_/B _5044_/A _4597_/C _4418_/X VGND VGND VPWR VPWR _4827_/C sky130_fd_sc_hd__a31oi_2
Xclkbuf_leaf_66_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7015_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _4786_/B _4939_/B _4756_/C _4755_/B _4774_/B VGND VGND VPWR VPWR _4757_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3708_ _6766_/Q _5485_/B _4139_/C _3452_/X _6962_/Q VGND VGND VPWR VPWR _3708_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4688_ _4688_/A _4688_/B _4688_/C VGND VGND VPWR VPWR _4688_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6427_ _6746_/Q _6446_/B _6347_/C _6097_/X _6761_/Q VGND VGND VPWR VPWR _6427_/X
+ sky130_fd_sc_hd__a32o_1
X_3639_ _3350_/B hold56/A _3446_/X _4092_/S input58/X VGND VGND VPWR VPWR _3639_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_122_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6358_ _6673_/Q _6129_/A _6098_/X _6748_/Q _6357_/X VGND VGND VPWR VPWR _6365_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5309_ _5309_/A0 hold2/X hold40/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__mux2_1
X_6289_ _7140_/Q _6115_/X _6119_/X _7052_/Q _6288_/X VGND VGND VPWR VPWR _6290_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6875_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3990_ _3918_/B hold532/X _3992_/S VGND VGND VPWR VPWR _3990_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5660_ hold8/X _3474_/X _3918_/X _5665_/S hold828/X VGND VGND VPWR VPWR _5660_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4611_ _4611_/A _4611_/B _4611_/C VGND VGND VPWR VPWR _4617_/A sky130_fd_sc_hd__nand3_1
XFILLER_176_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5591_ _4051_/B hold841/X hold44/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4542_ _4698_/A _4657_/C VGND VGND VPWR VPWR _4674_/D sky130_fd_sc_hd__and2b_4
XFILLER_190_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold404 hold404/A VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold415 _6900_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlygate4sd3_1
X_7261_ _7278_/CLK _7261_/D fanout597/X VGND VGND VPWR VPWR _7261_/Q sky130_fd_sc_hd__dfrtp_4
Xhold426 _7014_/Q VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4632_/B _4489_/C VGND VGND VPWR VPWR _4473_/Y sky130_fd_sc_hd__nand2_2
Xhold437 _6821_/Q VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _6747_/Q VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _6634_/Q VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _7105_/Q _6112_/X _6145_/X _7009_/Q _6211_/X VGND VGND VPWR VPWR _6212_/X
+ sky130_fd_sc_hd__a221o_1
X_3424_ _5476_/C _5494_/C _5575_/C VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__and3_4
XFILLER_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7192_ _7237_/CLK _7192_/D fanout578/X VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6143_ _6141_/B _6444_/C _6143_/C _6143_/D VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__and4b_4
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3355_ hold71/X hold26/X hold65/A VGND VGND VPWR VPWR _3355_/X sky130_fd_sc_hd__and3b_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6662_/Q _5794_/X _6072_/X _6073_/X _6071_/X VGND VGND VPWR VPWR _6074_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold1104 _5632_/X VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 hold1383/X VGND VGND VPWR VPWR _5296_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _4729_/A VGND VGND VPWR VPWR _4860_/B sky130_fd_sc_hd__inv_8
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _6564_/Q VGND VGND VPWR VPWR _3380_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1137 hold1385/X VGND VGND VPWR VPWR _5540_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5025_ _4575_/B _4589_/C _5012_/X _4918_/X VGND VGND VPWR VPWR _5027_/B sky130_fd_sc_hd__a31o_1
Xhold1148 hold1433/X VGND VGND VPWR VPWR _5576_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1159 _6763_/Q VGND VGND VPWR VPWR _4140_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6976_ _6976_/CLK _6976_/D fanout590/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_159_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5927_ _6948_/Q _5779_/X _5782_/X _6940_/Q _5926_/X VGND VGND VPWR VPWR _5927_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5858_ _6905_/Q _5774_/X _5794_/X _6921_/Q _5857_/X VGND VGND VPWR VPWR _5858_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _4507_/Y _4621_/Y _4808_/Y _4206_/Y VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__a31oi_1
X_5789_ _7181_/Q _7180_/Q _5814_/C _5795_/D VGND VGND VPWR VPWR _5789_/X sky130_fd_sc_hd__and4_4
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold960 _7174_/Q VGND VGND VPWR VPWR hold960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 hold971/A VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold982 _6765_/Q VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _4067_/X VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6830_ _6855_/CLK _6830_/D fanout583/X VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6761_ _6761_/CLK _6761_/D fanout572/X VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3973_ hold475/X _3921_/B _3974_/S VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__mux2_1
X_5712_ _6800_/Q _5759_/B VGND VGND VPWR VPWR _5712_/Y sky130_fd_sc_hd__nor2_4
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6692_ _7264_/CLK _6692_/D fanout579/X VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5643_ hold24/X hold52/X hold9/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__mux2_1
XFILLER_148_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5574_ _5692_/A1 hold909/X _5574_/S VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__mux2_1
X_7313_ _7313_/A VGND VGND VPWR VPWR _7313_/X sky130_fd_sc_hd__clkbuf_2
Xhold201 _3911_/X VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _5090_/A _5090_/B _4606_/B _4606_/D VGND VGND VPWR VPWR _4525_/Y sky130_fd_sc_hd__nand4_2
Xhold212 _5323_/X VGND VGND VPWR VPWR _5324_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _5533_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _6874_/Q VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _5517_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7244_ _7244_/CLK _7244_/D fanout580/X VGND VGND VPWR VPWR _7244_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold256 _7140_/Q VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4456_/A _4456_/B _4456_/C VGND VGND VPWR VPWR _4456_/Y sky130_fd_sc_hd__nand3_1
Xhold267 _5589_/X VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold278 _7011_/Q VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _5425_/X VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ hold75/X hold16/X hold54/X _5324_/B VGND VGND VPWR VPWR _3407_/X sky130_fd_sc_hd__and4b_4
X_7175_ _7219_/CLK _7175_/D fanout577/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4387_ _4632_/A _4511_/A _4789_/B VGND VGND VPWR VPWR _5255_/B sky130_fd_sc_hd__and3_2
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6126_ _7187_/Q _6136_/A _6143_/C _7188_/Q VGND VGND VPWR VPWR _6126_/X sky130_fd_sc_hd__and4b_4
X_3338_ input1/X _6874_/Q _3337_/Y VGND VGND VPWR VPWR _3338_/Y sky130_fd_sc_hd__o21ai_4
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6057_ _7273_/Q _5780_/X _5794_/X _6661_/Q VGND VGND VPWR VPWR _6057_/X sky130_fd_sc_hd__a22o_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3269_ _7002_/Q VGND VGND VPWR VPWR _3269_/Y sky130_fd_sc_hd__inv_2
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ _5128_/A _5128_/B _4732_/C _4970_/B _4689_/C VGND VGND VPWR VPWR _5008_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_107 _6136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_118 _6246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _6984_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ _7135_/CLK _6959_/D fanout588/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_179_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold790 _3983_/X VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1490 _6617_/Q VGND VGND VPWR VPWR _3951_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput306 _3343_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
Xoutput317 hold643/X VGND VGND VPWR VPWR hold644/A sky130_fd_sc_hd__buf_12
Xoutput328 hold548/X VGND VGND VPWR VPWR hold549/A sky130_fd_sc_hd__buf_12
X_4310_ _4747_/A _4310_/B _4310_/C _4310_/D VGND VGND VPWR VPWR _4318_/B sky130_fd_sc_hd__nand4_2
X_5290_ hold372/X _6538_/A0 _5294_/S VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__mux2_1
Xoutput339 hold577/X VGND VGND VPWR VPWR hold578/A sky130_fd_sc_hd__buf_12
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4241_ _4734_/B _4416_/B VGND VGND VPWR VPWR _4346_/A sky130_fd_sc_hd__and2b_2
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ _4187_/S _3539_/X _4171_/Y _4076_/X VGND VGND VPWR VPWR _4188_/S sky130_fd_sc_hd__o211a_4
XFILLER_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6813_ _7267_/CLK _6813_/D fanout572/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3956_ _6538_/A0 hold461/X _3959_/S VGND VGND VPWR VPWR _3956_/X sky130_fd_sc_hd__mux2_1
X_6744_ _7263_/CLK _6744_/D fanout578/X VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6675_ _7265_/CLK _6675_/D fanout575/X VGND VGND VPWR VPWR _6675_/Q sky130_fd_sc_hd__dfrtp_2
X_3887_ _7166_/Q _3509_/X _3559_/X _6910_/Q _3886_/X VGND VGND VPWR VPWR _3887_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5626_ _6505_/A1 hold833/X _5628_/S VGND VGND VPWR VPWR _5626_/X sky130_fd_sc_hd__mux2_1
X_5557_ _6548_/B _5557_/B VGND VGND VPWR VPWR _5565_/S sky130_fd_sc_hd__nand2_8
XFILLER_3_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4508_ _4523_/C _4523_/A _4336_/X VGND VGND VPWR VPWR _4586_/B sky130_fd_sc_hd__a21oi_2
X_5488_ _5488_/A0 _3918_/X _5493_/S VGND VGND VPWR VPWR _5488_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7227_ _7259_/CLK _7227_/D VGND VGND VPWR VPWR _7227_/Q sky130_fd_sc_hd__dfxtp_1
X_4439_ _5042_/A _5060_/C _5042_/B _4439_/D VGND VGND VPWR VPWR _4440_/D sky130_fd_sc_hd__nand4_1
Xfanout500 _5959_/C VGND VGND VPWR VPWR _5934_/C sky130_fd_sc_hd__buf_8
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout511 hold32/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__buf_12
Xfanout522 hold24/X VGND VGND VPWR VPWR _3921_/B sky130_fd_sc_hd__buf_6
Xfanout533 _7188_/Q VGND VGND VPWR VPWR _6143_/D sky130_fd_sc_hd__buf_8
XFILLER_76_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7158_ _7173_/CLK _7158_/D fanout603/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout544 hold64/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__buf_12
XFILLER_59_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout577 fanout579/X VGND VGND VPWR VPWR fanout577/X sky130_fd_sc_hd__buf_8
X_6109_ _6138_/A _6444_/C _6425_/B VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__and3_4
Xfanout588 fanout589/X VGND VGND VPWR VPWR fanout588/X sky130_fd_sc_hd__buf_8
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7089_/CLK _7089_/D fanout596/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout599 input75/X VGND VGND VPWR VPWR fanout599/X sky130_fd_sc_hd__buf_8
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _3810_/A _3810_/B _3810_/C _3810_/D VGND VGND VPWR VPWR _3811_/C sky130_fd_sc_hd__nor4_2
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ _4788_/X _4790_/B _4790_/C VGND VGND VPWR VPWR _4790_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_18 _3757_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _5611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _6595_/Q _5684_/B _3466_/X _3738_/X _3740_/X VGND VGND VPWR VPWR _3751_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_158_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6460_ _6601_/Q _6109_/X _6110_/X _6558_/Q _6459_/X VGND VGND VPWR VPWR _6460_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3672_ _6745_/Q _3368_/X _5485_/B _3548_/X _7049_/Q VGND VGND VPWR VPWR _3672_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5411_ _5404_/B _4073_/X _5412_/S hold839/X VGND VGND VPWR VPWR _5411_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6391_ _6689_/Q _6466_/A1 _5759_/A VGND VGND VPWR VPWR _6391_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5342_ _5342_/A0 _5649_/A0 _5349_/S VGND VGND VPWR VPWR _5342_/X sky130_fd_sc_hd__mux2_1
X_5273_ _6524_/A _6524_/B _6530_/D _5273_/D VGND VGND VPWR VPWR _5278_/S sky130_fd_sc_hd__nand4_4
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7012_ _7156_/CLK _7012_/D fanout602/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_4
X_4224_ _4255_/A _4600_/B _4612_/C _4647_/C VGND VGND VPWR VPWR _4427_/D sky130_fd_sc_hd__nand4_4
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4155_ _4152_/C _3919_/X _4156_/S hold858/X VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4086_ hold69/X _3924_/X _4092_/S VGND VGND VPWR VPWR _4086_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _4716_/A _5128_/B _4945_/B _5255_/A VGND VGND VPWR VPWR _4988_/X sky130_fd_sc_hd__o211a_1
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6727_ _6855_/CLK _6727_/D fanout583/X VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfstp_2
X_3939_ _6524_/A _6536_/B _6530_/C _4127_/C VGND VGND VPWR VPWR _3944_/S sky130_fd_sc_hd__nand4_4
XFILLER_177_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6658_ _6827_/CLK _6658_/D fanout573/X VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5609_ hold21/X hold132/X _5610_/S VGND VGND VPWR VPWR _5609_/X sky130_fd_sc_hd__mux2_1
X_6589_ _6761_/CLK _6589_/D fanout572/X VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5960_ _7038_/Q _5826_/B _5773_/X _5959_/X VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__a31o_1
XFILLER_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4911_ _4601_/Y _5248_/A3 _4648_/Y _4560_/B _4909_/X VGND VGND VPWR VPWR _4914_/B
+ sky130_fd_sc_hd__o311a_1
X_5891_ _5934_/C _6072_/C _6891_/Q _5776_/X _6955_/Q VGND VGND VPWR VPWR _5891_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_45_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_290 _5814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4842_ _5060_/A _5060_/B _5055_/D _5128_/B VGND VGND VPWR VPWR _4843_/C sky130_fd_sc_hd__and4_1
XFILLER_178_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4773_ _4773_/A _4773_/B _4773_/C VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__nor3_1
XFILLER_21_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6512_ _7249_/Q _7253_/D _6512_/A3 _4206_/B wire406/X VGND VGND VPWR VPWR _7237_/D
+ sky130_fd_sc_hd__o41ai_2
X_3724_ _7066_/Q _5512_/B hold39/A _3488_/X _7074_/Q VGND VGND VPWR VPWR _3724_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6443_ _6442_/X _6467_/A2 _6443_/S VGND VGND VPWR VPWR _7218_/D sky130_fd_sc_hd__mux2_1
X_3655_ _7041_/Q _5512_/B _5684_/C _5503_/B _7009_/Q VGND VGND VPWR VPWR _3655_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6374_ _6560_/Q _6446_/B _6446_/C _6138_/X _6608_/Q VGND VGND VPWR VPWR _6374_/X
+ sky130_fd_sc_hd__a32o_1
X_3586_ _7152_/Q _3550_/X _3553_/X _6679_/Q VGND VGND VPWR VPWR _3586_/X sky130_fd_sc_hd__a22o_1
X_5325_ _6524_/B _5666_/C _5325_/C VGND VGND VPWR VPWR _5326_/S sky130_fd_sc_hd__and3_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5256_ _4939_/A _5255_/A _5263_/C _5255_/X _4872_/D VGND VGND VPWR VPWR _5257_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4207_ _4600_/B _4612_/C VGND VGND VPWR VPWR _4970_/D sky130_fd_sc_hd__and2_4
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _5187_/A _5234_/B _5234_/C VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__and3_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4138_ _6535_/A0 _4138_/A1 _4138_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4069_ hold8/X _3539_/X _3918_/X hold57/X hold542/X VGND VGND VPWR VPWR _4069_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold608 _5582_/X VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _6999_/Q hold39/A _3407_/X _3439_/X VGND VGND VPWR VPWR _3440_/X sky130_fd_sc_hd__a31o_1
Xhold619 _7303_/A VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_3371_ _5476_/B _6536_/A _6536_/C VGND VGND VPWR VPWR _3372_/B sky130_fd_sc_hd__and3_2
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5110_ _4754_/B _4255_/A _4789_/B _4939_/A VGND VGND VPWR VPWR _5110_/X sky130_fd_sc_hd__a31o_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _6442_/S _6090_/A2 _6443_/S VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__a21o_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _4557_/B _4860_/B _4751_/A _4860_/C VGND VGND VPWR VPWR _5143_/C sky130_fd_sc_hd__a211o_2
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 _5658_/X VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1319 _7001_/Q VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6992_ _7122_/CLK _6992_/D fanout606/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5943_ _7125_/Q _5826_/B _5911_/C _5940_/X _5942_/X VGND VGND VPWR VPWR _5943_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5874_ _6890_/Q _5815_/B _5815_/C _5826_/B _5873_/X VGND VGND VPWR VPWR _5874_/X
+ sky130_fd_sc_hd__a311o_1
X_4825_ _4271_/Y _4514_/Y _4423_/Y _4348_/X VGND VGND VPWR VPWR _4827_/B sky130_fd_sc_hd__a211o_1
XFILLER_138_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4756_ _4760_/C _4786_/B _4756_/C _4760_/B VGND VGND VPWR VPWR _4756_/Y sky130_fd_sc_hd__nand4_1
X_3707_ _6845_/Q _5323_/S _3700_/X _3703_/X _3706_/X VGND VGND VPWR VPWR _3717_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4687_ _4939_/A _4687_/B VGND VGND VPWR VPWR _4688_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3638_ _6897_/Q _5377_/C _3636_/X _3637_/X VGND VGND VPWR VPWR _3652_/A sky130_fd_sc_hd__a211o_1
X_6426_ _6641_/Q _6177_/X _6425_/X _6424_/X _6423_/X VGND VGND VPWR VPWR _6431_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6357_ _7244_/Q _6465_/A2 _6106_/C _6129_/D _6668_/Q VGND VGND VPWR VPWR _6357_/X
+ sky130_fd_sc_hd__a32o_1
X_3569_ _3568_/Y _3569_/A1 _3906_/S VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5308_ hold312/X _3916_/C hold40/X VGND VGND VPWR VPWR _5308_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6288_ _7020_/Q _6177_/C _6110_/C _6135_/X _6940_/Q VGND VGND VPWR VPWR _6288_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_103_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5239_ _4753_/A _4753_/B _4549_/D _5036_/B VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__a211o_1
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__buf_12
XFILLER_94_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4610_ _4333_/A _4484_/D _5216_/A VGND VGND VPWR VPWR _4611_/C sky130_fd_sc_hd__a21oi_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ _6505_/A1 hold830/X hold44/X VGND VGND VPWR VPWR _5590_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4541_ _4606_/B _4584_/B _4544_/B _4544_/D VGND VGND VPWR VPWR _4541_/Y sky130_fd_sc_hd__nand4_1
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold405 _6819_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
X_7260_ _7260_/CLK _7260_/D fanout572/X VGND VGND VPWR VPWR _7260_/Q sky130_fd_sc_hd__dfrtp_4
Xhold416 _5383_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4472_ _4632_/A _4600_/B _5036_/B VGND VGND VPWR VPWR _4557_/B sky130_fd_sc_hd__nor3_2
Xhold427 _5511_/X VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold438 _5286_/X VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _6743_/Q _3418_/X _3422_/X _3417_/X _3415_/X VGND VGND VPWR VPWR _3437_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold449 _4120_/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6211_ _6993_/Q _6176_/B _6143_/C _6137_/X _7097_/Q VGND VGND VPWR VPWR _6211_/X
+ sky130_fd_sc_hd__a32o_1
X_7191_ _7219_/CLK _7191_/D fanout578/X VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _7187_/Q _6177_/A _6143_/C _6143_/D VGND VGND VPWR VPWR _6142_/X sky130_fd_sc_hd__and4b_4
X_3354_ _7249_/Q _3354_/B VGND VGND VPWR VPWR _7255_/D sky130_fd_sc_hd__and2_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6752_/Q _5842_/C _6028_/C _6757_/Q _6073_/B2 VGND VGND VPWR VPWR _6073_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1105 _7009_/Q VGND VGND VPWR VPWR _5506_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_3285_ _4511_/A VGND VGND VPWR VPWR _5036_/B sky130_fd_sc_hd__inv_6
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _6569_/Q VGND VGND VPWR VPWR _3389_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _3380_/X VGND VGND VPWR VPWR _6564_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5024_ _5264_/C _5024_/B _5174_/C _5265_/B VGND VGND VPWR VPWR _5027_/A sky130_fd_sc_hd__nand4_1
Xhold1138 _6789_/Q VGND VGND VPWR VPWR _4184_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _7275_/Q VGND VGND VPWR VPWR _6549_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _7071_/CLK _6975_/D fanout585/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfstp_2
X_5926_ _7092_/Q _5826_/B wire398/X _5795_/X _6900_/Q VGND VGND VPWR VPWR _5926_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5857_ _7001_/Q _5782_/C _5795_/C _5971_/A2 hold59/A VGND VGND VPWR VPWR _5857_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_179_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4808_ _4808_/A _4808_/B VGND VGND VPWR VPWR _4808_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5788_ _5911_/C _5795_/D VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__and2_4
XFILLER_166_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4739_ _5128_/A _5128_/C _5263_/B _4738_/X VGND VGND VPWR VPWR _4739_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6409_ _6675_/Q _6129_/A _6129_/D _6670_/Q _6408_/X VGND VGND VPWR VPWR _6414_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold950 _6825_/Q VGND VGND VPWR VPWR hold950/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold961 _5692_/X VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 _6879_/Q VGND VGND VPWR VPWR hold972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _4142_/X VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold994 _7079_/Q VGND VGND VPWR VPWR hold994/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7165_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7037_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6760_ _7267_/CLK _6760_/D _3291_/A VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfstp_2
X_3972_ hold224/X hold2/X _3974_/S VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ _5711_/A _5711_/B _5711_/C VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__and3_1
X_6691_ _6761_/CLK _6691_/D fanout572/X VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfstp_1
X_5642_ _3918_/B hold641/X hold9/X VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5573_ _4051_/B hold720/X _5574_/S VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7312_ _7312_/A VGND VGND VPWR VPWR _7312_/X sky130_fd_sc_hd__buf_2
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 _6651_/Q VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _4606_/B _4923_/A _4606_/D VGND VGND VPWR VPWR _4592_/B sky130_fd_sc_hd__and3_1
Xhold213 _5324_/X VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _6635_/Q VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7099_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold235 _5354_/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7243_ _7248_/CLK _7243_/D fanout580/X VGND VGND VPWR VPWR _7243_/Q sky130_fd_sc_hd__dfrtp_1
Xhold246 _7107_/Q VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4455_ _5128_/B _4689_/A VGND VGND VPWR VPWR _4456_/C sky130_fd_sc_hd__nand2_1
Xhold257 _5654_/X VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold268 _6992_/Q VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _5508_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _6530_/D _5666_/C _5476_/C VGND VGND VPWR VPWR _3406_/X sky130_fd_sc_hd__and3_1
XFILLER_132_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7174_ _7174_/CLK _7174_/D fanout602/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
X_4386_ _4600_/B _4612_/C VGND VGND VPWR VPWR _4753_/B sky130_fd_sc_hd__nand2b_2
XFILLER_131_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3337_ input1/X input2/X VGND VGND VPWR VPWR _3337_/Y sky130_fd_sc_hd__nand2_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6125_ _6444_/C _6124_/Y _6143_/C _7188_/Q VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__o211a_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6056_ _6052_/X _6053_/X _6055_/X _6051_/X _6049_/X VGND VGND VPWR VPWR _6056_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3268_ _7010_/Q VGND VGND VPWR VPWR _3268_/Y sky130_fd_sc_hd__inv_2
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5007_ _5007_/A _5007_/B _5007_/C _5225_/B VGND VGND VPWR VPWR _5009_/C sky130_fd_sc_hd__nor4b_1
XFILLER_39_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _6136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_119 _6371_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _7053_/CLK _6958_/D fanout603/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5909_ _5909_/A1 _5761_/X _5908_/X VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__o21a_1
X_6889_ _6889_/CLK _6889_/D fanout584/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 hold780/A VGND VGND VPWR VPWR hold780/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 hold791/A VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1480 _6628_/Q VGND VGND VPWR VPWR _3964_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 _6739_/Q VGND VGND VPWR VPWR hold206/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput307 _3342_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
Xoutput318 hold534/X VGND VGND VPWR VPWR hold535/A sky130_fd_sc_hd__buf_12
Xoutput329 hold601/X VGND VGND VPWR VPWR hold602/A sky130_fd_sc_hd__buf_12
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _4760_/B _4637_/A VGND VGND VPWR VPWR _4416_/B sky130_fd_sc_hd__nand2_2
XFILLER_113_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4171_ _5326_/A0 _3249_/A _3346_/D _4187_/S VGND VGND VPWR VPWR _4171_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6812_ _6812_/CLK _6812_/D fanout580/X VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ _7267_/CLK _6743_/D _3291_/A VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfrtp_2
X_3955_ _3370_/B _3955_/A1 _3959_/S VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__mux2_1
X_6674_ _6843_/CLK _6674_/D fanout576/X VGND VGND VPWR VPWR _6674_/Q sky130_fd_sc_hd__dfrtp_2
X_3886_ _7038_/Q _3547_/X _5593_/B _7094_/Q VGND VGND VPWR VPWR _3886_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5625_ _3924_/B hold708/X _5628_/S VGND VGND VPWR VPWR _5625_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5556_ _5692_/A1 hold901/X _5556_/S VGND VGND VPWR VPWR _5556_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4507_ _4505_/X _4504_/Y _4266_/Y VGND VGND VPWR VPWR _4507_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_132_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5487_ hold268/X _3915_/B _5493_/S VGND VGND VPWR VPWR _5487_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7226_ _7259_/CLK _7226_/D VGND VGND VPWR VPWR _7226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4438_ _5042_/A _5042_/B _5260_/A _4438_/D VGND VGND VPWR VPWR _4440_/C sky130_fd_sc_hd__nand4_1
Xfanout501 _5959_/C VGND VGND VPWR VPWR _5795_/D sky130_fd_sc_hd__buf_12
Xfanout512 _4049_/B VGND VGND VPWR VPWR _6505_/A1 sky130_fd_sc_hd__buf_8
Xfanout523 hold50/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__buf_6
XFILLER_132_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7157_ _7157_/CLK _7157_/D fanout593/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout534 _7187_/Q VGND VGND VPWR VPWR _6141_/B sky130_fd_sc_hd__buf_6
Xfanout545 hold237/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__buf_8
X_4369_ _4632_/A _4255_/A _4632_/C _4612_/C _4647_/C VGND VGND VPWR VPWR _4369_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_86_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6108_ _6143_/D _7190_/Q _7189_/Q _6141_/B VGND VGND VPWR VPWR _6108_/X sky130_fd_sc_hd__and4bb_4
Xfanout567 _4211_/X VGND VGND VPWR VPWR _4751_/A sky130_fd_sc_hd__buf_8
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout578 fanout579/X VGND VGND VPWR VPWR fanout578/X sky130_fd_sc_hd__buf_4
XFILLER_112_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 input75/X VGND VGND VPWR VPWR fanout589/X sky130_fd_sc_hd__buf_6
XFILLER_59_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7088_ _7088_/CLK _7088_/D fanout590/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6039_ _6760_/Q _5771_/X _6027_/X _6038_/X VGND VGND VPWR VPWR _6039_/X sky130_fd_sc_hd__a211o_1
XFILLER_100_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_19 _3427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3740_ _6577_/Q _3987_/A _6548_/D _5684_/B _3739_/X VGND VGND VPWR VPWR _3740_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3671_ _6831_/Q _5325_/C _5311_/C _7121_/Q _3525_/X VGND VGND VPWR VPWR _3671_/X
+ sky130_fd_sc_hd__a32o_1
X_5410_ hold83/X hold168/X _5412_/S VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6390_ _6369_/X _6371_/X _6390_/C _6390_/D VGND VGND VPWR VPWR _6390_/X sky130_fd_sc_hd__and4bb_1
XFILLER_127_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5341_ _5341_/A hold56/X _5341_/C VGND VGND VPWR VPWR _5349_/S sky130_fd_sc_hd__and3_4
XFILLER_127_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ _5272_/A1 wire442/X _5271_/Y _5268_/Y VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__a211o_1
XFILLER_141_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7011_ _7131_/CLK _7011_/D fanout606/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4223_ _4255_/A _4494_/C _4557_/A _4647_/C VGND VGND VPWR VPWR _4225_/C sky130_fd_sc_hd__and4_1
X_4154_ _3916_/C hold326/X _4156_/S VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ _4085_/A0 _4084_/X _4093_/S VGND VGND VPWR VPWR _4085_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4987_ _4987_/A _4987_/B _4987_/C VGND VGND VPWR VPWR _4987_/X sky130_fd_sc_hd__and3_1
XFILLER_149_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6726_ _6855_/CLK _6726_/D fanout583/X VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfstp_2
X_3938_ _3934_/S hold822/X _3432_/X _3925_/X VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6657_ _6855_/CLK _6657_/D fanout584/X VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfrtp_4
X_3869_ input50/X _3368_/X _5684_/B _5350_/B _6877_/Q VGND VGND VPWR VPWR _3869_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5608_ _6505_/A1 hold816/X _5610_/S VGND VGND VPWR VPWR _5608_/X sky130_fd_sc_hd__mux2_1
X_6588_ _7279_/CLK _6588_/D fanout597/X VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfrtp_4
X_5539_ _5620_/A _6548_/B _5548_/C hold28/X VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__nand4_4
XFILLER_132_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7209_ _7251_/CLK _7209_/D fanout595/X VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout375 _6343_/S VGND VGND VPWR VPWR _6443_/S sky130_fd_sc_hd__buf_8
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _3353_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_155_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4910_ _5263_/A _4746_/A _4755_/B _4581_/B _4557_/X VGND VGND VPWR VPWR _4910_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5890_ _7035_/Q _6072_/B _6003_/C _5889_/X VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__a31o_1
X_4841_ _4841_/A _4841_/B _5165_/C VGND VGND VPWR VPWR _4843_/D sky130_fd_sc_hd__nand3_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 _5511_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_291 _5774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4772_ _5263_/B _5263_/C _4939_/B VGND VGND VPWR VPWR _4773_/B sky130_fd_sc_hd__and3_1
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6511_ _6510_/X _6511_/A1 _6511_/S VGND VGND VPWR VPWR _7236_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3723_ _6562_/Q _6536_/A _5311_/B _3722_/X VGND VGND VPWR VPWR _3723_/X sky130_fd_sc_hd__a31o_1
XFILLER_159_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6442_ _6441_/X _6442_/A1 _6442_/S VGND VGND VPWR VPWR _6442_/X sky130_fd_sc_hd__mux2_1
X_3654_ _7277_/Q _6536_/A _3466_/X _3653_/X VGND VGND VPWR VPWR _3654_/X sky130_fd_sc_hd__a31o_1
XFILLER_161_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6373_ _7276_/Q _6112_/X _6129_/D _6669_/Q _6372_/X VGND VGND VPWR VPWR _6380_/A
+ sky130_fd_sc_hd__a221o_1
X_3585_ input35/X _3469_/X _3471_/X input21/X VGND VGND VPWR VPWR _3585_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5324_ hold12/X _5324_/B _5324_/C VGND VGND VPWR VPWR _5324_/X sky130_fd_sc_hd__and3_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5255_ _5255_/A _5255_/B _5255_/C VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__and3_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4206_ _4206_/A _4206_/B VGND VGND VPWR VPWR _4206_/Y sky130_fd_sc_hd__nor2_1
X_5186_ _5040_/C _4265_/Y _4348_/X _5061_/C _5146_/B VGND VGND VPWR VPWR _5234_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4137_ _6546_/A0 hold555/X _4138_/S VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4068_ hold8/X _3539_/X _3915_/X hold57/X hold496/X VGND VGND VPWR VPWR _4068_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6709_ _7122_/CLK _6709_/D fanout606/X VGND VGND VPWR VPWR _7299_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_138_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold609 _6576_/Q VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3370_ _6536_/B _3370_/B _5311_/B VGND VGND VPWR VPWR _3370_/X sky130_fd_sc_hd__and3_4
XFILLER_170_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5040_ _5040_/A _5040_/B _5040_/C VGND VGND VPWR VPWR _5040_/X sky130_fd_sc_hd__and3_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1309 _6660_/Q VGND VGND VPWR VPWR hold791/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6991_ _7077_/CLK _6991_/D fanout587/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_92_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5942_ _7053_/Q _5826_/B _5815_/C _5814_/C _5941_/X VGND VGND VPWR VPWR _5942_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ _6986_/Q _7183_/Q _7182_/Q _5815_/C _5872_/X VGND VGND VPWR VPWR _5873_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4824_ _4299_/Y _5040_/A _4403_/X _4398_/X VGND VGND VPWR VPWR _4827_/A sky130_fd_sc_hd__a211o_1
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4755_ _4755_/A _4755_/B _4939_/B _4755_/D VGND VGND VPWR VPWR _4755_/Y sky130_fd_sc_hd__nand4_1
XFILLER_147_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3706_ _6994_/Q _3496_/X _5557_/B _7058_/Q _3705_/X VGND VGND VPWR VPWR _3706_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4686_ _4712_/B _4641_/B _4685_/Y VGND VGND VPWR VPWR _4688_/A sky130_fd_sc_hd__a21oi_1
XFILLER_119_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6425_ _7263_/Q _6425_/B _6425_/C VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and3_1
XFILLER_147_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3637_ _6889_/Q _5440_/C _3533_/C _3513_/X _6670_/Q VGND VGND VPWR VPWR _3637_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6356_ _6356_/A _6356_/B _6356_/C _6356_/D VGND VGND VPWR VPWR _6356_/Y sky130_fd_sc_hd__nor4_1
X_3568_ _3568_/A _3568_/B _3568_/C VGND VGND VPWR VPWR _3568_/Y sky130_fd_sc_hd__nand3_4
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ _5307_/A0 _5649_/A0 hold40/X VGND VGND VPWR VPWR _5307_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6287_ _7060_/Q _6118_/X _6137_/X _7100_/Q _6286_/X VGND VGND VPWR VPWR _6290_/C
+ sky130_fd_sc_hd__a221o_1
X_3499_ _3563_/A _5548_/D _5657_/D VGND VGND VPWR VPWR _3499_/X sky130_fd_sc_hd__and3_4
XFILLER_76_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5238_ _5238_/A _5238_/B _5238_/C _5238_/D VGND VGND VPWR VPWR _5238_/Y sky130_fd_sc_hd__nor4_1
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5169_ hold42/A wire442/X _5168_/Y _5150_/X VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__a211o_1
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4540_ _4284_/A _4308_/Y _4689_/C _4754_/B _4314_/X VGND VGND VPWR VPWR _4540_/Y
+ sky130_fd_sc_hd__o2111ai_1
Xwire370 _5869_/Y VGND VGND VPWR VPWR _5883_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold406 _5284_/X VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire392 wire392/A VGND VGND VPWR VPWR wire392/X sky130_fd_sc_hd__buf_2
X_4471_ _4549_/D _4600_/B VGND VGND VPWR VPWR _4489_/C sky130_fd_sc_hd__nor2_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold417 hold417/A VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold428 _6934_/Q VGND VGND VPWR VPWR hold428/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 hold439/A VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6210_ _7065_/Q _6138_/B _6102_/X _6136_/X _7025_/Q VGND VGND VPWR VPWR _6210_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_144_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3422_ _7055_/Q _3563_/A _3902_/A3 _5566_/B _7063_/Q VGND VGND VPWR VPWR _3422_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7190_ _7259_/CLK _7190_/D fanout594/X VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6143_/D _6141_/B _6444_/C _6143_/C VGND VGND VPWR VPWR _6141_/X sky130_fd_sc_hd__and4_4
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _6856_/Q _3353_/B VGND VGND VPWR VPWR _3353_/X sky130_fd_sc_hd__and2_2
XFILLER_124_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6642_/Q _6072_/B _6072_/C VGND VGND VPWR VPWR _6072_/X sky130_fd_sc_hd__and3_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _4632_/A VGND VGND VPWR VPWR _4689_/B sky130_fd_sc_hd__inv_6
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _5506_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _3389_/X VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1128 hold1313/X VGND VGND VPWR VPWR _5531_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _4601_/Y _5248_/A3 _4643_/Y _5022_/Y _4565_/B VGND VGND VPWR VPWR _5265_/B
+ sky130_fd_sc_hd__o311a_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1139 _4184_/X VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6974_ _7006_/CLK _6974_/D fanout603/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5925_ _7116_/Q _5767_/X _5780_/X _7100_/Q _5924_/X VGND VGND VPWR VPWR _5925_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5856_ _7009_/Q _5783_/X _5795_/X _6897_/Q _5855_/X VGND VGND VPWR VPWR _5856_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4807_ _7255_/Q _7257_/Q _7258_/Q _7259_/Q _4806_/Y VGND VGND VPWR VPWR _4808_/A
+ sky130_fd_sc_hd__o41ai_1
X_5787_ _7181_/Q _7180_/Q _7183_/Q _7182_/Q VGND VGND VPWR VPWR _6025_/C sky130_fd_sc_hd__and4_4
X_4738_ _4738_/A _4738_/B _4859_/D VGND VGND VPWR VPWR _4738_/X sky130_fd_sc_hd__and3_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4669_ _4409_/C _4654_/B _4371_/Y _4870_/C _4848_/A VGND VGND VPWR VPWR _4669_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_107_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6408_ _6650_/Q _6177_/A _6106_/C _6177_/X _6640_/Q VGND VGND VPWR VPWR _6408_/X
+ sky130_fd_sc_hd__a32o_1
Xhold940 hold940/A VGND VGND VPWR VPWR hold940/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _5291_/X VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _6672_/Q VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold973 _5360_/X VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold984 _6883_/Q VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _6339_/A _6339_/B _6339_/C _6339_/D VGND VGND VPWR VPWR _6339_/Y sky130_fd_sc_hd__nor4_1
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold995 _5585_/X VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3971_ hold459/X _3916_/C _3974_/S VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5710_ _7177_/Q _7178_/Q _7179_/Q _5710_/D VGND VGND VPWR VPWR _5711_/C sky130_fd_sc_hd__nand4_1
X_6690_ _7268_/CLK _6690_/D fanout572/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5641_ _3915_/B hold391/X hold9/X VGND VGND VPWR VPWR _5641_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ _6505_/A1 hold835/X _5574_/S VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7311_ _7311_/A VGND VGND VPWR VPWR _7311_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4523_ _4523_/A _4656_/C _4523_/C VGND VGND VPWR VPWR _4606_/D sky130_fd_sc_hd__and3_4
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold203 _3991_/X VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _6942_/Q VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlygate4sd3_1
X_7242_ _7260_/CLK _7242_/D fanout579/X VGND VGND VPWR VPWR _7242_/Q sky130_fd_sc_hd__dfrtp_1
Xhold225 _3972_/X VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _6783_/Q VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4454_ _5255_/A _4691_/B _4848_/B _4878_/C VGND VGND VPWR VPWR _4689_/A sky130_fd_sc_hd__and4_2
Xhold247 _5616_/X VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold258 _6908_/Q VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold269 _5487_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ _5324_/B hold37/X _6807_/Q _5675_/D VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__and4_4
X_7173_ _7173_/CLK _7173_/D fanout603/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4385_ _4632_/C _4860_/B VGND VGND VPWR VPWR _4789_/B sky130_fd_sc_hd__nor2_8
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6124_ _7185_/Q _6141_/B VGND VGND VPWR VPWR _6124_/Y sky130_fd_sc_hd__nor2_1
X_3336_ _6717_/Q input3/X input1/X VGND VGND VPWR VPWR _3336_/X sky130_fd_sc_hd__mux2_4
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6562_/Q _6072_/B _6025_/C _6054_/X VGND VGND VPWR VPWR _6055_/X sky130_fd_sc_hd__a31o_1
XFILLER_85_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _7018_/Q VGND VGND VPWR VPWR _3267_/Y sky130_fd_sc_hd__inv_2
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5006_ _5089_/C _4308_/D _4480_/B _5005_/X VGND VGND VPWR VPWR _5225_/B sky130_fd_sc_hd__a31oi_2
XFILLER_94_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_109 _6136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _6957_/CLK _6957_/D fanout591/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ _6292_/S _7197_/Q _6443_/S _5907_/X VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__a211o_1
XFILLER_179_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6888_ _7152_/CLK _6888_/D fanout585/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5839_ _6442_/S _7194_/Q _6443_/S VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold770 _5597_/X VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _6885_/Q VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _6662_/Q VGND VGND VPWR VPWR hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1470 _6625_/Q VGND VGND VPWR VPWR _3961_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1481 _6631_/Q VGND VGND VPWR VPWR _3967_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 _6581_/Q VGND VGND VPWR VPWR _3694_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput308 _3350_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
Xoutput319 hold538/X VGND VGND VPWR VPWR hold539/A sky130_fd_sc_hd__buf_12
XFILLER_153_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4170_ _7253_/D _4170_/B _4170_/C _4170_/D VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__nand4b_1
XFILLER_83_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6811_ _7241_/CLK _6811_/D fanout576/X VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_91_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6742_ _6945_/CLK _6742_/D fanout583/X VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfstp_1
X_3954_ _6536_/B _3954_/B VGND VGND VPWR VPWR _3959_/S sky130_fd_sc_hd__nand2_4
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6673_ _6827_/CLK _6673_/D fanout574/X VGND VGND VPWR VPWR _6673_/Q sky130_fd_sc_hd__dfrtp_2
X_3885_ _7102_/Q _6548_/A _6548_/D _5675_/D VGND VGND VPWR VPWR _3885_/X sky130_fd_sc_hd__and4_1
XFILLER_176_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5624_ hold24/X _5624_/A1 _5628_/S VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__mux2_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5555_ hold21/X hold117/X _5556_/S VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4506_ _5060_/A _4597_/C VGND VGND VPWR VPWR _4506_/Y sky130_fd_sc_hd__nand2_1
X_5486_ _5486_/A0 _5667_/A0 _5493_/S VGND VGND VPWR VPWR _5486_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7225_ _7237_/CLK _7225_/D VGND VGND VPWR VPWR _7225_/Q sky130_fd_sc_hd__dfxtp_2
X_4437_ _4475_/B _4488_/C VGND VGND VPWR VPWR _4440_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout502 _3246_/Y VGND VGND VPWR VPWR _5759_/A sky130_fd_sc_hd__buf_8
Xfanout513 hold83/X VGND VGND VPWR VPWR _4049_/B sky130_fd_sc_hd__buf_6
Xfanout524 _3919_/C VGND VGND VPWR VPWR _6539_/A0 sky130_fd_sc_hd__buf_6
X_7156_ _7156_/CLK _7156_/D fanout602/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4368_ _4409_/C _4654_/B _4870_/C VGND VGND VPWR VPWR _4740_/C sky130_fd_sc_hd__a21oi_2
Xfanout535 _6072_/B VGND VGND VPWR VPWR _6025_/B sky130_fd_sc_hd__buf_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6107_ _6138_/B _6425_/B _6177_/C VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__and3_4
Xfanout557 _4730_/D VGND VGND VPWR VPWR _4786_/B sky130_fd_sc_hd__buf_6
Xfanout568 _4549_/D VGND VGND VPWR VPWR _4632_/A sky130_fd_sc_hd__buf_12
X_3319_ _4214_/A _3319_/B _3319_/C _3319_/D VGND VGND VPWR VPWR _3354_/B sky130_fd_sc_hd__and4b_1
X_7087_ _7087_/CLK _7087_/D fanout589/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfstp_1
Xfanout579 fanout580/X VGND VGND VPWR VPWR fanout579/X sky130_fd_sc_hd__buf_8
X_4299_ _4801_/A _5036_/C VGND VGND VPWR VPWR _4299_/Y sky130_fd_sc_hd__nand2_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6775_/Q _5779_/X _5782_/X _6655_/Q _6037_/X VGND VGND VPWR VPWR _6038_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _6957_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6945_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7129_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3670_ _6993_/Q _3496_/X _3661_/X _3662_/X _3669_/X VGND VGND VPWR VPWR _3692_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5340_ _6505_/A1 _5340_/A1 _5340_/S VGND VGND VPWR VPWR _5340_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5271_ _5210_/A _5252_/Y _5270_/X _5247_/Y VGND VGND VPWR VPWR _5271_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_99_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7010_ _7132_/CLK _7010_/D fanout610/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_4
X_4222_ _4222_/A _4222_/B VGND VGND VPWR VPWR _4307_/B sky130_fd_sc_hd__nor2_2
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4153_ _4153_/A1 _4156_/S _4152_/X VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4084_ hold121/X _3921_/X _4092_/S VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4986_ _5040_/B _4376_/Y _4849_/Y _4659_/Y _4985_/Y VGND VGND VPWR VPWR _5231_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_23_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6725_ _6945_/CLK _6725_/D fanout583/X VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfstp_1
X_3937_ _3934_/S hold860/X _3432_/X _3922_/X VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6656_ _6828_/CLK _6656_/D fanout573/X VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfrtp_4
X_3868_ _7141_/Q _3503_/X _3528_/X input18/X _3867_/X VGND VGND VPWR VPWR _3873_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5607_ _3924_/B hold714/X _5610_/S VGND VGND VPWR VPWR _5607_/X sky130_fd_sc_hd__mux2_1
X_6587_ _7274_/CLK _6587_/D fanout577/X VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfrtp_4
X_3799_ _3799_/A1 _4092_/S _3521_/X _7171_/Q _3798_/X VGND VGND VPWR VPWR _3799_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_152_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5538_ _5538_/A0 _5692_/A1 _5538_/S VGND VGND VPWR VPWR _5538_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5469_ hold89/X hold148/X _5475_/S VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7208_ _7256_/CLK _7208_/D fanout595/X VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7139_ _7145_/CLK _7139_/D fanout602/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout376 _5263_/A VGND VGND VPWR VPWR _4923_/A sky130_fd_sc_hd__buf_4
XFILLER_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4840_ _4356_/A _4848_/A _4259_/Y _4295_/A _4506_/Y VGND VGND VPWR VPWR _4841_/B
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_270 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 _5711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_292 _6009_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4771_ _4923_/B _5263_/C _4939_/B VGND VGND VPWR VPWR _4773_/A sky130_fd_sc_hd__and3_1
XFILLER_33_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6510_ _7257_/Q _6510_/A2 _6510_/B1 _4164_/Y _6509_/X VGND VGND VPWR VPWR _6510_/X
+ sky130_fd_sc_hd__a221o_1
X_3722_ _6821_/Q _5331_/C _5440_/C _5458_/B _6970_/Q VGND VGND VPWR VPWR _3722_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6441_ _6431_/Y _6440_/Y _6691_/Q _6466_/A1 VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__o2bb2a_1
X_3653_ _6589_/Q _6530_/C _3446_/X _3488_/X hold59/A VGND VGND VPWR VPWR _3653_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6372_ _6565_/Q _6136_/A _6465_/A3 _6452_/B1 _6754_/Q VGND VGND VPWR VPWR _6372_/X
+ sky130_fd_sc_hd__a32o_1
X_3584_ input15/X _3504_/X _3509_/X _7160_/Q _3583_/X VGND VGND VPWR VPWR _3584_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5323_ _6850_/Q hold211/X _5323_/S VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5254_ hold16/A wire442/X _5253_/Y _5243_/Y VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__a211o_1
X_4205_ _4205_/A0 _4204_/X _4205_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5185_ _5040_/C _4293_/Y _5146_/D _4841_/B VGND VGND VPWR VPWR _5234_/B sky130_fd_sc_hd__o211a_1
XFILLER_29_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_6_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_4136_ _6539_/A0 hold957/X _4138_/S VGND VGND VPWR VPWR _4136_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4067_ _6549_/A0 hold992/X hold57/X VGND VGND VPWR VPWR _4067_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4969_ _4632_/A _4511_/A _4208_/Y _4293_/Y VGND VGND VPWR VPWR _5165_/B sky130_fd_sc_hd__a211o_1
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6708_ _7053_/CLK _6708_/D fanout601/X VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6639_ _6875_/CLK _6639_/D fanout598/X VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6990_ _7160_/CLK _6990_/D fanout592/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ _7021_/Q _7184_/Q _6072_/C _5783_/X _7013_/Q VGND VGND VPWR VPWR _5941_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_18_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5872_ _6906_/Q _5782_/C _5814_/C _6028_/B _6914_/Q VGND VGND VPWR VPWR _5872_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4823_ _4277_/Y _5040_/A _4403_/X _4358_/X VGND VGND VPWR VPWR _4827_/D sky130_fd_sc_hd__a211o_1
XFILLER_178_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4754_ _4755_/A _4754_/B _5036_/B VGND VGND VPWR VPWR _4754_/X sky130_fd_sc_hd__and3_1
X_3705_ _7026_/Q _5548_/C _6548_/D hold28/A _3704_/X VGND VGND VPWR VPWR _3705_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_147_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4685_ _4681_/Y _4685_/B _4685_/C _4685_/D VGND VGND VPWR VPWR _4685_/Y sky130_fd_sc_hd__nand4b_1
XFILLER_174_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3636_ _6660_/Q _3447_/X _3502_/X _6655_/Q _3635_/X VGND VGND VPWR VPWR _3636_/X
+ sky130_fd_sc_hd__a221o_1
X_6424_ _6562_/Q _6446_/B _6446_/C _6129_/B _6661_/Q VGND VGND VPWR VPWR _6424_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6355_ _6559_/Q _5750_/X _6454_/B1 _6768_/Q _6354_/X VGND VGND VPWR VPWR _6356_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3567_ _5512_/B _5657_/D hold28/A VGND VGND VPWR VPWR _5503_/B sky130_fd_sc_hd__and3_4
X_5306_ _6524_/B _5666_/C hold39/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__and3_2
XFILLER_88_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6286_ _7156_/Q _6129_/C _6269_/X _6270_/X VGND VGND VPWR VPWR _6286_/X sky130_fd_sc_hd__a211o_1
X_3498_ _6536_/C _5273_/D _6536_/D VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__and3_2
XFILLER_170_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5237_ _5060_/B _4449_/A _5143_/C _5236_/X VGND VGND VPWR VPWR _5238_/D sky130_fd_sc_hd__a31o_1
XFILLER_124_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5168_ _5165_/X _5247_/B _5064_/X _5085_/X VGND VGND VPWR VPWR _5168_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ hold24/X hold226/X _4120_/S VGND VGND VPWR VPWR _4119_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5099_ _4792_/C _5090_/X _4591_/B VGND VGND VPWR VPWR _5100_/C sky130_fd_sc_hd__a21oi_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__buf_6
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire360 _3889_/Y VGND VGND VPWR VPWR _3905_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4470_ _5060_/B _5060_/C _5143_/A _4859_/C VGND VGND VPWR VPWR _4476_/A sky130_fd_sc_hd__and4_1
Xwire371 _3834_/Y VGND VGND VPWR VPWR _3844_/B sky130_fd_sc_hd__clkbuf_2
Xhold407 _6772_/Q VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold418 _6955_/Q VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3421_ hold65/X hold37/X hold42/X hold28/A VGND VGND VPWR VPWR _5629_/C sky130_fd_sc_hd__and4_4
Xhold429 _5421_/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6140_ _7071_/Q _6446_/C _6425_/C VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__and3_1
XFILLER_112_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3352_ _6855_/Q _3352_/B VGND VGND VPWR VPWR _3352_/X sky130_fd_sc_hd__and2_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6672_/Q _5774_/X _5795_/X _6677_/Q _6070_/X VGND VGND VPWR VPWR _6071_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _6025_/B VGND VGND VPWR VPWR _5959_/C sky130_fd_sc_hd__inv_6
XFILLER_112_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _7063_/Q VGND VGND VPWR VPWR _5567_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5022_ _4474_/X _4786_/B _5263_/A _4561_/B _4586_/B VGND VGND VPWR VPWR _5022_/Y
+ sky130_fd_sc_hd__o2111ai_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 hold1364/X VGND VGND VPWR VPWR _5667_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 _7160_/Q VGND VGND VPWR VPWR _5677_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6973_ _7143_/CLK _6973_/D fanout588/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5924_ _7108_/Q _5764_/X _5784_/X _7028_/Q _5923_/X VGND VGND VPWR VPWR _5924_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5855_ _6969_/Q _5771_/X _5813_/X _7057_/Q VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
X_4806_ _4633_/Y _4735_/Y _4804_/X _4803_/Y _4166_/B VGND VGND VPWR VPWR _4806_/Y
+ sky130_fd_sc_hd__o221ai_1
X_5786_ _5934_/C _5786_/B VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__and2_1
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4737_ _4737_/A _4737_/B _4737_/C VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__nor3_1
XFILLER_119_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4668_ _4848_/B _4668_/B _4668_/C _4691_/B VGND VGND VPWR VPWR _4732_/C sky130_fd_sc_hd__and4_2
XFILLER_174_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6407_ _6660_/Q _6129_/B _6143_/X _6775_/Q _6406_/X VGND VGND VPWR VPWR _6414_/A
+ sky130_fd_sc_hd__a221o_1
X_3619_ _6649_/Q _3565_/X _5503_/B _7008_/Q _3618_/X VGND VGND VPWR VPWR _3619_/X
+ sky130_fd_sc_hd__a221o_1
Xhold930 _4018_/X VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold941 _6748_/Q VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _4633_/B _5036_/B VGND VGND VPWR VPWR _4599_/Y sky130_fd_sc_hd__nand2_1
Xhold952 _6667_/Q VGND VGND VPWR VPWR hold952/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold963 _4016_/X VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold974 hold974/A VGND VGND VPWR VPWR hold974/X sky130_fd_sc_hd__dlygate4sd3_1
X_6338_ _7046_/Q _6109_/X _6335_/X _6337_/X VGND VGND VPWR VPWR _6339_/C sky130_fd_sc_hd__a211o_1
Xhold985 _5364_/X VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 _6767_/Q VGND VGND VPWR VPWR hold996/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6269_ _7108_/Q _6117_/C _5750_/C _6110_/X _7116_/Q VGND VGND VPWR VPWR _6269_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3970_ hold758/X _5649_/A0 _3974_/S VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5640_ _6543_/A0 hold824/X hold9/X VGND VGND VPWR VPWR _5640_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5571_ hold5/X hold104/X _5574_/S VGND VGND VPWR VPWR _5571_/X sky130_fd_sc_hd__mux2_1
X_7310_ _7310_/A VGND VGND VPWR VPWR _7310_/X sky130_fd_sc_hd__buf_2
XFILLER_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4522_ _4313_/A _4747_/A _4544_/B _4544_/A VGND VGND VPWR VPWR _4522_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_117_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold204 _6950_/Q VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _5430_/X VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7241_ _7241_/CLK _7241_/D fanout576/X VGND VGND VPWR VPWR _7241_/Q sky130_fd_sc_hd__dfstp_1
Xhold226 _6746_/Q VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _4761_/C _4320_/A _4280_/A _4683_/B _4870_/B VGND VGND VPWR VPWR _4878_/C
+ sky130_fd_sc_hd__o311a_2
Xhold237 hold63/X VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold248 hold248/A VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ hold26/X hold71/X hold65/A VGND VGND VPWR VPWR _3404_/X sky130_fd_sc_hd__and3b_1
Xhold259 _5392_/X VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7172_ _7174_/CLK _7172_/D fanout608/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_1
X_4384_ _5143_/A _4449_/B _5143_/D VGND VGND VPWR VPWR _4461_/A sky130_fd_sc_hd__and3_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6176_/B _6143_/C _6104_/X _6451_/B1 _6122_/X VGND VGND VPWR VPWR _6134_/D
+ sky130_fd_sc_hd__a2111oi_4
X_3335_ _6851_/Q _6898_/Q _3346_/D _6718_/Q VGND VGND VPWR VPWR _3335_/X sky130_fd_sc_hd__o31a_1
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6600_/Q _6025_/B _6028_/B _5784_/X _6623_/Q VGND VGND VPWR VPWR _6054_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3266_ _7026_/Q VGND VGND VPWR VPWR _3266_/Y sky130_fd_sc_hd__inv_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5005_ _4738_/A _4859_/C _4704_/B _4723_/A VGND VGND VPWR VPWR _5005_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6956_ _7143_/CLK hold84/X fanout588/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5907_ _6875_/Q _5726_/Y _5894_/X _5906_/X _5759_/A VGND VGND VPWR VPWR _5907_/X
+ sky130_fd_sc_hd__o221a_1
X_6887_ _7135_/CLK _6887_/D fanout588/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5838_ _6872_/Q _5726_/Y _5824_/X _5837_/X _5759_/A VGND VGND VPWR VPWR _5838_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_167_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5769_ _7181_/Q _7180_/Q _6010_/D VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__and3_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold760 _6596_/Q VGND VGND VPWR VPWR hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _6929_/Q VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 _5366_/X VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold793 _4004_/X VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1460 _7250_/Q VGND VGND VPWR VPWR _7256_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1471 _6579_/Q VGND VGND VPWR VPWR _3569_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1482 _6627_/Q VGND VGND VPWR VPWR _3963_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3250__1 _3250__1/A VGND VGND VPWR VPWR _6512_/A3 sky130_fd_sc_hd__inv_2
Xhold1493 _7216_/Q VGND VGND VPWR VPWR _6393_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput309 _7314_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6810_ _7254_/CLK _6810_/D fanout613/X VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__dfrtp_4
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6741_ _6945_/CLK _6741_/D fanout583/X VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ _3905_/Y _3953_/A1 _3953_/S VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6672_ _7239_/CLK _6672_/D fanout574/X VGND VGND VPWR VPWR _6672_/Q sky130_fd_sc_hd__dfrtp_4
X_3884_ _6902_/Q _5377_/C _3521_/X _7174_/Q VGND VGND VPWR VPWR _3884_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5623_ _3918_/B hold484/X _5628_/S VGND VGND VPWR VPWR _5623_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5554_ _6505_/A1 hold826/X _5556_/S VGND VGND VPWR VPWR _5554_/X sky130_fd_sc_hd__mux2_1
X_4505_ _5060_/A _4505_/B _4597_/C VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__and3_1
XFILLER_172_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5485_ hold13/X _5485_/B _5629_/C VGND VGND VPWR VPWR _5493_/S sky130_fd_sc_hd__and3_4
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7224_ _7251_/CLK _7224_/D VGND VGND VPWR VPWR _7224_/Q sky130_fd_sc_hd__dfxtp_1
X_4436_ _5060_/C _5143_/A _4438_/D VGND VGND VPWR VPWR _4441_/B sky130_fd_sc_hd__and3_1
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout503 _6542_/A VGND VGND VPWR VPWR _5494_/A sky130_fd_sc_hd__buf_12
Xfanout514 hold86/X VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__buf_12
X_7155_ _7171_/CLK _7155_/D fanout609/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_4
X_4367_ _4662_/B _4246_/Y _4280_/A _4657_/C VGND VGND VPWR VPWR _4668_/B sky130_fd_sc_hd__o31ai_1
Xfanout525 hold2/X VGND VGND VPWR VPWR _3919_/C sky130_fd_sc_hd__buf_8
XFILLER_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout536 _7184_/Q VGND VGND VPWR VPWR _6072_/B sky130_fd_sc_hd__buf_12
X_3318_ _4229_/A _4229_/B _3318_/C _3318_/D VGND VGND VPWR VPWR _3319_/D sky130_fd_sc_hd__and4bb_1
XFILLER_98_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6106_ _7186_/Q _7185_/Q _6106_/C VGND VGND VPWR VPWR _6106_/X sky130_fd_sc_hd__and3_4
X_7086_ _7163_/CLK _7086_/D fanout608/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4298_ _5036_/C _4689_/B _4511_/A VGND VGND VPWR VPWR _4298_/X sky130_fd_sc_hd__and3_1
Xfanout569 _4754_/B VGND VGND VPWR VPWR _4549_/D sky130_fd_sc_hd__buf_4
XFILLER_86_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3249_/A VGND VGND VPWR VPWR _3249_/Y sky130_fd_sc_hd__inv_2
X_6037_ _7267_/Q _6025_/B wire398/X _5795_/X _6675_/Q VGND VGND VPWR VPWR _6037_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _7135_/CLK _6939_/D fanout588/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_csclk _3347_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_135_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold590 hold590/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1290 _7082_/Q VGND VGND VPWR VPWR _5588_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_430 _6109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5270_ _5269_/X _5270_/B _5270_/C _5270_/D VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__and4b_1
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4221_ _4228_/C _4228_/D _4227_/A _4227_/B VGND VGND VPWR VPWR _4222_/B sky130_fd_sc_hd__nand4_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4152_ _6542_/A _4152_/B _4152_/C VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__and3_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4083_ _4083_/A0 _4082_/X _4093_/S VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4985_ _5255_/A _4804_/C _4659_/B _4857_/C _4987_/C VGND VGND VPWR VPWR _4985_/Y
+ sky130_fd_sc_hd__a32oi_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6724_ _6957_/CLK _6724_/D fanout591/X VGND VGND VPWR VPWR _7286_/A sky130_fd_sc_hd__dfrtp_1
X_3936_ _3934_/S hold796/X _3432_/X _3919_/X VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6655_ _6828_/CLK _6655_/D fanout573/X VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfstp_2
X_3867_ _7109_/Q _6536_/A _5281_/A2 _3452_/X _6965_/Q VGND VGND VPWR VPWR _3867_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5606_ hold24/X _5606_/A1 _5610_/S VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__mux2_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6586_ _7256_/CLK _6586_/D VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfxtp_1
X_3798_ input16/X _3528_/X _3559_/X _6907_/Q _3755_/X VGND VGND VPWR VPWR _3798_/X
+ sky130_fd_sc_hd__a221o_1
X_5537_ hold716/X _4051_/B _5538_/S VGND VGND VPWR VPWR _5537_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5468_ _5649_/A0 _5468_/A1 _5475_/S VGND VGND VPWR VPWR _5468_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7207_ _7219_/CLK _7207_/D fanout595/X VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfrtp_1
X_4419_ _4277_/Y _4358_/X _4403_/X _4415_/X _4391_/Y VGND VGND VPWR VPWR _5241_/C
+ sky130_fd_sc_hd__o32a_1
X_5399_ hold146/X _3922_/C _5403_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7138_ _7165_/CLK _7138_/D fanout602/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout377 _4521_/Y VGND VGND VPWR VPWR _5263_/A sky130_fd_sc_hd__buf_4
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7069_ _7093_/CLK _7069_/D fanout593/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _3969_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 _3536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_282 _5723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_293 _5777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4770_ _4598_/Y _4640_/Y _4769_/Y _4768_/Y VGND VGND VPWR VPWR _4773_/C sky130_fd_sc_hd__o211ai_1
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3721_ _6728_/Q hold38/A _3721_/A3 _3719_/X _3720_/X VGND VGND VPWR VPWR _3721_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6440_ _6440_/A _6440_/B _6440_/C _6440_/D VGND VGND VPWR VPWR _6440_/Y sky130_fd_sc_hd__nor4_1
XFILLER_174_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3652_ _3652_/A _3652_/B _3652_/C _3652_/D VGND VGND VPWR VPWR _3652_/Y sky130_fd_sc_hd__nor4_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3583_ _6603_/Q _5666_/C _4139_/C _3433_/X _6936_/Q VGND VGND VPWR VPWR _3583_/X
+ sky130_fd_sc_hd__a32o_1
X_6371_ _6659_/Q _6129_/B _6143_/X _6774_/Q _6370_/X VGND VGND VPWR VPWR _6371_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5322_ _3916_/C hold344/X _5322_/S VGND VGND VPWR VPWR _5322_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ _5249_/X _5252_/Y _5247_/Y VGND VGND VPWR VPWR _5253_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4204_ hold565/X _4053_/X _4204_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
X_5184_ _5238_/A _5238_/C _5184_/C VGND VGND VPWR VPWR _5187_/A sky130_fd_sc_hd__nor3_1
X_4135_ _6538_/A0 hold442/X _4138_/S VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_63_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7148_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4066_ _5620_/A _6548_/B hold56/X _5675_/D VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__nand4_4
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6835_/CLK sky130_fd_sc_hd__clkbuf_16
X_4968_ _4632_/B _4970_/D _4480_/B _4967_/X VGND VGND VPWR VPWR _4973_/A sky130_fd_sc_hd__a31o_1
X_6707_ _7168_/CLK _6707_/D fanout609/X VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfrtp_1
X_3919_ _5494_/A hold64/X _3919_/C VGND VGND VPWR VPWR _3919_/X sky130_fd_sc_hd__and3_4
XFILLER_149_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4899_ _5263_/A _4746_/A _5173_/C _4589_/B _4557_/X VGND VGND VPWR VPWR _4899_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6638_ _7269_/CLK _6638_/D fanout576/X VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6569_ _6687_/CLK _6569_/D fanout580/X VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7271_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire553 _4799_/C VGND VGND VPWR VPWR _4748_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5940_ _7085_/Q _5826_/B _6009_/C _5788_/X hold79/A VGND VGND VPWR VPWR _5940_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5871_ _7066_/Q _5723_/X _5773_/X _7034_/Q _5870_/X VGND VGND VPWR VPWR _5871_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4822_ _4277_/Y _4398_/X _4403_/X _4414_/X _4299_/Y VGND VGND VPWR VPWR _4829_/B
+ sky130_fd_sc_hd__o32a_1
X_4753_ _4753_/A _4753_/B VGND VGND VPWR VPWR _4755_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3704_ _6567_/Q _3368_/X _5548_/C _3547_/X _7034_/Q VGND VGND VPWR VPWR _3704_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4684_ _4939_/A _4849_/A _5255_/A _4878_/C VGND VGND VPWR VPWR _4685_/C sky130_fd_sc_hd__nand4_1
XFILLER_147_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6423_ _7247_/Q _6103_/X _6117_/X _6595_/Q _6422_/X VGND VGND VPWR VPWR _6423_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3635_ _6913_/Q _4158_/D _5281_/A2 _3492_/X _6665_/Q VGND VGND VPWR VPWR _3635_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6354_ _6587_/Q _6138_/A _6110_/C _6137_/X _7270_/Q VGND VGND VPWR VPWR _6354_/X
+ sky130_fd_sc_hd__a32o_1
X_3566_ _5512_/B _5630_/C hold28/A VGND VGND VPWR VPWR _5557_/B sky130_fd_sc_hd__and3_4
X_5305_ _5305_/A0 _5649_/A0 _5305_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3497_ _6524_/A _5327_/D _6536_/D VGND VGND VPWR VPWR _3497_/X sky130_fd_sc_hd__and3_2
X_6285_ _6285_/A _6285_/B VGND VGND VPWR VPWR _6285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5236_ _5060_/B _5060_/C _5133_/X _4813_/X VGND VGND VPWR VPWR _5236_/X sky130_fd_sc_hd__a31o_1
XFILLER_124_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5167_ _4480_/B _4718_/D _5166_/X VGND VGND VPWR VPWR _5247_/B sky130_fd_sc_hd__a21oi_1
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4118_ _3918_/B hold743/X _4120_/S VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__mux2_1
X_5098_ _5098_/A _5177_/C VGND VGND VPWR VPWR _5101_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4049_ hold65/X _4049_/B VGND VGND VPWR VPWR _4049_/X sky130_fd_sc_hd__and2_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire350 _3692_/Y VGND VGND VPWR VPWR _3693_/B sky130_fd_sc_hd__clkbuf_1
Xwire361 _3874_/Y VGND VGND VPWR VPWR _3875_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire372 _3523_/Y VGND VGND VPWR VPWR _3568_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_171_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold408 _4150_/X VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold419 _5445_/X VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3420_ hold26/X hold71/X hold65/A VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__o21ai_4
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3351_ input1/X _3351_/B VGND VGND VPWR VPWR _3351_/X sky130_fd_sc_hd__and2_2
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3282_/A VGND VGND VPWR VPWR _3282_/Y sky130_fd_sc_hd__inv_2
X_6070_ _6687_/Q _5768_/X _5814_/X _6591_/Q VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__a22o_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _5567_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5021_ _4786_/B _4561_/B _4581_/B _4910_/X _4562_/B VGND VGND VPWR VPWR _5174_/C
+ sky130_fd_sc_hd__a311oi_2
Xhold1119 _7265_/Q VGND VGND VPWR VPWR _6537_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6972_ _7015_/CLK _6972_/D fanout588/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5923_ _7076_/Q _5971_/A2 _5813_/X _7060_/Q _5922_/X VGND VGND VPWR VPWR _5923_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5854_ _6937_/Q _5782_/X _5852_/X _5934_/C _5853_/X VGND VGND VPWR VPWR _5854_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4805_ _4799_/C _4734_/X _7257_/Q _7258_/Q _7259_/Q VGND VGND VPWR VPWR _4805_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5785_ _6887_/Q _5795_/C _5815_/C _6028_/B _6911_/Q VGND VGND VPWR VPWR _5786_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_166_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4736_ _5128_/A _5128_/C _4923_/B VGND VGND VPWR VPWR _4737_/B sky130_fd_sc_hd__and3_1
XFILLER_159_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4667_ _4939_/A _4984_/B _4667_/C _4667_/D VGND VGND VPWR VPWR _4667_/Y sky130_fd_sc_hd__nand4_1
X_6406_ _6645_/Q _6444_/C wire392/A _6116_/X _6571_/Q VGND VGND VPWR VPWR _6406_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold920 _5678_/X VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3618_ _6928_/Q _5413_/B _3562_/X _6639_/Q _3617_/X VGND VGND VPWR VPWR _3618_/X
+ sky130_fd_sc_hd__a221o_1
Xhold931 _6890_/Q VGND VGND VPWR VPWR _3282_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4598_ _4494_/C _4754_/B _5036_/B VGND VGND VPWR VPWR _4598_/Y sky130_fd_sc_hd__nand3b_1
Xhold942 _4122_/X VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold953 _4010_/X VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6337_ _7118_/Q _6110_/X _6135_/X _6942_/Q _6336_/X VGND VGND VPWR VPWR _6337_/X
+ sky130_fd_sc_hd__a221o_1
Xhold964 _7134_/Q VGND VGND VPWR VPWR hold964/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold975 hold975/A VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlygate4sd3_1
X_3549_ _7047_/Q _3563_/A _3540_/B _3547_/X _7031_/Q VGND VGND VPWR VPWR _3549_/X
+ sky130_fd_sc_hd__a32o_1
Xhold986 _6597_/Q VGND VGND VPWR VPWR hold986/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold997 _4144_/X VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6268_ _6267_/X _6268_/A1 _6443_/S VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5219_ _4751_/A _4592_/B _4903_/A _4595_/A _5218_/X VGND VGND VPWR VPWR _5220_/D
+ sky130_fd_sc_hd__a221oi_1
X_6199_ hold59/A _6446_/C _6425_/C _6126_/X _6961_/Q VGND VGND VPWR VPWR _6199_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_29_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5570_ _3921_/B hold340/X _5574_/S VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4318_/A _4318_/B _4317_/Y VGND VGND VPWR VPWR _4521_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold205 _5439_/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7240_ _7240_/CLK _7240_/D fanout596/X VGND VGND VPWR VPWR _7240_/Q sky130_fd_sc_hd__dfrtp_2
Xhold216 _7142_/Q VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _4848_/A _4356_/A _4382_/Y _4295_/A _4349_/X VGND VGND VPWR VPWR _4456_/B
+ sky130_fd_sc_hd__a2111o_1
Xhold227 _4119_/X VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _5315_/X VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold249 _7051_/Q VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3403_ _6472_/A _7251_/Q VGND VGND VPWR VPWR _3906_/S sky130_fd_sc_hd__nand2_4
X_7171_ _7171_/CLK hold6/X fanout609/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_4
X_4383_ _4383_/A _4984_/A _4870_/B VGND VGND VPWR VPWR _4449_/B sky130_fd_sc_hd__and3_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6177_/A _6143_/C _6177_/C VGND VGND VPWR VPWR _6122_/X sky130_fd_sc_hd__and3_4
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _6723_/Q input77/X _3349_/A VGND VGND VPWR VPWR _3334_/X sky130_fd_sc_hd__mux2_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6053_ _6666_/Q _6028_/B _6072_/C _6681_/Q _6025_/B VGND VGND VPWR VPWR _6053_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _7034_/Q VGND VGND VPWR VPWR _3265_/Y sky130_fd_sc_hd__inv_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5128_/B _4945_/B _4675_/B _4719_/B _4788_/A VGND VGND VPWR VPWR _5007_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_39_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6955_ _7063_/CLK _6955_/D fanout590/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5906_ _7059_/Q _5813_/X _5898_/X _5902_/X _5905_/X VGND VGND VPWR VPWR _5906_/X
+ sky130_fd_sc_hd__a2111o_1
X_6886_ _6908_/CLK _6886_/D fanout609/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5837_ _7096_/Q _5780_/X _5829_/X _5833_/X _5836_/X VGND VGND VPWR VPWR _5837_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_179_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5768_ _5783_/C _5795_/D _5815_/B VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__and3_4
XFILLER_182_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4719_ _4788_/A _4719_/B VGND VGND VPWR VPWR _4720_/C sky130_fd_sc_hd__nand2_1
X_5699_ _6442_/S _3300_/B _6803_/Q _5697_/Y VGND VGND VPWR VPWR _5711_/A sky130_fd_sc_hd__a211o_1
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold750 _7138_/Q VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold761 _3926_/X VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _5416_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _6928_/Q VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1450 _7277_/Q VGND VGND VPWR VPWR hold959/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _7226_/Q VGND VGND VPWR VPWR _6478_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 _7227_/Q VGND VGND VPWR VPWR _6479_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1483 _6943_/Q VGND VGND VPWR VPWR hold1483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1494 _6614_/Q VGND VGND VPWR VPWR _3948_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6740_ _6835_/CLK _6740_/D fanout583/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfstp_4
X_3952_ _3875_/Y _3952_/A1 _3953_/S VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6671_ _6780_/CLK _6671_/D _3291_/A VGND VGND VPWR VPWR _6671_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3883_ _7126_/Q _3525_/X _3539_/X input60/X _3882_/X VGND VGND VPWR VPWR _3889_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5622_ _6550_/A0 hold712/X _5628_/S VGND VGND VPWR VPWR _5622_/X sky130_fd_sc_hd__mux2_1
X_5553_ _3924_/B hold249/X _5556_/S VGND VGND VPWR VPWR _5553_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4504_ _4504_/A _4504_/B _4504_/C VGND VGND VPWR VPWR _4504_/Y sky130_fd_sc_hd__nand3_1
XFILLER_144_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5484_ _4053_/B hold209/X _5484_/S VGND VGND VPWR VPWR _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7223_ _7259_/CLK _7223_/D VGND VGND VPWR VPWR _7223_/Q sky130_fd_sc_hd__dfxtp_1
X_4435_ _4427_/C _4429_/D _4277_/Y _4383_/A VGND VGND VPWR VPWR _4435_/X sky130_fd_sc_hd__a211o_1
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout504 hold12/X VGND VGND VPWR VPWR _6542_/A sky130_fd_sc_hd__buf_12
X_7154_ _7154_/CLK _7154_/D fanout593/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout515 _3925_/C VGND VGND VPWR VPWR _6535_/A0 sky130_fd_sc_hd__buf_8
XFILLER_160_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4366_ _4662_/B _4246_/Y _4280_/A _4870_/B VGND VGND VPWR VPWR _4654_/B sky130_fd_sc_hd__o31ai_4
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout526 hold2/X VGND VGND VPWR VPWR _3918_/B sky130_fd_sc_hd__buf_12
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout537 _6059_/S VGND VGND VPWR VPWR _5826_/B sky130_fd_sc_hd__buf_8
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6105_ _6117_/A _6136_/A _6177_/C VGND VGND VPWR VPWR _6105_/X sky130_fd_sc_hd__and3_4
X_3317_ _3317_/A _3317_/B _3317_/C VGND VGND VPWR VPWR _3318_/D sky130_fd_sc_hd__and3_1
Xfanout548 _4939_/B VGND VGND VPWR VPWR _4945_/C sky130_fd_sc_hd__buf_6
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7085_ _7148_/CLK _7085_/D fanout592/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout559 _4945_/B VGND VGND VPWR VPWR _5128_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_98_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4297_ _4612_/C _4600_/B VGND VGND VPWR VPWR _4753_/A sky130_fd_sc_hd__nand2b_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _7246_/Q _6025_/B _5723_/X _6025_/X _6035_/X VGND VGND VPWR VPWR _6036_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_86_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3248_ _6850_/Q VGND VGND VPWR VPWR _5694_/A sky130_fd_sc_hd__inv_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7152_/CLK _6938_/D fanout586/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _7071_/CLK _6869_/D fanout585/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold580 hold580/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_1_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold591 _6600_/Q VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1280 _7302_/A VGND VGND VPWR VPWR _4070_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 _6988_/Q VGND VGND VPWR VPWR _5482_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_420 _3918_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_431 _6425_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4220_ _4227_/C _4227_/D _4656_/C VGND VGND VPWR VPWR _4222_/A sky130_fd_sc_hd__nand3_1
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4151_ _6536_/B _4152_/C VGND VGND VPWR VPWR _4156_/S sky130_fd_sc_hd__nand2_2
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4082_ hold295/X _3918_/X _4092_/S VGND VGND VPWR VPWR _4082_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4984_ _4984_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _4987_/C sky130_fd_sc_hd__and3_2
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6723_ _7063_/CLK _6723_/D fanout584/X VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfrtp_2
X_3935_ _3934_/S hold787/X _3432_/X _3916_/X VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6654_ _6843_/CLK _6654_/D fanout584/X VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfrtp_4
X_3866_ _6973_/Q _5458_/B _3536_/X _6989_/Q _3865_/X VGND VGND VPWR VPWR _3873_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5605_ _3918_/B hold682/X _5610_/S VGND VGND VPWR VPWR _5605_/X sky130_fd_sc_hd__mux2_1
X_6585_ _7256_/CLK _6585_/D VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3797_ _6637_/Q _3969_/C _3794_/X _3796_/X VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__a211o_1
XFILLER_118_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5536_ hold868/X _6505_/A1 _5538_/S VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5467_ _5476_/B hold66/A _5485_/B _5575_/D VGND VGND VPWR VPWR _5475_/S sky130_fd_sc_hd__nand4_4
X_7206_ _7237_/CLK _7206_/D fanout578/X VGND VGND VPWR VPWR _7206_/Q sky130_fd_sc_hd__dfrtp_4
X_4418_ _4751_/A _5060_/B _5055_/D _4475_/B VGND VGND VPWR VPWR _4418_/X sky130_fd_sc_hd__and4_1
X_5398_ hold280/X _3919_/C _5403_/S VGND VGND VPWR VPWR _5398_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7137_ _7156_/CLK _7137_/D fanout602/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4349_ _4243_/A _4243_/B _4277_/Y _4346_/Y VGND VGND VPWR VPWR _4349_/X sky130_fd_sc_hd__a211o_2
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout378 _4862_/A VGND VGND VPWR VPWR _5255_/A sky130_fd_sc_hd__buf_4
X_7068_ _7171_/CLK _7068_/D fanout611/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6019_ _6759_/Q _5771_/X _6002_/X _6004_/X _6018_/X VGND VGND VPWR VPWR _6019_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_250 hold89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 _3433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 _3536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 _5723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_294 _5779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _7242_/Q _6536_/A _5325_/C _3564_/X _7268_/Q VGND VGND VPWR VPWR _3720_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3651_ _6905_/Q _3559_/X _3644_/X _3646_/X _3650_/X VGND VGND VPWR VPWR _3652_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6370_ _6649_/Q _6177_/A _6106_/C _6451_/B1 _6664_/Q VGND VGND VPWR VPWR _6370_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3582_ input62/X _5334_/B _3576_/X _3577_/X _3581_/X VGND VGND VPWR VPWR _3582_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_127_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5321_ _4051_/B hold583/X _5322_/S VGND VGND VPWR VPWR _5321_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ _4659_/B _4950_/X _5152_/X _5251_/X VGND VGND VPWR VPWR _5252_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_114_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4203_ _4203_/A0 _4202_/X _4205_/S VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5183_ _5040_/X _4414_/X _5182_/X _5142_/B VGND VGND VPWR VPWR _5184_/C sky130_fd_sc_hd__o211ai_1
X_4134_ _3370_/B hold943/X _4138_/S VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4065_ _4053_/X hold565/X _4065_/S VGND VGND VPWR VPWR _4065_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4967_ _4788_/A _4950_/X _4966_/Y _4938_/X VGND VGND VPWR VPWR _4967_/X sky130_fd_sc_hd__a211o_1
XFILLER_149_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3918_ hold65/X _3918_/B VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__and2_4
X_6706_ _7140_/CLK _6706_/D fanout609/X VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4898_ _4640_/A _4774_/B _4570_/B VGND VGND VPWR VPWR _4898_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6637_ _7035_/CLK _6637_/D fanout590/X VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3849_ input32/X _3504_/X _3544_/X _6949_/Q _3848_/X VGND VGND VPWR VPWR _3856_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_20_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6568_ _6781_/CLK _6568_/D _3291_/A VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5519_ hold21/X hold184/X _5520_/S VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__mux2_1
X_6499_ _6498_/X hold24/A _6511_/S VGND VGND VPWR VPWR _7232_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5870_ _7082_/Q _6010_/D _5815_/C _5795_/D VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__a31o_1
XFILLER_61_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4821_ _4299_/Y _4380_/X _4403_/X _4412_/Y _4349_/X VGND VGND VPWR VPWR _4829_/A
+ sky130_fd_sc_hd__o32a_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4752_ _4752_/A _4752_/B _4752_/C _4752_/D VGND VGND VPWR VPWR _4752_/Y sky130_fd_sc_hd__nand4_1
XFILLER_187_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3703_ _7122_/Q _3525_/X _3544_/X _6946_/Q _3702_/X VGND VGND VPWR VPWR _3703_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4683_ _4849_/A _4683_/B _4683_/C VGND VGND VPWR VPWR _4683_/X sky130_fd_sc_hd__and3_1
X_6422_ _6572_/Q _6116_/X _6129_/D _6671_/Q VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__a22o_1
X_3634_ _3987_/A _5657_/D _5313_/D VGND VGND VPWR VPWR _3634_/X sky130_fd_sc_hd__and3_1
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6353_ _6758_/Q _6097_/X _6101_/X _6683_/Q _6352_/X VGND VGND VPWR VPWR _6356_/C
+ sky130_fd_sc_hd__a221o_1
X_3565_ _3987_/A _6548_/A _5657_/D VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__and3_2
X_5304_ _5304_/A _5476_/B _5311_/C _6524_/B VGND VGND VPWR VPWR _5305_/S sky130_fd_sc_hd__and4_1
X_6284_ _7132_/Q _6116_/X _6276_/X _6280_/X _6283_/X VGND VGND VPWR VPWR _6285_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3496_ _5630_/C _5485_/B hold28/A VGND VGND VPWR VPWR _3496_/X sky130_fd_sc_hd__and3_4
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5235_ _4843_/B _5235_/B _5235_/C _5235_/D VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__and4b_1
XFILLER_69_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5166_ _4939_/A _4792_/A _5128_/C _4799_/X _4973_/C VGND VGND VPWR VPWR _5166_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_29_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4117_ _6538_/A0 hold385/X _4120_/S VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5097_ _4778_/C _5090_/X _4922_/B _4582_/A _5027_/B VGND VGND VPWR VPWR _5177_/C
+ sky130_fd_sc_hd__a2111o_1
X_4048_ hold369/X _3924_/B _4054_/S VGND VGND VPWR VPWR _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5999_ _6688_/Q _5726_/Y _5987_/X _5998_/X _5759_/A VGND VGND VPWR VPWR _5999_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput290 _6736_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_160_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__buf_6
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire351 _3652_/Y VGND VGND VPWR VPWR _3693_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_62_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7160_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire362 _3843_/Y VGND VGND VPWR VPWR _3844_/C sky130_fd_sc_hd__clkbuf_2
Xhold409 _6987_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3350_ _3350_/A _3350_/B VGND VGND VPWR VPWR _3350_/X sky130_fd_sc_hd__and2_2
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7067_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3281_/A VGND VGND VPWR VPWR _3281_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5020_ _5094_/A _5222_/D _5020_/C _5020_/D VGND VGND VPWR VPWR _5024_/B sky130_fd_sc_hd__and4b_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1109 _6855_/Q VGND VGND VPWR VPWR _5332_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6971_ _7071_/CLK hold62/X fanout585/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__dfrtp_4
X_5922_ _7044_/Q _5826_/B _5959_/B _5970_/B1 _6932_/Q VGND VGND VPWR VPWR _5922_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_179_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ _5795_/D _5782_/C _5795_/C _6086_/B1 _7105_/Q VGND VGND VPWR VPWR _5853_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4804_ _4804_/A _5128_/C _4804_/C VGND VGND VPWR VPWR _4804_/X sky130_fd_sc_hd__and3_1
X_5784_ _6059_/S _7181_/Q _7180_/Q _5815_/B VGND VGND VPWR VPWR _5784_/X sky130_fd_sc_hd__and4_4
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4735_ _4804_/A _5128_/C VGND VGND VPWR VPWR _4735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4666_ _5128_/B _5128_/C _4665_/Y _4661_/X VGND VGND VPWR VPWR _4666_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6405_ _6405_/A _6405_/B _6405_/C _6405_/D VGND VGND VPWR VPWR _6415_/B sky130_fd_sc_hd__nor4_1
XFILLER_134_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3617_ _7064_/Q _5512_/B hold39/A _3616_/X VGND VGND VPWR VPWR _3617_/X sky130_fd_sc_hd__a31o_1
XFILLER_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold910 _5574_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 _6880_/Q VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ _4606_/B _4597_/B _4597_/C _4923_/A VGND VGND VPWR VPWR _4604_/B sky130_fd_sc_hd__nand4_1
Xhold932 _6845_/Q VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _6758_/Q VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 hold954/A VGND VGND VPWR VPWR hold954/X sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ _7038_/Q _6138_/B _6108_/X _6137_/X _7102_/Q VGND VGND VPWR VPWR _6336_/X
+ sky130_fd_sc_hd__a32o_1
X_3548_ _5620_/A _3563_/A _5548_/D VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__and3_4
XFILLER_115_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold965 _5647_/X VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold976 _6677_/Q VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold987 _3928_/X VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold998 _6645_/Q VGND VGND VPWR VPWR hold998/X sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ _6292_/S _7210_/Q _6265_/Y _6266_/X VGND VGND VPWR VPWR _6267_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3479_ _3987_/A _5620_/A _5684_/B VGND VGND VPWR VPWR _5334_/B sky130_fd_sc_hd__and3_4
XFILLER_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5218_ _4595_/A _4923_/A _5263_/B _4596_/A VGND VGND VPWR VPWR _5218_/X sky130_fd_sc_hd__a31o_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6198_ _7121_/Q _5750_/X _6107_/X _7001_/Q _6197_/X VGND VGND VPWR VPWR _6205_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_97_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5149_ _4266_/Y _4503_/X _5149_/C _5149_/D VGND VGND VPWR VPWR _5235_/D sky130_fd_sc_hd__and4bb_1
XFILLER_84_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4520_ _4214_/A _4214_/B _4313_/A _4747_/A VGND VGND VPWR VPWR _4544_/B sky130_fd_sc_hd__a22oi_4
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold206 hold206/A VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _4451_/A _4451_/B VGND VGND VPWR VPWR _4456_/A sky130_fd_sc_hd__nor2_1
Xhold217 _5656_/X VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _6861_/Q VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 hold239/A VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _3924_/B hold786/X _3402_/S VGND VGND VPWR VPWR _3402_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7170_ _7170_/CLK _7170_/D fanout605/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4382_ _4383_/A _4870_/B VGND VGND VPWR VPWR _4382_/Y sky130_fd_sc_hd__nand2_2
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6121_ _7185_/Q _6143_/D _6141_/B _6143_/C VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__and4b_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3333_ _6860_/Q input81/X _3350_/A VGND VGND VPWR VPWR _3333_/X sky130_fd_sc_hd__mux2_4
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _7247_/Q _5723_/X _6003_/C _6610_/Q _6028_/C VGND VGND VPWR VPWR _6052_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3264_ _7042_/Q VGND VGND VPWR VPWR _3264_/Y sky130_fd_sc_hd__inv_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5003_/A _5194_/A _5003_/C _5228_/B VGND VGND VPWR VPWR _5007_/B sky130_fd_sc_hd__nand4_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6954_ _7156_/CLK _6954_/D fanout602/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_4
X_5905_ hold61/A _5771_/X _5888_/X _5891_/X _5904_/X VGND VGND VPWR VPWR _5905_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_81_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6885_ _7160_/CLK _6885_/D fanout592/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5836_ _6968_/Q _5771_/X _5818_/X _5821_/X _5835_/X VGND VGND VPWR VPWR _5836_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_22_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5767_ _6059_/S _7183_/Q _7182_/Q _5815_/C VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__and4_4
XFILLER_163_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4718_ _4859_/A _4984_/C _4788_/A _4718_/D VGND VGND VPWR VPWR _4720_/B sky130_fd_sc_hd__nand4_1
X_5698_ _3300_/B _6292_/S _6803_/Q VGND VGND VPWR VPWR _5698_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_175_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _4940_/C _4789_/B _4945_/C VGND VGND VPWR VPWR _4719_/B sky130_fd_sc_hd__and3_4
XFILLER_135_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold740 _5682_/X VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold751 _5652_/X VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold762 hold762/A VGND VGND VPWR VPWR hold762/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold773 _6655_/Q VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold784 _6649_/Q VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ _7086_/Q _6177_/A _6102_/X _6130_/X _6934_/Q VGND VGND VPWR VPWR _6319_/X
+ sky130_fd_sc_hd__a32o_1
X_7299_ _7299_/A VGND VGND VPWR VPWR _7299_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold795 _5415_/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1440 _6804_/Q VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1451 _6551_/X VGND VGND VPWR VPWR _7277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1462 _6976_/Q VGND VGND VPWR VPWR hold148/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1473 _7085_/Q VGND VGND VPWR VPWR hold841/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 _6618_/Q VGND VGND VPWR VPWR _3952_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _7195_/Q VGND VGND VPWR VPWR _5861_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3951_ _3844_/Y _3951_/A1 _3953_/S VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6670_ _6827_/CLK _6670_/D fanout574/X VGND VGND VPWR VPWR _6670_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3882_ input51/X _3368_/X hold56/A _3463_/X _7118_/Q VGND VGND VPWR VPWR _3882_/X
+ sky130_fd_sc_hd__a32o_1
X_5621_ _6549_/A0 _5621_/A1 _5628_/S VGND VGND VPWR VPWR _5621_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5552_ _3921_/B hold330/X _5556_/S VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4503_ _4505_/B _4804_/A _4804_/C VGND VGND VPWR VPWR _4503_/X sky130_fd_sc_hd__and3_1
X_5483_ _4051_/B hold463/X _5484_/S VGND VGND VPWR VPWR _5483_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7222_ _7259_/CLK _7222_/D VGND VGND VPWR VPWR _7222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4434_ _4247_/Y _4248_/X _4984_/A _4256_/Y VGND VGND VPWR VPWR _4438_/D sky130_fd_sc_hd__o211a_1
XFILLER_172_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7153_ _7165_/CLK _7153_/D fanout601/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4365_ _4662_/B _4246_/Y _4280_/A _4870_/B VGND VGND VPWR VPWR _4683_/C sky130_fd_sc_hd__o31a_1
Xfanout505 hold12/X VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__buf_12
Xfanout516 hold5/X VGND VGND VPWR VPWR _3925_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout527 hold35/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__buf_12
X_6104_ _6117_/A _6130_/A _6138_/B VGND VGND VPWR VPWR _6104_/X sky130_fd_sc_hd__and3_4
X_3316_ _4227_/C _4227_/D _3316_/C VGND VGND VPWR VPWR _3317_/C sky130_fd_sc_hd__nor3_1
Xfanout538 _6059_/S VGND VGND VPWR VPWR _5965_/B sky130_fd_sc_hd__buf_4
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7084_ _7168_/CLK _7084_/D fanout608/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout549 _4637_/Y VGND VGND VPWR VPWR _4939_/B sky130_fd_sc_hd__buf_6
XFILLER_58_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4296_ _4612_/C _4600_/B VGND VGND VPWR VPWR _5036_/C sky130_fd_sc_hd__and2b_4
X_6035_ _6589_/Q _5814_/X _5815_/X _6640_/Q _6034_/X VGND VGND VPWR VPWR _6035_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3247_ _4747_/A VGND VGND VPWR VPWR _4760_/B sky130_fd_sc_hd__clkinv_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6937_ _7067_/CLK _6937_/D fanout582/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6868_ _7077_/CLK _6868_/D fanout591/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5819_ _6912_/Q _6028_/B _5934_/C VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__and3_1
X_6799_ _7168_/CLK _6799_/D fanout608/X VGND VGND VPWR VPWR _7298_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_10_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold570 _4060_/X VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold581 hold581/A VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold592 _3931_/X VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1270 _6475_/A1 VGND VGND VPWR VPWR hold676/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1281 _7131_/Q VGND VGND VPWR VPWR _5644_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 _7171_/Q VGND VGND VPWR VPWR _5689_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_410 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_421 hold64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_432 _6446_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4150_ hold407/X _3925_/C _4150_/S VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4081_ _4081_/A0 _4080_/X _4093_/S VGND VGND VPWR VPWR _4081_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4983_ _4678_/A _4983_/B _4983_/C VGND VGND VPWR VPWR _5120_/B sky130_fd_sc_hd__and3b_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6722_ _7148_/CLK _6722_/D fanout591/X VGND VGND VPWR VPWR _7285_/A sky130_fd_sc_hd__dfrtp_1
X_3934_ _4152_/B _3934_/A1 _3934_/S VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3865_ _7085_/Q _6536_/A _5440_/C _3571_/X _6731_/Q VGND VGND VPWR VPWR _3865_/X
+ sky130_fd_sc_hd__a32o_1
X_6653_ _7265_/CLK _6653_/D fanout575/X VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5604_ _6550_/A0 hold783/X _5610_/S VGND VGND VPWR VPWR _5604_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3796_ _7147_/Q _3474_/X _3502_/X _6657_/Q _3795_/X VGND VGND VPWR VPWR _3796_/X
+ sky130_fd_sc_hd__a221o_1
X_6584_ _7256_/CLK _6584_/D VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5535_ hold142/X hold5/X _5538_/S VGND VGND VPWR VPWR _5535_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5466_ _4053_/B hold198/X _5466_/S VGND VGND VPWR VPWR _5466_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7205_ _7218_/CLK _7205_/D fanout594/X VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4417_ _4734_/B _4416_/A _4670_/D _4416_/Y VGND VGND VPWR VPWR _4475_/B sky130_fd_sc_hd__o211a_2
XFILLER_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5397_ hold398/X _3916_/C _5403_/S VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7136_ _7156_/CLK _7136_/D fanout603/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfstp_1
X_4348_ _4214_/A _4214_/B _4284_/A _4488_/B VGND VGND VPWR VPWR _4348_/X sky130_fd_sc_hd__a211o_2
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7067_ _7067_/CLK _7067_/D fanout584/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_4
X_4279_ _4698_/A _4657_/C _4656_/C _4647_/C VGND VGND VPWR VPWR _4280_/B sky130_fd_sc_hd__nand4_2
Xfanout379 _4375_/X VGND VGND VPWR VPWR _4862_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6018_ _6774_/Q _5779_/X _5782_/X _6654_/Q _6017_/X VGND VGND VPWR VPWR _6018_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_240 hold2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 hold89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 _3446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_273 _3544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_284 _5764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 _5783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3650_ input37/X _4187_/S _3649_/X _3634_/X _3648_/X VGND VGND VPWR VPWR _3650_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3581_ _6904_/Q _3559_/X _3572_/X _3579_/X _3580_/X VGND VGND VPWR VPWR _3581_/X
+ sky130_fd_sc_hd__a2111o_1
X_5320_ hold83/X hold140/X _5322_/S VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5251_ _4716_/A _4945_/C _4903_/B _5066_/X _5250_/X VGND VGND VPWR VPWR _5251_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4202_ hold599/X _4051_/X _4204_/S VGND VGND VPWR VPWR _4202_/X sky130_fd_sc_hd__mux2_1
X_5182_ _4262_/X _4403_/X _5132_/Y _4829_/A VGND VGND VPWR VPWR _5182_/X sky130_fd_sc_hd__o31a_1
XFILLER_142_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4133_ _6542_/A _4133_/B VGND VGND VPWR VPWR _4138_/S sky130_fd_sc_hd__nand2_4
XFILLER_95_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4064_ _4051_/X hold599/X _4065_/S VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4966_ _4946_/X _4709_/Y _4965_/X _4964_/X VGND VGND VPWR VPWR _4966_/Y sky130_fd_sc_hd__o211ai_1
X_6705_ _7168_/CLK _6705_/D fanout608/X VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfrtp_1
X_3917_ hold13/X _3913_/B _3915_/X _3914_/S hold623/X VGND VGND VPWR VPWR _3917_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4897_ _5140_/C _4589_/B _4589_/C _4746_/X VGND VGND VPWR VPWR _4897_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6636_ _7117_/CLK _6636_/D fanout608/X VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfrtp_4
X_3848_ _6981_/Q _5494_/C _5281_/A2 _3499_/X _7021_/Q VGND VGND VPWR VPWR _3848_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3779_ _6601_/Q _3927_/B _5557_/B _7059_/Q _3778_/X VGND VGND VPWR VPWR _3779_/X
+ sky130_fd_sc_hd__a221o_1
X_6567_ _6676_/CLK _6567_/D fanout577/X VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5518_ _6505_/A1 hold812/X _5520_/S VGND VGND VPWR VPWR _5518_/X sky130_fd_sc_hd__mux2_1
X_6498_ _7257_/Q _6498_/A2 _6498_/B1 _4164_/Y _6497_/X VGND VGND VPWR VPWR _6498_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5449_ hold66/A _5449_/B _5494_/C _5575_/D VGND VGND VPWR VPWR _5457_/S sky130_fd_sc_hd__and4_4
XFILLER_154_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7119_ _7119_/CLK _7119_/D fanout593/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3347_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4820_ _4403_/X _4262_/X _4349_/X _4815_/Y _4358_/X VGND VGND VPWR VPWR _4820_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4751_/A _4945_/B VGND VGND VPWR VPWR _4752_/D sky130_fd_sc_hd__nand2_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3702_ _6686_/Q _6548_/C _5630_/C _5331_/C _3701_/X VGND VGND VPWR VPWR _3702_/X
+ sky130_fd_sc_hd__a41o_1
X_4682_ _4853_/C _4682_/B VGND VGND VPWR VPWR _4685_/B sky130_fd_sc_hd__nand2_1
X_6421_ _6623_/Q _6136_/X _6452_/B1 _6756_/Q _6420_/X VGND VGND VPWR VPWR _6431_/A
+ sky130_fd_sc_hd__a221o_1
X_3633_ _3632_/Y _3633_/A1 _3906_/S VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3564_ _6536_/A _6536_/C _6536_/D VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__and3_2
X_6352_ _6773_/Q _6347_/C _6425_/C _6117_/X _6592_/Q VGND VGND VPWR VPWR _6352_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5303_ _4053_/B _5303_/A1 hold73/X VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
X_6283_ _7164_/Q _6104_/X _6129_/D _6908_/Q _6282_/X VGND VGND VPWR VPWR _6283_/X
+ sky130_fd_sc_hd__a221o_1
X_3495_ _6620_/Q _3954_/B _3492_/X _6663_/Q _3494_/X VGND VGND VPWR VPWR _3507_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5234_ _5234_/A _5234_/B _5234_/C _5234_/D VGND VGND VPWR VPWR _5235_/B sky130_fd_sc_hd__and4_1
XFILLER_69_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5165_ _5165_/A _5165_/B _5165_/C VGND VGND VPWR VPWR _5165_/X sky130_fd_sc_hd__and3_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4116_ _4120_/S _4116_/A2 _3370_/X _5273_/D VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5096_ _5265_/A _5265_/B _5096_/C _5265_/C VGND VGND VPWR VPWR _5098_/A sky130_fd_sc_hd__nand4_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4047_ hold494/X _3921_/B _4054_/S VGND VGND VPWR VPWR _4047_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6773_/Q _5779_/X _5993_/X _5995_/X _5997_/X VGND VGND VPWR VPWR _5998_/X
+ sky130_fd_sc_hd__a2111o_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4949_ _4948_/X _4947_/X _4742_/C _4760_/B VGND VGND VPWR VPWR _4954_/A sky130_fd_sc_hd__o211a_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6619_ _7251_/CLK _6619_/D VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput280 _6831_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
XFILLER_160_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput291 _6737_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_181_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire352 _6365_/Y VGND VGND VPWR VPWR wire352/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire363 _3825_/Y VGND VGND VPWR VPWR _3844_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _6914_/Q VGND VGND VPWR VPWR _3280_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6970_ _7152_/CLK _6970_/D fanout587/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5921_ _7068_/Q _5965_/B _5723_/X _5911_/X _5920_/X VGND VGND VPWR VPWR _5921_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_81_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5852_ _6889_/Q _5795_/C _5815_/C _6028_/B _6913_/Q VGND VGND VPWR VPWR _5852_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4803_ _4735_/Y _4802_/X _4801_/Y _4800_/X VGND VGND VPWR VPWR _4803_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5783_ _6059_/S _5815_/B _5783_/C VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__and3_4
XFILLER_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4734_ _4940_/A _4734_/B _5128_/C VGND VGND VPWR VPWR _4734_/X sky130_fd_sc_hd__and3_1
XFILLER_159_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _4496_/Y _4663_/Y _4664_/Y VGND VGND VPWR VPWR _4665_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6404_ _6765_/Q _6126_/X _6136_/X _6622_/Q _6403_/X VGND VGND VPWR VPWR _6405_/D
+ sky130_fd_sc_hd__a221o_1
Xhold900 _4157_/X VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3616_ _7104_/Q _6548_/A _5281_/A2 _5350_/B _6872_/Q VGND VGND VPWR VPWR _3616_/X
+ sky130_fd_sc_hd__a32o_1
Xhold911 _7022_/Q VGND VGND VPWR VPWR hold911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 _5361_/X VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4596_ _4596_/A _4596_/B _4596_/C VGND VGND VPWR VPWR _4604_/A sky130_fd_sc_hd__nor3_1
XFILLER_134_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold933 _5318_/X VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 _4134_/X VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ _7142_/Q _6177_/C _6114_/X _6116_/X _7134_/Q VGND VGND VPWR VPWR _6335_/X
+ sky130_fd_sc_hd__a32o_1
Xhold955 _6648_/Q VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__dlygate4sd3_1
X_3547_ _5512_/B _6548_/D _5675_/D VGND VGND VPWR VPWR _3547_/X sky130_fd_sc_hd__and3_4
Xhold966 hold966/A VGND VGND VPWR VPWR hold966/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold977 _4022_/X VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 _6778_/Q VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__dlygate4sd3_1
X_3478_ _6967_/Q _5458_/B _5350_/B _6871_/Q _3475_/X VGND VGND VPWR VPWR _3485_/C
+ sky130_fd_sc_hd__a221o_1
Xhold999 _3984_/X VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _6875_/Q _6466_/A1 _5759_/A VGND VGND VPWR VPWR _6266_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5217_ _5102_/Y _5180_/A _5217_/C _5217_/D VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__and4bb_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6197_ _7033_/Q _6138_/B _6108_/X _6109_/X _7041_/Q VGND VGND VPWR VPWR _6197_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5148_ _5147_/X _5235_/C _5148_/C VGND VGND VPWR VPWR _5148_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_84_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5079_ _5079_/A _5079_/B _5079_/C VGND VGND VPWR VPWR _5082_/B sky130_fd_sc_hd__and3_1
XFILLER_56_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ _4450_/A _4450_/B _4450_/C _4450_/D VGND VGND VPWR VPWR _4451_/B sky130_fd_sc_hd__nand4_1
XFILLER_171_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold207 _6641_/Q VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold218 _6966_/Q VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold229 _5339_/X VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ hold24/X hold239/X _3402_/S VGND VGND VPWR VPWR _3401_/X sky130_fd_sc_hd__mux2_1
X_4381_ _4761_/C _4209_/Y _4320_/A _4249_/Y _4870_/B VGND VGND VPWR VPWR _4460_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_98_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3332_ _6858_/Q input78/X _3350_/A VGND VGND VPWR VPWR _3332_/X sky130_fd_sc_hd__mux2_4
X_6120_ _6130_/A _6444_/C _6143_/C VGND VGND VPWR VPWR _6120_/X sky130_fd_sc_hd__and3_2
XFILLER_171_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _7278_/Q _6086_/B1 _5813_/X _6567_/Q _6050_/X VGND VGND VPWR VPWR _6051_/X
+ sky130_fd_sc_hd__a221o_1
X_3263_ _7050_/Q VGND VGND VPWR VPWR _3263_/Y sky130_fd_sc_hd__inv_2
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A _5002_/B VGND VGND VPWR VPWR _5228_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6953_ _7067_/CLK _6953_/D fanout582/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5904_ _6947_/Q _5779_/X _5782_/X _6939_/Q _5903_/X VGND VGND VPWR VPWR _5904_/X
+ sky130_fd_sc_hd__a221o_1
X_6884_ _7168_/CLK _6884_/D fanout608/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _6944_/Q _5779_/X _5782_/X _6936_/Q _5834_/X VGND VGND VPWR VPWR _5835_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5766_ _7183_/Q _7182_/Q _5815_/C VGND VGND VPWR VPWR _5842_/C sky130_fd_sc_hd__and3_4
XFILLER_147_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4717_ _4717_/A _4717_/B _4717_/C VGND VGND VPWR VPWR _4720_/A sky130_fd_sc_hd__nor3_1
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5697_ _6803_/Q _6442_/S _5759_/B _3307_/Y VGND VGND VPWR VPWR _5697_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_108_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4648_ _4777_/B _4674_/D VGND VGND VPWR VPWR _4648_/Y sky130_fd_sc_hd__nand2_2
XFILLER_162_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold730 _6520_/X VGND VGND VPWR VPWR _7240_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _7005_/Q VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4579_ _4579_/A _4579_/B _4579_/C VGND VGND VPWR VPWR _4582_/C sky130_fd_sc_hd__nand3_1
Xhold752 _6573_/Q VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _6570_/Q VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _3996_/X VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _6317_/X _6318_/A1 _6343_/S VGND VGND VPWR VPWR _7213_/D sky130_fd_sc_hd__mux2_1
Xhold785 _3989_/X VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 _6604_/Q VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7298_ _7298_/A VGND VGND VPWR VPWR _7298_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6249_ _7083_/Q _6177_/A _6102_/X _6323_/B1 _6963_/Q VGND VGND VPWR VPWR _6249_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1430 _6968_/Q VGND VGND VPWR VPWR hold343/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _3355_/X VGND VGND VPWR VPWR hold1441/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1452 _7032_/Q VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1463 _6626_/Q VGND VGND VPWR VPWR _3962_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1474 _7215_/Q VGND VGND VPWR VPWR _6392_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7157_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1485 _6802_/Q VGND VGND VPWR VPWR _5752_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1496 _5840_/X VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6889_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_csclk _7277_/CLK VGND VGND VPWR VPWR _7278_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_29_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7017_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3950_ _6477_/A0 _3950_/A1 _3953_/S VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3881_ _6740_/Q _3441_/X _3489_/X _6918_/Q _3880_/X VGND VGND VPWR VPWR _3889_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_189_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5620_ _5620_/A _5630_/A _6548_/B _5675_/D VGND VGND VPWR VPWR _5628_/S sky130_fd_sc_hd__nand4_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ hold2/X hold166/X _5556_/S VGND VGND VPWR VPWR _5551_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4502_ _4319_/X _4423_/Y _4490_/Y _4497_/Y _4501_/Y VGND VGND VPWR VPWR _4504_/C
+ sky130_fd_sc_hd__o32a_1
X_5482_ hold83/X _5482_/A1 _5484_/S VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__mux2_1
XFILLER_184_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7221_ _7251_/CLK _7221_/D VGND VGND VPWR VPWR _7221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4433_ _4427_/C _4429_/D _4383_/A _4391_/Y _4395_/Y VGND VGND VPWR VPWR _4442_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_144_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7152_ _7152_/CLK _7152_/D fanout587/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_98_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4364_ _4698_/A _4657_/C _4722_/A _4984_/A VGND VGND VPWR VPWR _4409_/C sky130_fd_sc_hd__nand4_4
Xfanout506 hold7/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__buf_4
Xfanout517 hold5/X VGND VGND VPWR VPWR _3924_/B sky130_fd_sc_hd__clkbuf_16
X_6103_ _7187_/Q _6138_/B _6425_/B _7188_/Q VGND VGND VPWR VPWR _6103_/X sky130_fd_sc_hd__and4b_4
X_3315_ _4228_/C _4228_/D _4227_/A _4227_/B VGND VGND VPWR VPWR _3317_/B sky130_fd_sc_hd__nor4_1
Xfanout528 hold89/X VGND VGND VPWR VPWR _6538_/A0 sky130_fd_sc_hd__buf_8
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7083_ _7123_/CLK _7083_/D fanout610/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout539 _7184_/Q VGND VGND VPWR VPWR _6059_/S sky130_fd_sc_hd__buf_8
XFILLER_112_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4295_ _4295_/A _4356_/A VGND VGND VPWR VPWR _5055_/D sky130_fd_sc_hd__and2_4
XFILLER_113_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3246_ _6442_/S VGND VGND VPWR VPWR _3246_/Y sky130_fd_sc_hd__clkinv_4
X_6034_ _6645_/Q _6059_/S _5815_/B _5783_/C _6033_/X VGND VGND VPWR VPWR _6034_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _6967_/CLK _6936_/D fanout586/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfstp_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6867_ _7143_/CLK hold70/X fanout587/X VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__dfrtp_1
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5818_ _7000_/Q _5934_/C _5782_/C _5795_/C VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__o211a_1
X_6798_ _7163_/CLK _6798_/D fanout610/X VGND VGND VPWR VPWR _7297_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_10_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5749_ _6143_/D _6141_/B _6425_/B VGND VGND VPWR VPWR _5750_/C sky130_fd_sc_hd__and3_4
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold560 _5579_/X VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold571 _6705_/Q VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 hold582/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
Xhold593 hold593/A VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1260 _3963_/A1 VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _3968_/A1 VGND VGND VPWR VPWR hold686/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _7117_/Q VGND VGND VPWR VPWR _5627_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1293 _6565_/Q VGND VGND VPWR VPWR _3381_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_411 _6451_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_422 _4139_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_433 _6425_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4080_ hold346/X _3915_/X _4092_/S VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4982_ _4984_/A _4984_/B _4984_/C _4982_/D VGND VGND VPWR VPWR _4983_/C sky130_fd_sc_hd__nand4_1
X_6721_ _7143_/CLK _6721_/D fanout587/X VGND VGND VPWR VPWR _7284_/A sky130_fd_sc_hd__dfrtp_1
X_3933_ _6524_/B _6548_/C _5666_/C _5575_/C VGND VGND VPWR VPWR _3934_/S sky130_fd_sc_hd__nand4_4
XFILLER_149_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6652_ _7245_/CLK _6652_/D fanout596/X VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3864_ hold79/A _3496_/X _3861_/X _3863_/X VGND VGND VPWR VPWR _3874_/C sky130_fd_sc_hd__a211o_2
X_5603_ _6549_/A0 _5603_/A1 _5610_/S VGND VGND VPWR VPWR _5603_/X sky130_fd_sc_hd__mux2_1
X_6583_ _7237_/CLK _6583_/D VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3795_ _6782_/Q _5311_/B _5422_/D _3471_/X input24/X VGND VGND VPWR VPWR _3795_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5534_ hold373/X _3921_/B _5538_/S VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5465_ _4051_/B hold480/X _5466_/S VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7204_ _7218_/CLK _7204_/D fanout577/X VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
X_4416_ _4416_/A _4416_/B VGND VGND VPWR VPWR _4416_/Y sky130_fd_sc_hd__nand2_1
X_5396_ _5396_/A0 _5649_/A0 _5403_/S VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7135_ _7135_/CLK _7135_/D fanout588/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4347_ _4243_/A _4243_/B _4346_/Y VGND VGND VPWR VPWR _5044_/A sky130_fd_sc_hd__a21oi_4
XFILLER_160_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7066_ _7122_/CLK _7066_/D fanout607/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_4
X_4278_ _4698_/A _4657_/C _4656_/C _4647_/C VGND VGND VPWR VPWR _4282_/C sky130_fd_sc_hd__and4_1
X_6017_ _7266_/Q _6025_/B wire398/X _5795_/X _6674_/Q VGND VGND VPWR VPWR _6017_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3250__1/A sky130_fd_sc_hd__clkbuf_16
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6919_ _7071_/CLK _6919_/D fanout585/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_168_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold390 _3942_/X VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1090 _5635_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _3916_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_241 hold2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_252 hold211/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 _3446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _3547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _5764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 _5783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3580_ input72/X _5684_/B _5629_/C _4204_/S input44/X VGND VGND VPWR VPWR _3580_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5250_ _4718_/D _4945_/C _4903_/B _4763_/Y VGND VGND VPWR VPWR _5250_/X sky130_fd_sc_hd__a31o_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4201_ _4201_/A0 _4200_/X _4205_/S VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5181_ _4262_/X _4382_/Y _5132_/Y _5055_/Y _4816_/X VGND VGND VPWR VPWR _5238_/C
+ sky130_fd_sc_hd__o311ai_2
XFILLER_96_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4132_ _6535_/A0 hold934/X _4132_/S VGND VGND VPWR VPWR _4132_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4063_ _4049_/X hold645/X _4065_/S VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4965_ _4271_/Y _4344_/Y _5248_/A3 _4707_/Y _4745_/Y VGND VGND VPWR VPWR _4965_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6704_ _7168_/CLK _6704_/D fanout609/X VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_1
X_3916_ _5494_/A hold64/X _3916_/C VGND VGND VPWR VPWR _3916_/X sky130_fd_sc_hd__and3_4
X_4896_ _4894_/X _4732_/X _4893_/X _5200_/B VGND VGND VPWR VPWR _4896_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6635_ _7167_/CLK _6635_/D fanout604/X VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ _6901_/Q _5377_/C _3550_/X _7157_/Q _3846_/X VGND VGND VPWR VPWR _3856_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ _6781_/CLK _6566_/D _3291_/A VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3778_ _6568_/Q _5311_/B _6530_/C _5566_/B _7067_/Q VGND VGND VPWR VPWR _3778_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5517_ _3924_/B hold244/X _5520_/S VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6497_ _7259_/Q _6497_/A2 _6497_/B1 _7258_/Q VGND VGND VPWR VPWR _6497_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5448_ _5448_/A0 _5692_/A1 _5448_/S VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5379_ hold492/X _3916_/C _5385_/S VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7118_ _7162_/CLK _7118_/D fanout605/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7049_ _7065_/CLK _7049_/D fanout599/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _5263_/B _4750_/B VGND VGND VPWR VPWR _4752_/C sky130_fd_sc_hd__nand2_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3701_ _6746_/Q _3368_/X _5485_/B _3438_/X _7002_/Q VGND VGND VPWR VPWR _3701_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4681_ _4681_/A _4681_/B _4681_/C _4681_/D VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__nand4_1
XFILLER_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6420_ _6666_/Q _6451_/B1 _6130_/X _6781_/Q _6419_/X VGND VGND VPWR VPWR _6420_/X
+ sky130_fd_sc_hd__a221o_1
X_3632_ _3582_/X _3632_/B _3632_/C VGND VGND VPWR VPWR _3632_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6351_ _6811_/Q _6107_/X _6347_/X _6348_/X _6350_/X VGND VGND VPWR VPWR _6356_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3563_ _3563_/A _6548_/D hold28/A VGND VGND VPWR VPWR _3563_/X sky130_fd_sc_hd__and3_1
XFILLER_115_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5302_ hold21/X hold115/X hold73/X VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6282_ _7172_/Q _6130_/A _6114_/X _6281_/X VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__a31o_1
X_3494_ _6851_/Q _5666_/C _5325_/C _3493_/X VGND VGND VPWR VPWR _3494_/X sky130_fd_sc_hd__a31o_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5233_ _4970_/B _4730_/D _5190_/X VGND VGND VPWR VPWR _5234_/D sky130_fd_sc_hd__a21oi_1
XFILLER_102_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5164_ _5164_/A _5249_/A _5247_/A VGND VGND VPWR VPWR _5165_/A sky130_fd_sc_hd__and3_1
X_4115_ _5476_/B _6524_/B _6536_/C _5273_/D VGND VGND VPWR VPWR _4120_/S sky130_fd_sc_hd__nand4_4
XFILLER_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5095_ _4640_/A _5090_/X _4570_/A VGND VGND VPWR VPWR _5265_/C sky130_fd_sc_hd__a21oi_1
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4046_ hold301/X _3918_/B _4054_/S VGND VGND VPWR VPWR _4046_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _7275_/Q _6086_/B1 _5771_/X _6758_/Q _5996_/X VGND VGND VPWR VPWR _5997_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4948_ _4751_/A _4730_/A _4699_/B _4923_/B _4755_/B VGND VGND VPWR VPWR _4948_/X
+ sky130_fd_sc_hd__a32o_1
X_4879_ _4879_/A _4879_/B _4879_/C _4879_/D VGND VGND VPWR VPWR _4881_/A sky130_fd_sc_hd__nor4_1
X_6618_ _7251_/CLK _6618_/D VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6549_ _6549_/A0 _6549_/A1 _6553_/S VGND VGND VPWR VPWR _6549_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput270 _6825_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
XFILLER_133_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput281 _6832_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
Xoutput292 hold93/A VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_87_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire353 _6339_/Y VGND VGND VPWR VPWR _6340_/C sky130_fd_sc_hd__clkbuf_1
Xwire364 _3592_/Y VGND VGND VPWR VPWR _3632_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ _7052_/Q _5814_/X _5815_/X _7020_/Q _5919_/X VGND VGND VPWR VPWR _5920_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5851_ _7065_/Q _5723_/X wire398/X _7089_/Q _5850_/X VGND VGND VPWR VPWR _5851_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _4632_/A _5036_/B _4753_/B _4496_/Y VGND VGND VPWR VPWR _4802_/X sky130_fd_sc_hd__o31a_1
XFILLER_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5782_ _6010_/D _5795_/D _5782_/C VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__and3_4
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4733_ _4675_/A _5128_/A _4732_/C _4732_/X _4729_/A VGND VGND VPWR VPWR _4737_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_175_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4664_ _4557_/A _4761_/C _4792_/B _4750_/B VGND VGND VPWR VPWR _4664_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6403_ _7262_/Q _6446_/C _6425_/C _6138_/X _6609_/Q VGND VGND VPWR VPWR _6403_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3615_ _7096_/Q _3510_/X _3570_/X _3573_/X _3614_/X VGND VGND VPWR VPWR _3615_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_134_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4595_ _4595_/A _5140_/C _4923_/A VGND VGND VPWR VPWR _4596_/B sky130_fd_sc_hd__and3_1
Xhold901 _7054_/Q VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 _5520_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold923 _7153_/Q VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold934 _6757_/Q VGND VGND VPWR VPWR hold934/X sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ _6958_/Q _6142_/X _6177_/X _7022_/Q _6333_/X VGND VGND VPWR VPWR _6339_/B
+ sky130_fd_sc_hd__a221o_1
Xhold945 hold945/A VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__dlygate4sd3_1
X_3546_ _6927_/Q _5413_/B _3543_/X _3545_/X _3541_/X VGND VGND VPWR VPWR _3561_/B
+ sky130_fd_sc_hd__a2111o_4
Xhold956 _3988_/X VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _6675_/Q VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold978 hold978/A VGND VGND VPWR VPWR hold978/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold989 _4159_/X VGND VGND VPWR VPWR _6778_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _6246_/X _6265_/B _6265_/C VGND VGND VPWR VPWR _6265_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3477_ _5630_/C _5675_/D _5331_/C VGND VGND VPWR VPWR _5350_/B sky130_fd_sc_hd__and3_4
X_5216_ _5216_/A _5216_/B _5216_/C _5216_/D VGND VGND VPWR VPWR _5217_/D sky130_fd_sc_hd__nor4_1
X_6196_ _7089_/Q _6106_/X _6110_/X _7113_/Q _6195_/X VGND VGND VPWR VPWR _6196_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5147_ _5060_/A _4505_/B _4815_/A _4488_/X _4843_/B VGND VGND VPWR VPWR _5147_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5078_ _4946_/X _4633_/Y _4613_/Y _5248_/A3 _4707_/Y VGND VGND VPWR VPWR _5079_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4029_ _6542_/A _4029_/B VGND VGND VPWR VPWR _4034_/S sky130_fd_sc_hd__nand2_4
XFILLER_72_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold208 _3979_/X VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 _5457_/X VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3400_ _3918_/B hold609/X _3402_/S VGND VGND VPWR VPWR _3400_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4380_ _4243_/A _4243_/B _4262_/X _4346_/Y VGND VGND VPWR VPWR _4380_/X sky130_fd_sc_hd__a211o_2
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3331_ _6857_/Q input80/X _3350_/A VGND VGND VPWR VPWR _3331_/X sky130_fd_sc_hd__mux2_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6746_/Q _6028_/C _6025_/C _5774_/X _6671_/Q VGND VGND VPWR VPWR _6050_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _7058_/Q VGND VGND VPWR VPWR _3262_/Y sky130_fd_sc_hd__inv_2
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _4984_/A _4704_/B _5255_/A _4719_/B _4792_/C VGND VGND VPWR VPWR _5002_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6952_ _7087_/CLK _6952_/D fanout584/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5903_ _7091_/Q _6072_/B wire398/X _5795_/X _6899_/Q VGND VGND VPWR VPWR _5903_/X
+ sky130_fd_sc_hd__a32o_1
X_6883_ _6957_/CLK _6883_/D fanout591/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5834_ _7088_/Q _6072_/B wire398/X _5795_/X _6896_/Q VGND VGND VPWR VPWR _5834_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_179_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5765_ _7180_/Q _7181_/Q VGND VGND VPWR VPWR _5815_/C sky130_fd_sc_hd__and2b_4
X_4716_ _4716_/A _4862_/A _4729_/D VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__and3_1
X_5696_ _6803_/Q _6442_/S _5759_/B _3307_/Y VGND VGND VPWR VPWR _5706_/D sky130_fd_sc_hd__o31a_1
XFILLER_147_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4647_ _4698_/A _4656_/C _4647_/C _4657_/C VGND VGND VPWR VPWR _4755_/B sky130_fd_sc_hd__and4bb_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold720 _7069_/Q VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _6575_/Q VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ _4751_/A _4597_/B _4923_/A _4589_/C VGND VGND VPWR VPWR _4579_/C sky130_fd_sc_hd__nand4_1
Xhold742 _5501_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold753 _3393_/X VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6317_ _6292_/S _7212_/Q _6315_/Y _6316_/X VGND VGND VPWR VPWR _6317_/X sky130_fd_sc_hd__a22o_1
Xhold764 _3390_/X VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ _6773_/Q _4152_/C _3528_/X input11/X _3526_/X VGND VGND VPWR VPWR _3529_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold775 _6676_/Q VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlygate4sd3_1
X_7297_ _7297_/A VGND VGND VPWR VPWR _7297_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold786 hold786/A VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _3936_/X VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6248_ _6899_/Q _6129_/A _6107_/X hold91/A _6247_/X VGND VGND VPWR VPWR _6255_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6179_ _7064_/Q _6103_/X _6144_/X _7080_/Q _6178_/X VGND VGND VPWR VPWR _6179_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1420 _3401_/X VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 _5460_/X VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 _4108_/S VGND VGND VPWR VPWR _4111_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _5532_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 _6740_/Q VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1475 _6368_/X VGND VGND VPWR VPWR _7215_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1486 _7193_/Q VGND VGND VPWR VPWR _5758_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _7208_/Q VGND VGND VPWR VPWR _6217_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3880_ _6982_/Q _5273_/D _5281_/A2 _3471_/X input28/X VGND VGND VPWR VPWR _3880_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_71_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5550_ _6550_/A0 hold779/X _5550_/S VGND VGND VPWR VPWR _5550_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4501_ _4729_/A _4792_/B VGND VGND VPWR VPWR _4501_/Y sky130_fd_sc_hd__nand2_2
X_5481_ _3925_/C hold409/X _5484_/S VGND VGND VPWR VPWR _5481_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7220_ _7256_/CLK _7220_/D _6472_/A VGND VGND VPWR VPWR _7220_/Q sky130_fd_sc_hd__dfrtp_4
X_4432_ _4427_/C _4429_/D _4383_/A _4388_/Y _4395_/Y VGND VGND VPWR VPWR _4442_/C
+ sky130_fd_sc_hd__a2111o_1
X_7151_ _7151_/CLK _7151_/D fanout586/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfstp_1
X_4363_ _4363_/A _4722_/A _4984_/A VGND VGND VPWR VPWR _4721_/C sky130_fd_sc_hd__and3_1
XFILLER_113_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout507 _6511_/A1 VGND VGND VPWR VPWR _5692_/A1 sky130_fd_sc_hd__buf_6
X_6102_ _6141_/B _7190_/Q _7189_/Q _6143_/D VGND VGND VPWR VPWR _6102_/X sky130_fd_sc_hd__and4bb_4
X_3314_ _4229_/C _4229_/D _4228_/A _4228_/B VGND VGND VPWR VPWR _3318_/C sky130_fd_sc_hd__nor4_1
Xfanout518 hold47/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__buf_12
Xfanout529 hold89/X VGND VGND VPWR VPWR _3916_/C sky130_fd_sc_hd__buf_8
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7082_ _7170_/CLK hold45/X fanout605/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4294_ _4939_/A _4294_/B _4804_/A VGND VGND VPWR VPWR _4843_/A sky130_fd_sc_hd__and3_1
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6033_ _6650_/Q _6059_/S _6009_/C _5788_/X _6745_/Q VGND VGND VPWR VPWR _6033_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7071_/CLK _6935_/D fanout585/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6866_ _7077_/CLK _6866_/D fanout587/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5817_ _5817_/A1 _6443_/S _5816_/X VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__a21o_1
X_6797_ _7163_/CLK _6797_/D fanout608/X VGND VGND VPWR VPWR _7296_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ _7190_/Q _7189_/Q VGND VGND VPWR VPWR _6134_/C sky130_fd_sc_hd__nand2b_2
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5679_ hold8/X _3509_/X _3921_/X _5683_/S hold631/X VGND VGND VPWR VPWR _5679_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_175_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold550 _6978_/Q VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _6704_/Q VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold572 _4062_/X VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _6848_/Q VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold594 hold594/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1250 _3694_/A1 VGND VGND VPWR VPWR hold519/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 _3953_/A1 VGND VGND VPWR VPWR hold601/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 _6480_/A1 VGND VGND VPWR VPWR hold694/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _6555_/Q VGND VGND VPWR VPWR _3363_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1294 _7091_/Q VGND VGND VPWR VPWR _5598_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_401 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_412 _6072_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_423 _5723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_434 _6425_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput170 wb_we_i VGND VGND VPWR VPWR _6514_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4981_ _4290_/Y _4423_/Y _4501_/Y _4740_/Y _5200_/B VGND VGND VPWR VPWR _4981_/X
+ sky130_fd_sc_hd__o311a_1
X_6720_ _7077_/CLK _6720_/D fanout587/X VGND VGND VPWR VPWR _7283_/A sky130_fd_sc_hd__dfrtp_1
X_3932_ _6535_/A0 _3932_/A1 _3932_/S VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6651_ _7275_/CLK _6651_/D fanout596/X VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfrtp_4
X_3863_ input59/X _3539_/X _5413_/B _6933_/Q _3862_/X VGND VGND VPWR VPWR _3863_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5602_ _5630_/A _6548_/B _6548_/D _5675_/D VGND VGND VPWR VPWR _5610_/S sky130_fd_sc_hd__nand4_4
X_6582_ _7218_/CLK _6582_/D VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfxtp_1
X_3794_ _6939_/Q hold39/A _3542_/B _3539_/X input56/X VGND VGND VPWR VPWR _3794_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5533_ hold222/X hold2/X _5538_/S VGND VGND VPWR VPWR _5533_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5464_ hold83/X hold164/X _5466_/S VGND VGND VPWR VPWR _5464_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7154_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7203_ _7218_/CLK _7203_/D fanout594/X VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4415_ _4427_/C _4429_/D _4383_/A _4398_/X VGND VGND VPWR VPWR _4415_/X sky130_fd_sc_hd__a211o_1
XFILLER_132_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5395_ _5476_/B _6524_/B _5422_/D _5575_/D VGND VGND VPWR VPWR _5403_/S sky130_fd_sc_hd__and4_4
X_7134_ _7173_/CLK _7134_/D fanout603/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfrtp_1
X_4346_ _4346_/A _4670_/D VGND VGND VPWR VPWR _4346_/Y sky130_fd_sc_hd__nand2_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7087_/CLK sky130_fd_sc_hd__clkbuf_16
X_7065_ _7065_/CLK _7065_/D fanout590/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4277_ _4632_/A _4632_/B _4600_/B _4612_/C VGND VGND VPWR VPWR _4277_/Y sky130_fd_sc_hd__nand4_4
X_6016_ _7271_/Q _5780_/X _6013_/X _6015_/X VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__a211o_1
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _7154_/CLK _6918_/D fanout592/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7279_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6849_ _6889_/CLK _6849_/D fanout584/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7167_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_182_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold380 hold380/A VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 hold391/A VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1080 _5342_/X VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1091 _7047_/Q VGND VGND VPWR VPWR _5549_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_220 _3925_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _6550_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 hold5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 hold211/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _5639_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_275 _3678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _5842_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_297 _5783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4200_ hold645/X _4049_/X _4204_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
X_5180_ _5180_/A _5180_/B VGND VGND VPWR VPWR _5180_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4131_ _6546_/A0 hold508/X _4132_/S VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4062_ _3924_/X hold571/X _4065_/S VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4964_ _5248_/A3 _4946_/X _4699_/Y _4963_/X _4962_/X VGND VGND VPWR VPWR _4964_/X
+ sky130_fd_sc_hd__o311a_1
X_6703_ _7168_/CLK _6703_/D fanout609/X VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3915_ hold65/X _3915_/B VGND VGND VPWR VPWR _3915_/X sky130_fd_sc_hd__and2_4
X_4895_ _5128_/A _5128_/C _5263_/B _4623_/Y VGND VGND VPWR VPWR _5200_/B sky130_fd_sc_hd__a31oi_2
XFILLER_60_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6634_ _6843_/CLK _6634_/D fanout584/X VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_4
X_3846_ _6957_/Q _3424_/X _3521_/X _7173_/Q _3573_/X VGND VGND VPWR VPWR _3846_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6565_ _7260_/CLK hold90/X fanout579/X VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3777_ _7279_/Q _6548_/A _3466_/X _5639_/B _7131_/Q VGND VGND VPWR VPWR _3777_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5516_ hold13/X _3499_/X _3921_/X _5520_/S hold490/X VGND VGND VPWR VPWR _5516_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_180_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6496_ _6495_/X _3918_/B _6511_/S VGND VGND VPWR VPWR _7231_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5447_ hold690/X _4051_/B _5448_/S VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5378_ hold724/X _5667_/A0 _5385_/S VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7117_ _7117_/CLK hold22/X fanout608/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_2
X_4329_ _4940_/C _4320_/B _4523_/A VGND VGND VPWR VPWR _4509_/B sky130_fd_sc_hd__o21ai_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7048_ _7129_/CLK _7048_/D fanout598/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3700_ _7082_/Q _5630_/A _5440_/C _5350_/B _6874_/Q VGND VGND VPWR VPWR _3700_/X
+ sky130_fd_sc_hd__a32o_1
X_4680_ _4804_/C _4682_/B VGND VGND VPWR VPWR _4681_/C sky130_fd_sc_hd__nand2_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3631_ _3631_/A _3631_/B _3631_/C _3631_/D VGND VGND VPWR VPWR _3631_/Y sky130_fd_sc_hd__nor4_1
X_6350_ _6763_/Q _6126_/X _6130_/X _6778_/Q _6349_/X VGND VGND VPWR VPWR _6350_/X
+ sky130_fd_sc_hd__a221o_1
X_3562_ _3987_/A _5512_/B _5657_/D VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__and3_4
X_5301_ hold83/X hold96/X hold73/X VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6281_ _7028_/Q _6136_/A _6328_/A3 _6113_/X _7148_/Q VGND VGND VPWR VPWR _6281_/X
+ sky130_fd_sc_hd__a32o_1
X_3493_ _7239_/Q hold17/A _5325_/C VGND VGND VPWR VPWR _3493_/X sky130_fd_sc_hd__and3_1
XFILLER_115_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5232_ _5125_/B _5197_/B _5228_/X _5258_/C _5226_/Y VGND VGND VPWR VPWR _5243_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_130_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5163_ _4788_/A _4950_/X _5162_/X VGND VGND VPWR VPWR _5247_/A sky130_fd_sc_hd__a21oi_1
X_4114_ hold362/X _3916_/C _4114_/S VGND VGND VPWR VPWR _4114_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5094_ _5094_/A _5094_/B _5175_/B VGND VGND VPWR VPWR _5096_/C sky130_fd_sc_hd__nor3b_1
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4045_ hold360/X _3916_/C _4054_/S VGND VGND VPWR VPWR _4045_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _7265_/Q _6025_/B wire398/X _5795_/X _6673_/Q VGND VGND VPWR VPWR _5996_/X
+ sky130_fd_sc_hd__a32o_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4947_ _4804_/C _4923_/B _4750_/B _4761_/C VGND VGND VPWR VPWR _4947_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4878_ _4878_/A _4878_/B _4878_/C VGND VGND VPWR VPWR _4879_/B sky130_fd_sc_hd__and3_1
XFILLER_20_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6617_ _7259_/CLK _6617_/D VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3829_ _7132_/Q _5639_/B _3539_/X input57/X _3828_/X VGND VGND VPWR VPWR _3834_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6548_ _6548_/A _6548_/B _6548_/C _6548_/D VGND VGND VPWR VPWR _6553_/S sky130_fd_sc_hd__nand4_4
XFILLER_192_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6479_ _3875_/Y _6479_/A1 _6480_/S VGND VGND VPWR VPWR _7227_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput260 _6837_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
Xoutput271 _6733_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
Xoutput282 _6734_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
Xoutput293 _6739_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_87_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire354 _6314_/Y VGND VGND VPWR VPWR _6315_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_128_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire365 _6305_/Y VGND VGND VPWR VPWR _6315_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_183_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire398 _5769_/X VGND VGND VPWR VPWR wire398/X sky130_fd_sc_hd__buf_12
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5850_ _7033_/Q _6010_/C _5814_/C _6009_/C _7081_/Q VGND VGND VPWR VPWR _5850_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_34_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _4801_/A _4801_/B _5036_/C _5128_/C VGND VGND VPWR VPWR _4801_/Y sky130_fd_sc_hd__nand4_1
X_5781_ _7180_/Q _5795_/C _7181_/Q VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__and3b_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4732_ _5128_/A _4860_/C _4732_/C VGND VGND VPWR VPWR _4732_/X sky130_fd_sc_hd__and3_1
XFILLER_159_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4663_ _4674_/C _4674_/D VGND VGND VPWR VPWR _4663_/Y sky130_fd_sc_hd__nand2_4
XFILLER_175_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6402_ _6561_/Q _5750_/X _6103_/X _7246_/Q _6401_/X VGND VGND VPWR VPWR _6405_/C
+ sky130_fd_sc_hd__a221o_1
X_3614_ _6759_/Q _4133_/B _3418_/X _6744_/Q _3613_/X VGND VGND VPWR VPWR _3614_/X
+ sky130_fd_sc_hd__a221o_2
X_4594_ _4815_/A _4595_/A _4923_/A VGND VGND VPWR VPWR _4596_/A sky130_fd_sc_hd__and3_1
Xhold902 _5556_/X VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _7086_/Q VGND VGND VPWR VPWR hold913/X sky130_fd_sc_hd__dlygate4sd3_1
X_3545_ _6643_/Q _5485_/B _3457_/X _3544_/X _6943_/Q VGND VGND VPWR VPWR _3545_/X
+ sky130_fd_sc_hd__a32o_1
Xhold924 _5669_/X VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6333_ _7078_/Q _6425_/B _6139_/X _6117_/X _7174_/Q VGND VGND VPWR VPWR _6333_/X
+ sky130_fd_sc_hd__a32o_1
Xhold935 _4132_/X VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _6674_/Q VGND VGND VPWR VPWR hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _6760_/Q VGND VGND VPWR VPWR hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _4020_/X VGND VGND VPWR VPWR _6675_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6264_ _6264_/A _6264_/B _6264_/C _6339_/D VGND VGND VPWR VPWR _6265_/C sky130_fd_sc_hd__nor4_2
X_3476_ _4127_/C _5476_/C _5494_/C VGND VGND VPWR VPWR _5458_/B sky130_fd_sc_hd__and3_4
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5215_ _4620_/A _4595_/A _4620_/C _4615_/X _5214_/X VGND VGND VPWR VPWR _5216_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_130_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6195_ _7145_/Q _6113_/X _6141_/X _6977_/Q _6194_/X VGND VGND VPWR VPWR _6195_/X
+ sky130_fd_sc_hd__a221o_1
X_5146_ _5234_/A _5146_/B _5146_/C _5146_/D VGND VGND VPWR VPWR _5148_/C sky130_fd_sc_hd__and4_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5077_ _4946_/X _4633_/Y _4613_/Y _5248_/A3 _4699_/Y VGND VGND VPWR VPWR _5079_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4028_ hold938/X _6535_/A0 _4028_/S VGND VGND VPWR VPWR _4028_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5979_ _6811_/Q _6028_/C _5782_/C _5795_/C VGND VGND VPWR VPWR _5979_/X sky130_fd_sc_hd__o211a_1
XFILLER_52_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 _6990_/Q VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3330_ _7154_/Q _3350_/A _3329_/Y VGND VGND VPWR VPWR _3330_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _7066_/Q VGND VGND VPWR VPWR _3261_/Y sky130_fd_sc_hd__inv_2
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5000_ _4501_/Y _4638_/Y _4699_/Y _4999_/X _4881_/B VGND VGND VPWR VPWR _5003_/C
+ sky130_fd_sc_hd__o311a_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6951_ _7087_/CLK _6951_/D fanout589/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5902_ _7075_/Q _5971_/A2 _5899_/X _5901_/X VGND VGND VPWR VPWR _5902_/X sky130_fd_sc_hd__a211o_1
X_6882_ _7171_/CLK _6882_/D fanout610/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5833_ _7104_/Q _5764_/X _5784_/X _7024_/Q _5832_/X VGND VGND VPWR VPWR _5833_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5764_ _6059_/S _7183_/Q _7182_/Q _5783_/C VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__and4_4
XFILLER_148_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4715_ _4740_/C _4987_/B VGND VGND VPWR VPWR _4715_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5695_ _3297_/Y _5694_/B _5695_/A3 _5694_/Y VGND VGND VPWR VPWR _7175_/D sky130_fd_sc_hd__a31o_1
XFILLER_148_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4646_ _4718_/D _4682_/B VGND VGND VPWR VPWR _4681_/D sky130_fd_sc_hd__nand2_1
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold710 _6893_/Q VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _5573_/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4577_ _4597_/B _4597_/C _4923_/A _4589_/C VGND VGND VPWR VPWR _4579_/B sky130_fd_sc_hd__nand4_1
Xhold732 _3399_/X VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap451 _3757_/D VGND VGND VPWR VPWR _5313_/D sky130_fd_sc_hd__buf_2
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold743 hold743/A VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 hold754/A VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ _6877_/Q _6134_/Y _3246_/Y VGND VGND VPWR VPWR _6316_/X sky130_fd_sc_hd__o21a_1
X_3528_ _5304_/A _4127_/C _3528_/C VGND VGND VPWR VPWR _3528_/X sky130_fd_sc_hd__and3_4
Xhold765 _6639_/Q VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 _4021_/X VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7296_ _7296_/A VGND VGND VPWR VPWR _7296_/X sky130_fd_sc_hd__clkbuf_2
Xhold787 _6603_/Q VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold798 hold798/A VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3459_ _6536_/C _6536_/D _4158_/D VGND VGND VPWR VPWR _4017_/B sky130_fd_sc_hd__and3_4
X_6247_ _7075_/Q _6425_/B _6139_/X _6119_/X _7051_/Q VGND VGND VPWR VPWR _6247_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1410 _7246_/Q VGND VGND VPWR VPWR hold404/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6178_ _7008_/Q _6117_/C _6096_/Y _6118_/X _7056_/Q VGND VGND VPWR VPWR _6178_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1421 _7241_/Q VGND VGND VPWR VPWR hold1421/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1432 _7103_/Q VGND VGND VPWR VPWR hold1432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 _4109_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5129_ _4675_/A _5128_/A _4732_/C _4732_/X _5128_/X VGND VGND VPWR VPWR _5129_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1454 _6630_/Q VGND VGND VPWR VPWR _3966_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 _6831_/Q VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1476 _6619_/Q VGND VGND VPWR VPWR _3953_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _7217_/Q VGND VGND VPWR VPWR _6442_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _6808_/Q VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4500_ _4789_/B _5036_/B _4689_/B VGND VGND VPWR VPWR _4804_/C sky130_fd_sc_hd__and3_4
X_5480_ _3921_/B hold658/X _5484_/S VGND VGND VPWR VPWR _5480_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4431_ _4427_/C _4429_/D _4383_/A _5040_/B _4395_/Y VGND VGND VPWR VPWR _4442_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7150_ _7150_/CLK _7150_/D fanout603/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfrtp_1
X_4362_ _4761_/C _4320_/A _4280_/A _4683_/B VGND VGND VPWR VPWR _4668_/C sky130_fd_sc_hd__o31ai_4
XFILLER_153_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6101_ _6117_/C _6347_/C _6177_/C VGND VGND VPWR VPWR _6101_/X sky130_fd_sc_hd__and3_4
X_3313_ input123/X input122/X _3313_/C _3313_/D VGND VGND VPWR VPWR _3319_/C sky130_fd_sc_hd__and4bb_1
Xfanout508 _4053_/B VGND VGND VPWR VPWR _6511_/A1 sky130_fd_sc_hd__buf_6
X_7081_ _7167_/CLK _7081_/D fanout604/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout519 _3922_/C VGND VGND VPWR VPWR _6546_/A0 sky130_fd_sc_hd__buf_8
XFILLER_113_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4293_ _4294_/B _4804_/A VGND VGND VPWR VPWR _4293_/Y sky130_fd_sc_hd__nand2_2
XFILLER_86_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6032_ _6765_/Q _5770_/X _5793_/X _6750_/Q _6031_/X VGND VGND VPWR VPWR _6032_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6934_ _7173_/CLK _6934_/D fanout602/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6865_ _7143_/CLK _6865_/D fanout587/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_1
X_5816_ _6871_/Q _5726_/Y _5802_/X _5812_/X _5759_/X VGND VGND VPWR VPWR _5816_/X
+ sky130_fd_sc_hd__o221a_1
X_6796_ _7163_/CLK _6796_/D fanout610/X VGND VGND VPWR VPWR _7295_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5747_ _7190_/Q _7189_/Q VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__and2b_1
X_5678_ _5683_/S hold919/X _3509_/X _3919_/X VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4629_ _4777_/A _4674_/C VGND VGND VPWR VPWR _4629_/Y sky130_fd_sc_hd__nand2_4
XFILLER_190_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 _6766_/Q VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold551 _5471_/X VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold562 _4061_/X VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold573 _6999_/Q VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold584 _5321_/X VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold595/A VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__dlygate4sd3_1
X_7279_ _7279_/CLK _7279_/D fanout597/X VGND VGND VPWR VPWR _7279_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1240 _6823_/Q VGND VGND VPWR VPWR _5289_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1251 _3845_/A1 VGND VGND VPWR VPWR hold534/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1262 _6473_/A1 VGND VGND VPWR VPWR hold597/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 _6478_/A1 VGND VGND VPWR VPWR hold706/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 _6844_/Q VGND VGND VPWR VPWR _5317_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_402 _6115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 _7109_/Q VGND VGND VPWR VPWR _5618_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_413 hold39/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_424 _5776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_435 _6425_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6507_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4980_ _4979_/X _4846_/X _4206_/B _4980_/B2 VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3931_ _6546_/A0 hold591/X _3932_/S VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6650_ _6650_/CLK _6650_/D fanout596/X VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfstp_1
X_3862_ _7149_/Q _5684_/B _5440_/C _5404_/B _6925_/Q VGND VGND VPWR VPWR _3862_/X
+ sky130_fd_sc_hd__a32o_1
X_5601_ _5692_/A1 hold925/X hold14/X VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6581_ _7218_/CLK _6581_/D VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfxtp_1
X_3793_ _7011_/Q _5503_/B _3788_/X _3789_/X _3792_/X VGND VGND VPWR VPWR _3810_/C
+ sky130_fd_sc_hd__a2111o_2
X_5532_ hold163/X hold89/X _5538_/S VGND VGND VPWR VPWR _5532_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_csclk _7277_/CLK VGND VGND VPWR VPWR _7089_/CLK sky130_fd_sc_hd__clkbuf_16
X_5463_ hold5/X hold61/X _5466_/S VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__mux2_1
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7202_ _7218_/CLK _7202_/D fanout577/X VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_1
X_4414_ _4427_/C _4429_/D _4383_/A _4395_/Y VGND VGND VPWR VPWR _4414_/X sky130_fd_sc_hd__a211o_1
X_5394_ _5394_/A0 _5692_/A1 _5394_/S VGND VGND VPWR VPWR _5394_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7133_ _7133_/CLK _7133_/D fanout601/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4345_ _4214_/A _4214_/B _4284_/A VGND VGND VPWR VPWR _5042_/B sky130_fd_sc_hd__a21oi_4
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7064_ _7108_/CLK _7064_/D fanout606/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_113_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4276_ _4632_/A _4511_/A _4632_/C _4729_/A VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__and4_4
XFILLER_86_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6015_ _7261_/Q _5777_/X _5813_/X _6565_/Q _6014_/X VGND VGND VPWR VPWR _6015_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6917_ _7015_/CLK _6917_/D fanout588/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6848_ _6889_/CLK _6848_/D fanout582/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6779_ _6781_/CLK _6779_/D _3291_/A VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 _4048_/X VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold381 _7026_/Q VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _7269_/Q VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1070 _5665_/X VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 _6726_/Q VGND VGND VPWR VPWR _4096_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 _5549_/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _5512_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 _3924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_232 _6550_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_243 hold5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 hold211/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _3466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 _3685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 _5842_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_298 _5795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4130_ _6539_/A0 _4130_/A1 _4132_/S VGND VGND VPWR VPWR _4130_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4061_ _3921_/X hold561/X _4065_/S VGND VGND VPWR VPWR _4061_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4963_ _4699_/Y _4745_/Y _4939_/Y _4707_/Y VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__o22a_1
X_6702_ _7140_/CLK _6702_/D fanout609/X VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfrtp_1
X_3914_ _6549_/A0 _3914_/A1 _3914_/S VGND VGND VPWR VPWR _3914_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4894_ _5128_/A _5128_/C _4718_/D _4738_/X VGND VGND VPWR VPWR _4894_/X sky130_fd_sc_hd__a31o_1
XFILLER_189_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6633_ _6835_/CLK _6633_/D fanout583/X VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfrtp_2
X_3845_ _3844_/Y _3845_/A1 _3906_/S VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6564_ _6751_/CLK _6564_/D _3291_/A VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfrtp_4
X_3776_ _7091_/Q _5593_/B _3768_/X _3770_/X _3775_/X VGND VGND VPWR VPWR _3776_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5515_ hold13/X _3499_/X _3918_/X _5520_/S hold990/X VGND VGND VPWR VPWR _5515_/X
+ sky130_fd_sc_hd__a32o_1
X_6495_ _7258_/Q _6495_/A2 _6495_/B1 _4164_/Y _6494_/X VGND VGND VPWR VPWR _6495_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5446_ _5446_/A0 hold83/X _5448_/S VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__mux2_1
XFILLER_172_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5377_ _5494_/A hold64/X _5377_/C VGND VGND VPWR VPWR _5385_/S sky130_fd_sc_hd__and3_4
XFILLER_87_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7116_ _7122_/CLK _7116_/D fanout607/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_1
X_4328_ _4208_/Y _4940_/C _4761_/C VGND VGND VPWR VPWR _4523_/A sky130_fd_sc_hd__o21ai_4
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7047_ _7117_/CLK _7047_/D fanout608/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfstp_2
X_4259_ _4429_/A _4429_/D VGND VGND VPWR VPWR _4259_/Y sky130_fd_sc_hd__nand2_2
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire558 _4792_/B VGND VGND VPWR VPWR _4712_/B sky130_fd_sc_hd__buf_2
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7135_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3630_ _7271_/Q _6542_/B _3626_/X _3627_/X _3629_/X VGND VGND VPWR VPWR _3631_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_186_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3561_ _3561_/A _3561_/B _3561_/C _3561_/D VGND VGND VPWR VPWR _3568_/C sky130_fd_sc_hd__nor4_4
XFILLER_127_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5300_ hold5/X _5300_/A1 hold73/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_89_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7244_/CLK sky130_fd_sc_hd__clkbuf_16
X_3492_ _6536_/C _4127_/C _3533_/C VGND VGND VPWR VPWR _3492_/X sky130_fd_sc_hd__and3_2
X_6280_ _6924_/Q _6129_/B _6454_/B1 _6956_/Q _6279_/X VGND VGND VPWR VPWR _6280_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5231_ _5231_/A _5231_/B _5231_/C _5231_/D VGND VGND VPWR VPWR _5258_/C sky130_fd_sc_hd__and4_1
XFILLER_102_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5162_ _4945_/B _4804_/C _4789_/D _4788_/X _5161_/X VGND VGND VPWR VPWR _5162_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_csclk _7277_/CLK VGND VGND VPWR VPWR _6650_/CLK sky130_fd_sc_hd__clkbuf_16
X_4113_ _4113_/A0 _5649_/A0 _4114_/S VGND VGND VPWR VPWR _4113_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5093_ _4522_/Y _4613_/Y _4648_/Y _4560_/C _4909_/C VGND VGND VPWR VPWR _5175_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4044_ _5667_/A0 _4187_/S _5341_/C hold654/X VGND VGND VPWR VPWR _4044_/X sky130_fd_sc_hd__a31o_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7114_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5995_ _6653_/Q _6028_/C _5723_/X _5994_/X VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__a31o_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4946_ _4689_/B _4255_/A _4753_/A _4501_/Y VGND VGND VPWR VPWR _4946_/X sky130_fd_sc_hd__o31a_4
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4877_ _4689_/A _4860_/B _4860_/C _4708_/A _4778_/C VGND VGND VPWR VPWR _4879_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_178_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6616_ _7237_/CLK _6616_/D VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_138_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3828_ input49/X _5311_/B hold56/A _5359_/B _6884_/Q VGND VGND VPWR VPWR _3828_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6547_ _3925_/C hold383/X _6547_/S VGND VGND VPWR VPWR _6547_/X sky130_fd_sc_hd__mux2_1
X_3759_ _6955_/Q _5485_/B _5440_/C _3452_/X _6963_/Q VGND VGND VPWR VPWR _3759_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6478_ _3844_/Y _6478_/A1 _6480_/S VGND VGND VPWR VPWR _7226_/D sky130_fd_sc_hd__mux2_1
X_5429_ _4051_/B hold452/X _5430_/S VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput250 _7309_/X VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
Xoutput261 _6817_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
Xoutput272 _6727_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
Xoutput283 _6833_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput294 _6740_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XFILLER_114_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire355 _6239_/Y VGND VGND VPWR VPWR _6240_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_99_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire366 _6255_/Y VGND VGND VPWR VPWR _6265_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_183_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4729_/A _4970_/A _4293_/Y _4798_/X VGND VGND VPWR VPWR _4800_/X sky130_fd_sc_hd__o31a_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5780_ _6059_/S _7183_/Q _7182_/Q _6010_/C VGND VGND VPWR VPWR _5780_/X sky130_fd_sc_hd__and4_4
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4731_/A _4731_/B _4731_/C VGND VGND VPWR VPWR _4737_/C sky130_fd_sc_hd__nand3_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4662_ _4674_/C _4662_/B _4662_/C VGND VGND VPWR VPWR _4903_/B sky130_fd_sc_hd__and3_4
X_6401_ _6745_/Q _6446_/B _6143_/C _6117_/X _6594_/Q VGND VGND VPWR VPWR _6401_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3613_ _6644_/Q _5485_/B _3457_/X _3907_/B _6588_/Q VGND VGND VPWR VPWR _3613_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_175_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4593_ _4473_/Y _4525_/Y _4592_/Y _4591_/Y VGND VGND VPWR VPWR _4596_/C sky130_fd_sc_hd__o211ai_1
Xhold903 _7126_/Q VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__dlygate4sd3_1
X_6332_ _6902_/Q _6129_/A _6129_/B _6926_/Q _6331_/X VGND VGND VPWR VPWR _6339_/A
+ sky130_fd_sc_hd__a221o_1
Xhold914 _5592_/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3544_ _5494_/C _5575_/C _5575_/D VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__and3_4
Xhold925 _7094_/Q VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _6780_/Q VGND VGND VPWR VPWR hold936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 _4019_/X VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _4136_/X VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 _6822_/Q VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6263_ _7107_/Q _6112_/X _6260_/X _6262_/X VGND VGND VPWR VPWR _6264_/C sky130_fd_sc_hd__a211o_1
X_3475_ _7281_/A _3540_/B _3528_/C _3474_/X _7143_/Q VGND VGND VPWR VPWR _3475_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_142_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5214_ _4632_/B _5036_/C _4333_/A _5089_/X VGND VGND VPWR VPWR _5214_/X sky130_fd_sc_hd__a31o_1
XFILLER_130_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6194_ _7081_/Q _6177_/A _6102_/X _6104_/X _7161_/Q VGND VGND VPWR VPWR _6194_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5145_ _5238_/A _5145_/B _5238_/B VGND VGND VPWR VPWR _5146_/C sky130_fd_sc_hd__nor3_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5076_ _5073_/Y _5076_/B _5076_/C VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__and3b_1
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4027_ hold515/X _6546_/A0 _4028_/S VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5978_ _6743_/Q _6028_/C _6025_/C _5768_/X _6683_/Q VGND VGND VPWR VPWR _5978_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_40_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4929_ _4751_/A _4592_/B _4903_/A _4595_/A _4928_/Y VGND VGND VPWR VPWR _4929_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmgmt_gpio_9_buff_inst _6785_/Q VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3260_ _7074_/Q VGND VGND VPWR VPWR _3260_/Y sky130_fd_sc_hd__inv_2
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6950_ _7148_/CLK _6950_/D fanout591/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5901_ _7107_/Q _5764_/X _5784_/X _7027_/Q _5900_/X VGND VGND VPWR VPWR _5901_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6881_ _7063_/CLK _6881_/D fanout590/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5832_ _7112_/Q _5826_/B _5842_/C _5831_/X VGND VGND VPWR VPWR _5832_/X sky130_fd_sc_hd__a31o_1
XFILLER_179_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5763_ _7183_/Q _7182_/Q _5783_/C _5795_/D VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__and4_2
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4714_ _4721_/C _4683_/C _4987_/B _4668_/C VGND VGND VPWR VPWR _4729_/D sky130_fd_sc_hd__o211a_2
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5694_ _5694_/A _5694_/B VGND VGND VPWR VPWR _5694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4645_ _4645_/A _4756_/C VGND VGND VPWR VPWR _4645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold700 hold700/A VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 _5375_/X VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4576_ _4576_/A _4576_/B _4576_/C VGND VGND VPWR VPWR _4579_/A sky130_fd_sc_hd__nor3_1
Xhold722 _7149_/Q VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 _6567_/Q VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap441 _4252_/Y VGND VGND VPWR VPWR _4427_/C sky130_fd_sc_hd__buf_4
X_6315_ _6296_/X _6315_/B _6315_/C VGND VGND VPWR VPWR _6315_/Y sky130_fd_sc_hd__nand3b_4
Xhold744 _7136_/Q VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3527_ _6536_/C _6530_/D _3533_/C VGND VGND VPWR VPWR _4152_/C sky130_fd_sc_hd__and3_2
Xhold755 hold755/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_89_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7295_ _7295_/A VGND VGND VPWR VPWR _7295_/X sky130_fd_sc_hd__clkbuf_2
Xhold766 _3977_/X VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _7147_/Q VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 _3935_/X VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _7091_/Q _6106_/X _6135_/X _6939_/Q _6245_/X VGND VGND VPWR VPWR _6246_/X
+ sky130_fd_sc_hd__a221o_1
Xhold799 hold799/A VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3458_ _6829_/Q _5325_/C _3721_/A3 _7103_/Q _5611_/B VGND VGND VPWR VPWR _3458_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6177_ _6177_/A _6425_/B _6177_/C VGND VGND VPWR VPWR _6177_/X sky130_fd_sc_hd__and3_4
XFILLER_162_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1400 _6967_/Q VGND VGND VPWR VPWR hold1400/X sky130_fd_sc_hd__dlygate4sd3_1
X_3389_ _6549_/A0 _3389_/A1 _3393_/S VGND VGND VPWR VPWR _3389_/X sky130_fd_sc_hd__mux2_1
Xhold1411 _6527_/X VGND VGND VPWR VPWR _7246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _6521_/X VGND VGND VPWR VPWR _7241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _7071_/Q VGND VGND VPWR VPWR hold1433/X sky130_fd_sc_hd__dlygate4sd3_1
X_5128_ _5128_/A _5128_/B _5128_/C VGND VGND VPWR VPWR _5128_/X sky130_fd_sc_hd__and3_1
XFILLER_29_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1444 _7056_/Q VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 _6585_/Q VGND VGND VPWR VPWR _3876_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1466 _6580_/Q VGND VGND VPWR VPWR _3633_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1477 _7222_/Q VGND VGND VPWR VPWR _6474_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1488 _6418_/X VGND VGND VPWR VPWR _7217_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5059_ _4259_/Y _4356_/Y _4506_/Y _4482_/C VGND VGND VPWR VPWR _5061_/C sky130_fd_sc_hd__o31a_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1499 _3542_/B VGND VGND VPWR VPWR hold1499/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold85/X VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4430_ _4428_/Y _5044_/B _5044_/A VGND VGND VPWR VPWR _4440_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_2 _5390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4361_ _4761_/C _4320_/A _4280_/A _4683_/B VGND VGND VPWR VPWR _4870_/C sky130_fd_sc_hd__o31a_2
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6100_ _6177_/A _6130_/A _6143_/C VGND VGND VPWR VPWR _6129_/B sky130_fd_sc_hd__and3_4
X_3312_ input118/X input119/X _3312_/C _3312_/D VGND VGND VPWR VPWR _3319_/B sky130_fd_sc_hd__and4bb_1
Xfanout509 hold158/X VGND VGND VPWR VPWR hold126/A sky130_fd_sc_hd__buf_8
X_7080_ _7170_/CLK _7080_/D fanout605/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfstp_2
X_4292_ _4940_/A _4734_/B _4294_/B VGND VGND VPWR VPWR _4970_/B sky130_fd_sc_hd__and3_2
XFILLER_140_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6031_ _6755_/Q _6073_/B2 _5774_/X _6670_/Q _6030_/X VGND VGND VPWR VPWR _6031_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6933_ _7150_/CLK _6933_/D fanout602/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6864_ _7152_/CLK _6864_/D fanout587/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5815_ _6059_/S _5815_/B _5815_/C VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__and3_4
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ _7171_/CLK _6795_/D fanout610/X VGND VGND VPWR VPWR _7294_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_179_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5746_ _5746_/A _5746_/B VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__nand2_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5677_ _5494_/A _3509_/X _3915_/X _5683_/S _5677_/B2 VGND VGND VPWR VPWR _5677_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4628_ _4656_/C _4777_/A _4761_/C VGND VGND VPWR VPWR _5263_/C sky130_fd_sc_hd__and3_4
XFILLER_163_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold530 _6869_/Q VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold541 _4143_/X VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _4584_/B _5140_/C _5263_/A _4561_/B VGND VGND VPWR VPWR _4560_/B sky130_fd_sc_hd__nand4_1
XFILLER_190_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold552 _7059_/Q VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold563 _7163_/Q VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _5495_/X VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold585 hold585/A VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlygate4sd3_1
X_7278_ _7278_/CLK _7278_/D fanout595/X VGND VGND VPWR VPWR _7278_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_173_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold596 hold596/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
X_6229_ _7122_/Q _5750_/X _6117_/X _7170_/Q _6228_/X VGND VGND VPWR VPWR _6230_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1230 _6838_/Q VGND VGND VPWR VPWR _5307_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 _5289_/X VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _3876_/A1 VGND VGND VPWR VPWR hold538/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1263 _3967_/A1 VGND VGND VPWR VPWR hold621/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1274 _6479_/A1 VGND VGND VPWR VPWR hold725/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 _7045_/Q VGND VGND VPWR VPWR _5546_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_403 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1296 _7114_/Q VGND VGND VPWR VPWR _5624_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 _6028_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_425 _5815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6494_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6510_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3930_ _6539_/A0 _3930_/A1 _3932_/S VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3861_ _7045_/Q _5548_/C _5684_/C _3463_/X _7117_/Q VGND VGND VPWR VPWR _3861_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_31_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5600_ _4051_/B hold727/X hold14/X VGND VGND VPWR VPWR _5600_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6580_ _7256_/CLK _6580_/D VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfxtp_1
X_3792_ _6752_/Q _4121_/B _3562_/X _6642_/Q _3791_/X VGND VGND VPWR VPWR _3792_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5531_ _5531_/A0 _6549_/A0 _5538_/S VGND VGND VPWR VPWR _5531_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5462_ _3922_/C hold112/X _5466_/S VGND VGND VPWR VPWR _5462_/X sky130_fd_sc_hd__mux2_1
X_7201_ _7259_/CLK _7201_/D fanout595/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4413_ _4751_/A _5055_/D _5143_/A _5140_/B VGND VGND VPWR VPWR _4413_/Y sky130_fd_sc_hd__nand4_1
X_5393_ hold669/X _4051_/B _5394_/S VGND VGND VPWR VPWR _5393_/X sky130_fd_sc_hd__mux2_1
X_7132_ _7132_/CLK _7132_/D fanout610/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_1
X_4344_ _4730_/A _4674_/C VGND VGND VPWR VPWR _4344_/Y sky130_fd_sc_hd__nand2_2
X_7063_ _7063_/CLK _7063_/D fanout590/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfstp_2
X_4275_ _4632_/A _4511_/A VGND VGND VPWR VPWR _5089_/C sky130_fd_sc_hd__nand2_8
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6014_ _6598_/Q _6072_/B _6028_/B _5789_/X _6779_/Q VGND VGND VPWR VPWR _6014_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_100_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _7015_/CLK _6916_/D fanout588/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6847_ _6889_/CLK _6847_/D fanout582/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6778_ _6780_/CLK _6778_/D _3291_/A VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5729_ _5795_/D _5728_/X _5727_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__o21ai_1
XFILLER_182_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold360 _6694_/Q VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 hold371/A VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _5525_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _6541_/X VGND VGND VPWR VPWR _7269_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1060 _3986_/X VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 _6791_/Q VGND VGND VPWR VPWR _4188_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1082 _4096_/X VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _6446_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1093 _6815_/Q VGND VGND VPWR VPWR _5278_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_211 _6536_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _3922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _3915_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 hold5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _6802_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_266 _3466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 _3832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 _5767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 _5917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4060_ _3918_/X hold569/X _4065_/S VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4962_ _4692_/Y _4951_/X _4960_/X _4961_/X VGND VGND VPWR VPWR _4962_/X sky130_fd_sc_hd__o211a_1
X_6701_ _6957_/CLK _6701_/D fanout591/X VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_1
X_3913_ _6548_/B _3913_/B VGND VGND VPWR VPWR _3914_/S sky130_fd_sc_hd__nand2_2
X_4893_ _5036_/B _4970_/D _4970_/B _4892_/X VGND VGND VPWR VPWR _4893_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6632_ _7256_/CLK _6632_/D VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3844_ _3844_/A _3844_/B _3844_/C VGND VGND VPWR VPWR _3844_/Y sky130_fd_sc_hd__nand3_4
XFILLER_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6563_ _7269_/CLK _6563_/D fanout576/X VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3775_ _7264_/Q _6530_/C _3457_/X _3771_/X _3774_/X VGND VGND VPWR VPWR _3775_/X
+ sky130_fd_sc_hd__a311o_1
X_5514_ _6550_/A0 hold253/X _5520_/S VGND VGND VPWR VPWR _5514_/X sky130_fd_sc_hd__mux2_1
X_6494_ _7259_/Q _6494_/A2 _6494_/B1 _7257_/Q VGND VGND VPWR VPWR _6494_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5445_ hold418/X _3925_/C _5448_/S VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5376_ _5376_/A0 _5692_/A1 _5376_/S VGND VGND VPWR VPWR _5376_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7115_ _7129_/CLK _7115_/D fanout598/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4327_ _4320_/B _4940_/C _4691_/B VGND VGND VPWR VPWR _4327_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7046_ _7140_/CLK _7046_/D fanout609/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_2
X_4258_ _4691_/B _4427_/D _4254_/Y _4252_/Y _4427_/A VGND VGND VPWR VPWR _5060_/B
+ sky130_fd_sc_hd__o311a_4
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4189_ _4204_/S _3539_/X _4056_/Y _3369_/Y _4076_/X VGND VGND VPWR VPWR _4205_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold190 _7061_/Q VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6687_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ _6607_/Q _3558_/X _3559_/X _6903_/Q _3557_/X VGND VGND VPWR VPWR _3561_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3491_ _6536_/C _6530_/C _6536_/D VGND VGND VPWR VPWR _3954_/B sky130_fd_sc_hd__and3_4
XFILLER_127_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5230_ _4376_/Y _4633_/Y _4658_/Y _4663_/Y _4667_/Y VGND VGND VPWR VPWR _5231_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5161_ _4970_/D _4633_/B _5128_/C _4789_/D _4940_/C VGND VGND VPWR VPWR _5161_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4112_ _6524_/B _5331_/C _6536_/D _5575_/D VGND VGND VPWR VPWR _4114_/S sky130_fd_sc_hd__and4_1
XFILLER_96_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5092_ _4271_/Y _4546_/Y _5020_/C _5091_/X VGND VGND VPWR VPWR _5094_/B sky130_fd_sc_hd__o211ai_1
XFILLER_68_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4043_ _4187_/S _5341_/C hold653/X VGND VGND VPWR VPWR _4043_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5994_ _6559_/Q _6025_/B _6025_/C _5783_/X _6643_/Q VGND VGND VPWR VPWR _5994_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_64_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4945_ _4984_/A _4945_/B _4945_/C VGND VGND VPWR VPWR _4945_/X sky130_fd_sc_hd__and3_1
XFILLER_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4876_ _4876_/A _4876_/B _5109_/A VGND VGND VPWR VPWR _4879_/D sky130_fd_sc_hd__nand3_1
XFILLER_138_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6615_ _7256_/CLK _6615_/D VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfxtp_1
X_3827_ _6876_/Q _5350_/B _3499_/X _7020_/Q _3826_/X VGND VGND VPWR VPWR _3834_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6546_ _6546_/A0 hold536/X _6547_/S VGND VGND VPWR VPWR _6546_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3758_ _6672_/Q _3513_/X _5377_/C _6899_/Q VGND VGND VPWR VPWR _3758_/X sky130_fd_sc_hd__a22o_2
XFILLER_145_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6477_ _6477_/A0 _6477_/A1 _6480_/S VGND VGND VPWR VPWR _7225_/D sky130_fd_sc_hd__mux2_1
X_3689_ _6813_/Q _5341_/A _5273_/D _3498_/X _6765_/Q VGND VGND VPWR VPWR _3689_/X
+ sky130_fd_sc_hd__a32o_1
X_5428_ hold83/X hold106/X _5430_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
Xoutput240 _3324_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput251 _7310_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput262 _6818_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput273 _6728_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_160_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput284 _6834_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
X_5359_ hold13/X _5359_/B VGND VGND VPWR VPWR _5367_/S sky130_fd_sc_hd__nand2_8
Xoutput295 _6725_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7029_ _7161_/CLK _7029_/D fanout600/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_55_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__1184_ clkbuf_0__1184_/X VGND VGND VPWR VPWR _6477_/A0 sky130_fd_sc_hd__clkbuf_16
Xwire356 _6214_/Y VGND VGND VPWR VPWR _6215_/C sky130_fd_sc_hd__clkbuf_1
Xwire367 _6230_/Y VGND VGND VPWR VPWR _6240_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_137_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4730_ _4730_/A _4777_/B _4730_/C _4730_/D VGND VGND VPWR VPWR _4731_/C sky130_fd_sc_hd__nand4_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ _4970_/D _5128_/C _4755_/D VGND VGND VPWR VPWR _4661_/X sky130_fd_sc_hd__and3_1
X_6400_ _6680_/Q _6122_/X _6452_/B1 _6755_/Q _6399_/X VGND VGND VPWR VPWR _6405_/B
+ sky130_fd_sc_hd__a221o_1
X_3612_ _7072_/Q _3488_/X _3603_/X _3604_/X _3611_/X VGND VGND VPWR VPWR _3631_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4592_ _4751_/A _4592_/B VGND VGND VPWR VPWR _4592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6331_ _7094_/Q _6136_/A _6102_/X _6113_/X _7150_/Q VGND VGND VPWR VPWR _6331_/X
+ sky130_fd_sc_hd__a32o_1
Xhold904 _5638_/X VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3543_ _7260_/Q _6530_/C _5325_/C VGND VGND VPWR VPWR _3543_/X sky130_fd_sc_hd__and3_1
Xhold915 _6782_/Q VGND VGND VPWR VPWR hold915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _5601_/X VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _4161_/X VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold948 _6921_/Q VGND VGND VPWR VPWR hold948/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold959 hold959/A VGND VGND VPWR VPWR hold959/X sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _6923_/Q _6129_/B _6110_/X _7115_/Q _6261_/X VGND VGND VPWR VPWR _6262_/X
+ sky130_fd_sc_hd__a221o_1
X_3474_ _5666_/C _5476_/C _5575_/C VGND VGND VPWR VPWR _3474_/X sky130_fd_sc_hd__and3_4
X_5213_ _4333_/A _4786_/B _5036_/A _4738_/B _5036_/X VGND VGND VPWR VPWR _5216_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6193_ _6192_/X _6217_/A2 _6443_/S VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5144_ _4259_/Y _4356_/Y _5132_/Y _5143_/Y _4814_/Y VGND VGND VPWR VPWR _5238_/B
+ sky130_fd_sc_hd__o311ai_2
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5075_ _4946_/X _4633_/Y _4613_/Y _5248_/A3 _4692_/Y VGND VGND VPWR VPWR _5076_/C
+ sky130_fd_sc_hd__a311o_1
X_4026_ hold978/X _6539_/A0 _4028_/S VGND VGND VPWR VPWR _4026_/X sky130_fd_sc_hd__mux2_1
X_7191__627 VGND VGND VPWR VPWR _7191_/D _7191__627/LO sky130_fd_sc_hd__conb_1
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _5977_/A1 _5761_/X _5976_/X _5975_/X VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4928_ _4928_/A _5100_/A _4928_/C VGND VGND VPWR VPWR _4928_/Y sky130_fd_sc_hd__nand3_1
XFILLER_178_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4859_ _4859_/A _4984_/C _4859_/C _4859_/D VGND VGND VPWR VPWR _4859_/Y sky130_fd_sc_hd__nand4_1
XFILLER_21_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6529_ _6535_/A0 _6529_/A1 _6529_/S VGND VGND VPWR VPWR _6529_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7073_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6768_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_csclk _7277_/CLK VGND VGND VPWR VPWR _7275_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7162_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5900_ _7115_/Q _6059_/S _5842_/C _5780_/X _7099_/Q VGND VGND VPWR VPWR _5900_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6880_ _7088_/CLK _6880_/D fanout591/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5831_ _7072_/Q _5971_/A2 _5813_/X _7056_/Q _5830_/X VGND VGND VPWR VPWR _5831_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5762_ _7181_/Q _7180_/Q VGND VGND VPWR VPWR _5783_/C sky130_fd_sc_hd__and2b_4
XFILLER_148_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4713_ _4208_/Y _4246_/Y _5089_/C _4371_/Y _4372_/Y VGND VGND VPWR VPWR _4987_/B
+ sky130_fd_sc_hd__o311a_4
X_5693_ _6803_/Q _6800_/Q VGND VGND VPWR VPWR _5694_/B sky130_fd_sc_hd__nand2b_1
XFILLER_187_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4644_ _4756_/C _4760_/B _4742_/C VGND VGND VPWR VPWR _4682_/B sky130_fd_sc_hd__and3_2
Xhold701 hold701/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
X_4575_ _5140_/C _4575_/B _4589_/C VGND VGND VPWR VPWR _4576_/B sky130_fd_sc_hd__and3_1
Xmax_cap420 _6025_/C VGND VGND VPWR VPWR _5911_/C sky130_fd_sc_hd__buf_8
Xhold712 _7112_/Q VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 _5664_/X VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3526_ _7119_/Q hold17/A _3902_/A3 _4121_/B _6748_/Q VGND VGND VPWR VPWR _3526_/X
+ sky130_fd_sc_hd__a32o_1
Xhold734 _3383_/X VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6314_ _6314_/A _6314_/B _6314_/C _6440_/D VGND VGND VPWR VPWR _6314_/Y sky130_fd_sc_hd__nor4_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold745 _5650_/X VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7294_ _7294_/A VGND VGND VPWR VPWR _7294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold756 _7137_/Q VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _6872_/Q VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold778 _5662_/X VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6245_ hold61/A _6097_/X _6452_/B1 _6979_/Q _6244_/X VGND VGND VPWR VPWR _6245_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3457_ _5324_/B hold37/X hold42/X _6548_/C VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__and4_4
Xhold789 _6644_/Q VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6176_ _6992_/Q _6176_/B _6347_/C VGND VGND VPWR VPWR _6176_/X sky130_fd_sc_hd__and3_1
X_3388_ _3987_/A _6548_/A _6548_/B _5630_/C VGND VGND VPWR VPWR _3393_/S sky130_fd_sc_hd__nand4_4
Xhold1401 _5459_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 _6951_/Q VGND VGND VPWR VPWR hold1412/X sky130_fd_sc_hd__dlygate4sd3_1
X_5127_ _5008_/X _5127_/B _5127_/C VGND VGND VPWR VPWR _5127_/Y sky130_fd_sc_hd__nand3b_1
Xhold1423 _7104_/Q VGND VGND VPWR VPWR hold762/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _5576_/X VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 _5559_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1456 _6632_/Q VGND VGND VPWR VPWR _3968_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1467 _6944_/Q VGND VGND VPWR VPWR hold375/A sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _5058_/A _5131_/B _5058_/C VGND VGND VPWR VPWR _5061_/A sky130_fd_sc_hd__and3_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1478 _6582_/Q VGND VGND VPWR VPWR _3754_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1489 _6615_/Q VGND VGND VPWR VPWR _3949_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ hold513/X _6546_/A0 _4010_/S VGND VGND VPWR VPWR _4009_/X sky130_fd_sc_hd__mux2_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__buf_12
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 _7085_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4360_ _4246_/Y _4280_/A _4662_/B VGND VGND VPWR VPWR _4683_/B sky130_fd_sc_hd__o21ai_2
X_3311_ _4637_/A _4747_/A _4747_/B _4747_/C VGND VGND VPWR VPWR _4214_/A sky130_fd_sc_hd__a211o_4
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4291_ _4637_/A _4747_/B _4747_/C _4760_/B VGND VGND VPWR VPWR _4799_/B sky130_fd_sc_hd__nor4_4
X_6030_ _6685_/Q _5768_/X _5794_/X _6660_/Q _6029_/X VGND VGND VPWR VPWR _6030_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6932_ _7117_/CLK _6932_/D fanout608/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6863_ _7071_/CLK _6863_/D fanout585/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5814_ _6059_/S _5815_/C _5814_/C VGND VGND VPWR VPWR _5814_/X sky130_fd_sc_hd__and3_4
X_6794_ _7171_/CLK _6794_/D fanout609/X VGND VGND VPWR VPWR _7293_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_167_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5745_ _5741_/Y _5752_/B2 _7189_/Q _5712_/Y VGND VGND VPWR VPWR _5746_/B sky130_fd_sc_hd__a211o_1
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5676_ _6549_/A0 _5676_/A1 _5683_/S VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__mux2_1
X_4627_ _4860_/C _4859_/D _4675_/B _4860_/B VGND VGND VPWR VPWR _4720_/D sky130_fd_sc_hd__nand4_1
Xhold520 hold520/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4558_ _5140_/C _4561_/B VGND VGND VPWR VPWR _4558_/Y sky130_fd_sc_hd__nand2_1
Xhold531 _5348_/X VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _7301_/A VGND VGND VPWR VPWR hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold553 _5562_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold564 _5680_/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3509_ _5449_/B _5684_/B _5675_/D VGND VGND VPWR VPWR _3509_/X sky130_fd_sc_hd__and3_4
Xhold575 _6652_/Q VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold586 hold586/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
X_7277_ _7277_/CLK _7277_/D fanout594/X VGND VGND VPWR VPWR _7277_/Q sky130_fd_sc_hd__dfstp_2
X_4489_ _4632_/B _4612_/C _4489_/C VGND VGND VPWR VPWR _5140_/C sky130_fd_sc_hd__and3_4
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold597 hold597/A VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6228_ _6946_/Q _6347_/C _6139_/X _6113_/X _7146_/Q VGND VGND VPWR VPWR _6228_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6159_ _6991_/Q _6176_/B _6347_/C _6113_/X _7143_/Q VGND VGND VPWR VPWR _6159_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 _6743_/Q VGND VGND VPWR VPWR _4116_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _5307_/X VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1242 _6678_/Q VGND VGND VPWR VPWR _4024_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 _3948_/A1 VGND VGND VPWR VPWR hold557/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1264 _3966_/A1 VGND VGND VPWR VPWR hold617/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 _3965_/A1 VGND VGND VPWR VPWR hold589/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _6956_/Q VGND VGND VPWR VPWR _5446_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_404 _6143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1297 _7098_/Q VGND VGND VPWR VPWR _5606_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_415 _5795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_426 _6109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6492_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6497_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6487_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3860_ input41/X _4187_/S _3469_/X input9/X _3859_/X VGND VGND VPWR VPWR _3874_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3791_ _6979_/Q _5494_/C _5281_/A2 _3790_/X VGND VGND VPWR VPWR _3791_/X sky130_fd_sc_hd__a31o_1
XFILLER_176_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ hold8/X _5548_/C _6548_/D _5675_/D VGND VGND VPWR VPWR _5538_/S sky130_fd_sc_hd__and4_4
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5461_ hold2/X _5461_/A1 _5466_/S VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__mux2_1
XFILLER_172_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7200_ _7259_/CLK _7200_/D fanout595/X VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_1
X_4412_ _5055_/D _5140_/B VGND VGND VPWR VPWR _4412_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5392_ hold258/X _4049_/B _5394_/S VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__mux2_1
X_4343_ _4656_/C _4730_/A _4761_/C VGND VGND VPWR VPWR _4788_/A sky130_fd_sc_hd__and3_4
XFILLER_98_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7131_ _7131_/CLK hold10/X fanout606/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7062_ _7157_/CLK _7062_/D fanout593/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4274_ _4698_/A _4657_/C _4656_/C _4647_/C VGND VGND VPWR VPWR _4799_/A sky130_fd_sc_hd__nor4b_4
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6013_ _7276_/Q _6086_/B1 _5784_/X _6621_/Q VGND VGND VPWR VPWR _6013_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6915_ _7063_/CLK _6915_/D fanout590/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_4
X_6846_ _7067_/CLK _6846_/D fanout582/X VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6777_ _7239_/CLK _6777_/D fanout574/X VGND VGND VPWR VPWR _6777_/Q sky130_fd_sc_hd__dfrtp_4
X_3989_ _6550_/A0 hold784/X _3992_/S VGND VGND VPWR VPWR _3989_/X sky130_fd_sc_hd__mux2_1
X_5728_ _6800_/Q _5759_/B _5782_/C _5795_/C VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__o211a_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5659_ _5494_/A _3474_/X _3915_/X _5665_/S _5659_/B2 VGND VGND VPWR VPWR _5659_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold350 _6587_/Q VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold361 _4045_/X VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold372 hold372/A VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _7274_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _6947_/Q VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1050 _7038_/Q VGND VGND VPWR VPWR _5538_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1061 _6642_/Q VGND VGND VPWR VPWR _3980_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _4188_/X VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 _6727_/Q VGND VGND VPWR VPWR _4097_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1094 _5278_/X VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _6446_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _6543_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _3922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_234 _3340_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _3246_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 _3466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 _3915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 _5768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4961_ _4271_/Y _5248_/A3 _4699_/Y _4745_/Y _4692_/Y VGND VGND VPWR VPWR _4961_/X
+ sky130_fd_sc_hd__o32a_1
X_6700_ _7077_/CLK _6700_/D fanout587/X VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_1
X_3912_ _3924_/B hold444/X _3912_/S VGND VGND VPWR VPWR _3912_/X sky130_fd_sc_hd__mux2_1
X_4892_ _5128_/A _4859_/C _4729_/D _4891_/X VGND VGND VPWR VPWR _4892_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6631_ _7219_/CLK _6631_/D VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3843_ _3843_/A _3843_/B _3843_/C _3843_/D VGND VGND VPWR VPWR _3843_/Y sky130_fd_sc_hd__nor4_1
X_6562_ _7268_/CLK _6562_/D fanout572/X VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfrtp_4
X_3774_ _6647_/Q _5273_/D _5325_/C _3773_/X VGND VGND VPWR VPWR _3774_/X sky130_fd_sc_hd__a31o_1
XFILLER_192_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5513_ _5667_/A0 _5513_/A1 _5520_/S VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__mux2_1
X_6493_ _6492_/X _6550_/A0 _6511_/S VGND VGND VPWR VPWR _7230_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ hold666/X _3921_/B _5448_/S VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__mux2_1
X_5375_ hold710/X _4051_/B _5376_/S VGND VGND VPWR VPWR _5375_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7114_ _7114_/CLK hold25/X fanout604/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4326_ _4321_/Y _4322_/Y _4325_/Y VGND VGND VPWR VPWR _4606_/B sky130_fd_sc_hd__a21oi_4
XFILLER_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7045_ _7162_/CLK hold78/X fanout602/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfrtp_4
X_4257_ _4427_/D _4320_/A _4657_/C _4249_/Y VGND VGND VPWR VPWR _4429_/A sky130_fd_sc_hd__o22ai_4
XFILLER_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4188_ _4188_/A0 _4187_/X _4188_/S VGND VGND VPWR VPWR _4188_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6829_ _6855_/CLK _6829_/D fanout584/X VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold180 _6916_/Q VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _5564_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3490_ _7071_/Q _3488_/X _3489_/X _6911_/Q _3487_/X VGND VGND VPWR VPWR _3507_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5160_ _5153_/X _4709_/Y _4963_/X _5079_/B VGND VGND VPWR VPWR _5249_/A sky130_fd_sc_hd__o211a_1
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4111_ _4053_/B hold160/X _4111_/S VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__mux2_1
X_5091_ _4522_/Y _4613_/Y _4658_/Y _4554_/B _4554_/C VGND VGND VPWR VPWR _5091_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4042_ _4055_/A1 _6898_/Q _3346_/D hold66/A _4187_/S VGND VGND VPWR VPWR _4054_/S
+ sky130_fd_sc_hd__o311a_4
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5993_ _6763_/Q _5770_/X _5979_/X _5989_/X _5992_/X VGND VGND VPWR VPWR _5993_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_18_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4944_ _4691_/B _4761_/C _4698_/A _4870_/B VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__a211o_1
X_4875_ _4376_/Y _4629_/Y _4633_/Y _4456_/C VGND VGND VPWR VPWR _5109_/A sky130_fd_sc_hd__o31a_1
X_6614_ _7256_/CLK _6614_/D VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3826_ _7044_/Q _5548_/C _5281_/A2 _3463_/X _7116_/Q VGND VGND VPWR VPWR _3826_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6545_ _3919_/C hold328/X _6547_/S VGND VGND VPWR VPWR _6545_/X sky130_fd_sc_hd__mux2_1
X_3757_ hold65/A _6805_/Q _5657_/D _3757_/D VGND VGND VPWR VPWR _3757_/X sky130_fd_sc_hd__and4_1
XFILLER_118_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6476_ _3753_/X _6476_/A1 _6480_/S VGND VGND VPWR VPWR _7224_/D sky130_fd_sc_hd__mux2_1
X_3688_ _6566_/Q _5311_/B _6530_/C _3687_/X VGND VGND VPWR VPWR _3688_/X sky130_fd_sc_hd__a31o_1
XFILLER_133_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput230 _7302_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
X_5427_ _3925_/C hold358/X _5430_/S VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__mux2_1
Xoutput241 _3323_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
Xoutput252 _3292_/Y VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput263 _6819_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
Xoutput274 _6729_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput285 _6835_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ _6511_/A1 hold264/X _5358_/S VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput296 _6726_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_102_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4309_ _4310_/B _4310_/C _4310_/D _4747_/A VGND VGND VPWR VPWR _4318_/A sky130_fd_sc_hd__a31o_1
X_5289_ _5289_/A0 _4152_/B _5294_/S VGND VGND VPWR VPWR _5289_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7028_ _7117_/CLK _7028_/D fanout608/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire346 _3631_/Y VGND VGND VPWR VPWR _3632_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_183_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire357 _6181_/Y VGND VGND VPWR VPWR wire357/X sky130_fd_sc_hd__clkbuf_1
Xwire368 _6165_/Y VGND VGND VPWR VPWR wire368/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout490 hold17/X VGND VGND VPWR VPWR _6536_/A sky130_fd_sc_hd__buf_12
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4660_ _4653_/B _4712_/B _4659_/B _4860_/B _5255_/A VGND VGND VPWR VPWR _4672_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_174_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3611_ _7048_/Q _3548_/X _3605_/X _3606_/X _3610_/X VGND VGND VPWR VPWR _3611_/X
+ sky130_fd_sc_hd__a2111o_1
X_4591_ _4591_/A _4591_/B _4591_/C VGND VGND VPWR VPWR _4591_/Y sky130_fd_sc_hd__nor3_1
X_6330_ _6330_/A _6330_/B _6330_/C _6330_/D VGND VGND VPWR VPWR _6340_/B sky130_fd_sc_hd__nor4_2
XFILLER_128_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3542_ _5630_/C _3542_/B hold28/A VGND VGND VPWR VPWR _5413_/B sky130_fd_sc_hd__and3_4
Xhold905 _7030_/Q VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 _4163_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _7046_/Q VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _6682_/Q VGND VGND VPWR VPWR hold938/X sky130_fd_sc_hd__dlygate4sd3_1
X_3473_ input34/X _3469_/X _3470_/X _7244_/Q _3472_/X VGND VGND VPWR VPWR _3485_/B
+ sky130_fd_sc_hd__a221o_1
Xhold949 _5407_/X VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6261_ _7011_/Q _6117_/C _6096_/Y _6137_/X _7099_/Q VGND VGND VPWR VPWR _6261_/X
+ sky130_fd_sc_hd__a32o_1
X_5212_ hold54/A wire442/X _5211_/Y _5202_/X VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__a211o_1
XFILLER_143_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6192_ _6191_/X _6192_/A1 _6292_/S VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5143_ _5143_/A _5260_/B _5143_/C _5143_/D VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__nand4_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5074_ _4946_/X _4633_/Y _4613_/Y _4629_/Y _5248_/A3 VGND VGND VPWR VPWR _5076_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4025_ hold478/X _6538_/A0 _4028_/S VGND VGND VPWR VPWR _4025_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5976_ _6292_/S _7200_/Q _6343_/S VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4927_ _4490_/Y _4601_/Y _4525_/Y VGND VGND VPWR VPWR _4928_/C sky130_fd_sc_hd__a21o_1
X_4858_ _5255_/A _4676_/X _4850_/X _4857_/X VGND VGND VPWR VPWR _4864_/B sky130_fd_sc_hd__a211oi_1
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ _3353_/B _4187_/S _3797_/X _3800_/X _3808_/X VGND VGND VPWR VPWR _3810_/D
+ sky130_fd_sc_hd__a2111o_2
XFILLER_119_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4789_ _4940_/C _4789_/B _5128_/C _4789_/D VGND VGND VPWR VPWR _4790_/B sky130_fd_sc_hd__nand4_1
XFILLER_165_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6528_ _6540_/A0 hold605/X _6529_/S VGND VGND VPWR VPWR _6528_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6689_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6459_ _7279_/Q _6444_/C _5750_/C _6105_/X _6606_/Q VGND VGND VPWR VPWR _6459_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5830_ _7040_/Q _5826_/B _6028_/B _5970_/B1 _6928_/Q VGND VGND VPWR VPWR _5830_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_179_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5761_ _6292_/S _3307_/B _5759_/X VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__a21o_4
X_4712_ _4862_/A _4712_/B _4792_/C _4860_/B VGND VGND VPWR VPWR _4717_/A sky130_fd_sc_hd__and4_1
XFILLER_187_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5692_ hold960/X _5692_/A1 _5692_/S VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4643_ _4699_/B _4674_/D VGND VGND VPWR VPWR _4643_/Y sky130_fd_sc_hd__nand2_2
XFILLER_162_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4574_ _4815_/A _4575_/B _4574_/C VGND VGND VPWR VPWR _4576_/A sky130_fd_sc_hd__and3_1
Xhold702 _6901_/Q VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _5622_/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold724 hold724/A VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _6973_/Q _6097_/X _6310_/X _6312_/X VGND VGND VPWR VPWR _6314_/C sky130_fd_sc_hd__a211o_1
XFILLER_143_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold735 _6858_/Q VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlygate4sd3_1
X_3525_ _5630_/A _5630_/C hold28/A VGND VGND VPWR VPWR _3525_/X sky130_fd_sc_hd__and3_4
Xmax_cap443 _4165_/Y VGND VGND VPWR VPWR _4170_/B sky130_fd_sc_hd__clkbuf_2
Xhold746 _7276_/Q VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__dlygate4sd3_1
X_7293_ _7293_/A VGND VGND VPWR VPWR _7293_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold757 _5651_/X VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 _5352_/X VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6244_ _6995_/Q _6176_/B _6347_/C _6113_/X _7147_/Q VGND VGND VPWR VPWR _6244_/X
+ sky130_fd_sc_hd__a32o_1
Xhold779 _7048_/Q VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap498 _6138_/A VGND VGND VPWR VPWR _6130_/A sky130_fd_sc_hd__buf_12
X_3456_ _5620_/A _5630_/A hold28/A VGND VGND VPWR VPWR _5611_/B sky130_fd_sc_hd__and3_4
XFILLER_103_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3387_ _5304_/A _6530_/D VGND VGND VPWR VPWR _3387_/Y sky130_fd_sc_hd__nand2_1
X_6175_ _6912_/Q _6451_/B1 _6122_/X _6888_/Q VGND VGND VPWR VPWR _6175_/X sky130_fd_sc_hd__a22o_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1402 _6566_/Q VGND VGND VPWR VPWR hold979/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _5441_/X VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5126_ _4271_/Y _4391_/Y _4715_/Y _4290_/Y VGND VGND VPWR VPWR _5127_/C sky130_fd_sc_hd__a211o_1
Xhold1424 _6745_/Q VGND VGND VPWR VPWR hold743/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1435 _6809_/Q VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 _7007_/Q VGND VGND VPWR VPWR hold1446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 _7221_/Q VGND VGND VPWR VPWR _6473_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _6613_/Q VGND VGND VPWR VPWR _3947_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5057_ _5040_/A _4466_/X _5056_/X VGND VGND VPWR VPWR _5131_/B sky130_fd_sc_hd__o21ba_1
Xhold1479 _7255_/Q VGND VGND VPWR VPWR _7252_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4008_ hold975/X _6539_/A0 _4010_/S VGND VGND VPWR VPWR _4008_/X sky130_fd_sc_hd__mux2_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ _6918_/Q _5959_/B _5959_/C VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__and3_1
XFILLER_187_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_4 _7232_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3310_ _4747_/B _4747_/C VGND VGND VPWR VPWR _4940_/A sky130_fd_sc_hd__nor2_2
X_4290_ _4859_/A _4667_/C _4667_/D VGND VGND VPWR VPWR _4290_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6931_ _7120_/CLK _6931_/D fanout610/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6862_ _7129_/CLK _6862_/D fanout606/X VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5813_ _6072_/B _7181_/Q _7180_/Q _5814_/C VGND VGND VPWR VPWR _5813_/X sky130_fd_sc_hd__and4_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6793_ _7171_/CLK _6793_/D fanout609/X VGND VGND VPWR VPWR _7292_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5744_ _5752_/B2 _6446_/B _7189_/Q VGND VGND VPWR VPWR _5746_/A sky130_fd_sc_hd__a21bo_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5675_ _6548_/B _6548_/D _5684_/B _5675_/D VGND VGND VPWR VPWR _5683_/S sky130_fd_sc_hd__nand4_4
Xclkbuf_leaf_72_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7071_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4626_ _4859_/C _4859_/D _4675_/B VGND VGND VPWR VPWR _4626_/X sky130_fd_sc_hd__and3_1
Xhold510 _7305_/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold521 hold521/A VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _4557_/A _4557_/B _4674_/D VGND VGND VPWR VPWR _4557_/X sky130_fd_sc_hd__and3_1
Xhold532 _6650_/Q VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold543 _4069_/X VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 hold554/A VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _3508_/A _3508_/B _3508_/C _3508_/D VGND VGND VPWR VPWR _3568_/A sky130_fd_sc_hd__and4_1
XFILLER_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold565 _6708_/Q VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_87_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7269_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7276_ _7279_/CLK _7276_/D fanout597/X VGND VGND VPWR VPWR _7276_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_171_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold576 _3992_/X VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _4760_/C _4488_/B _4488_/C VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__and3_1
Xhold587 _6671_/Q VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold598 hold598/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6227_ _7090_/Q _6106_/X _6118_/X _7058_/Q _6226_/X VGND VGND VPWR VPWR _6230_/C
+ sky130_fd_sc_hd__a221o_1
X_3439_ _6648_/Q _5304_/A hold17/A _6536_/D VGND VGND VPWR VPWR _3439_/X sky130_fd_sc_hd__and4_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6903_/Q _6129_/D _6146_/X _6148_/X _6157_/X VGND VGND VPWR VPWR _6158_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _7282_/A VGND VGND VPWR VPWR _4083_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _4116_/X VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_10_csclk _7277_/CLK VGND VGND VPWR VPWR _7240_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1232 _6723_/Q VGND VGND VPWR VPWR _4091_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 _4024_/X VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _5109_/A _5109_/B _5109_/C VGND VGND VPWR VPWR _5194_/B sky130_fd_sc_hd__and3_1
XFILLER_73_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6089_ _5726_/Y _6692_/Q _6088_/X _6078_/X _5759_/A VGND VGND VPWR VPWR _6089_/X
+ sky130_fd_sc_hd__o221a_1
Xhold1254 _3952_/A1 VGND VGND VPWR VPWR hold548/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1265 _3949_/A1 VGND VGND VPWR VPWR hold629/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1276 _3813_/A1 VGND VGND VPWR VPWR hold643/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 _6840_/Q VGND VGND VPWR VPWR _5309_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _6945_/Q VGND VGND VPWR VPWR _5434_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_405 _6143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_416 _4127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_427 _6636_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4229_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6494_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6500_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6491_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3790_ _7243_/Q _6536_/A _5325_/C _3470_/X _7248_/Q VGND VGND VPWR VPWR _3790_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_188_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5460_ _3916_/C hold343/X _5466_/S VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4411_ _4878_/A _4411_/B VGND VGND VPWR VPWR _4444_/B sky130_fd_sc_hd__nand2_1
X_5391_ hold473/X _3925_/C _5394_/S VGND VGND VPWR VPWR _5391_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7130_ _7130_/CLK hold53/X fanout600/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfrtp_4
X_4342_ _4647_/C _4656_/C VGND VGND VPWR VPWR _4674_/C sky130_fd_sc_hd__and2b_4
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7061_ _7160_/CLK _7061_/D fanout592/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_2
X_4273_ _4656_/C _4761_/C VGND VGND VPWR VPWR _4777_/B sky130_fd_sc_hd__nor2_2
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6012_ _6588_/Q _5814_/X _5815_/X _6639_/Q _6011_/X VGND VGND VPWR VPWR _6012_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_141_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

