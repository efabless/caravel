* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1 vccd2 vssd vssd1 vssd2 vccd2_uq0 vccd2_uq1
+ vccd2_uq2 vccd2_uq3 vccd2_uq4 vccd2_uq5 vccd2_uq6 vccd1_uq0 vccd1_uq1 vccd1_uq2
+ vccd1_uq3 vccd1_uq4 vccd1_uq5 vssd2_uq0 vssd2_uq1 vssd2_uq2 vssd2_uq3 vssd2_uq4
+ vssd2_uq5 vssd1_uq0 vssd1_uq1 vssd1_uq2 vssd1_uq4 vdda2_uq0 vdda1_uq0
XTAP_177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[72\] input229/X mprj_logic_high_inst/HI[402] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[72\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input127_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[50\] _642_/A la_buf_enable\[50\]/B vssd vssd vccd vccd la_buf\[50\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_501_ _501_/A vssd vssd vccd vccd _501_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ _432_/A vssd vssd vccd vccd _432_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_363_ _363_/A vssd vssd vccd vccd _363_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input92_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[36\] _500_/Y la_buf\[36\]/TE vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_6_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[108\] input141/X mprj_logic_high_inst/HI[438] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[108\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_10_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] user_to_mprj_in_gates\[25\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_47_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput467 output467/A vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_2
Xoutput478 output478/A vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_2
XFILLER_47_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput489 output489/A vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_2
XFILLER_9_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[76\] _339_/Y mprj_logic_high_inst/HI[278] vssd vssd vccd
+ vccd la_oenb_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_2_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[98\] _361_/A la_buf_enable\[98\]/B vssd vssd vccd vccd la_buf\[98\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[24\] _456_/Y mprj_dat_buf\[24\]/TE vssd vssd vccd vccd mprj_dat_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input244_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input411_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _415_/A vssd vssd vccd vccd _415_/Y sky130_fd_sc_hd__inv_12
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_346_ _346_/A vssd vssd vccd vccd _346_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_35_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[4\] _596_/A la_buf_enable\[4\]/B vssd vssd vccd vccd la_buf\[4\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[35\] input188/X mprj_logic_high_inst/HI[365] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[35\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[13\] _605_/A la_buf_enable\[13\]/B vssd vssd vccd vccd la_buf\[13\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input194_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input361_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input459_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input55_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[92\]_A_N _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[30\]_A_N _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_329_ _329_/A vssd vssd vccd vccd _329_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[45\]_A_N _637_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] user_to_mprj_in_gates\[92\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[109\] _372_/Y mprj_logic_high_inst/HI[311] vssd vssd vccd
+ vccd la_oenb_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_29_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[39\] _631_/Y mprj_logic_high_inst/HI[241] vssd vssd vccd
+ vccd la_oenb_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_28_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input207_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__402__A _402_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd vssd vccd vccd output549/A
+ sky130_fd_sc_hd__inv_2
XFILLER_50_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[20\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[80\] _343_/A la_buf_enable\[80\]/B vssd vssd vccd vccd la_buf\[80\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput301 la_oenb_mprj[21] vssd vssd vccd vccd _613_/A sky130_fd_sc_hd__buf_2
Xinput312 la_oenb_mprj[31] vssd vssd vccd vccd _623_/A sky130_fd_sc_hd__buf_2
XANTENNA_input157_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput345 la_oenb_mprj[61] vssd vssd vccd vccd _653_/A sky130_fd_sc_hd__buf_2
Xinput334 la_oenb_mprj[51] vssd vssd vccd vccd _643_/A sky130_fd_sc_hd__buf_2
Xinput323 la_oenb_mprj[41] vssd vssd vccd vccd _633_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput356 la_oenb_mprj[71] vssd vssd vccd vccd _334_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input324_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput367 la_oenb_mprj[81] vssd vssd vccd vccd _344_/A sky130_fd_sc_hd__buf_4
Xinput378 la_oenb_mprj[91] vssd vssd vccd vccd _354_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input18_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput389 mprj_adr_o_core[10] vssd vssd vccd vccd _410_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[66\] _530_/Y la_buf\[66\]/TE vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__einvp_8
XFILLER_44_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A vssd vssd vccd vccd _594_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_38_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _586_/Y la_buf\[122\]/TE vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__einvp_8
XFILLER_6_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] user_to_mprj_in_gates\[55\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input274_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input441_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput120 la_data_out_mprj[8] vssd vssd vccd vccd _472_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput131 la_data_out_mprj[9] vssd vssd vccd vccd _473_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput142 la_iena_mprj[109] vssd vssd vccd vccd input142/X sky130_fd_sc_hd__clkbuf_1
Xinput153 la_iena_mprj[119] vssd vssd vccd vccd input153/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput164 la_iena_mprj[13] vssd vssd vccd vccd input164/X sky130_fd_sc_hd__clkbuf_1
Xinput175 la_iena_mprj[23] vssd vssd vccd vccd input175/X sky130_fd_sc_hd__clkbuf_1
Xinput186 la_iena_mprj[33] vssd vssd vccd vccd input186/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput197 la_iena_mprj[43] vssd vssd vccd vccd input197/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_646_ _646_/A vssd vssd vccd vccd _646_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_577_ _577_/A vssd vssd vccd vccd _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[6\]_A _438_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd vssd vccd vccd output508/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput627 output627/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_2
Xoutput605 output605/A vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_2
Xoutput616 output616/A vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_2
XFILLER_12_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[65\] input221/X mprj_logic_high_inst/HI[395] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[65\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_500_ _500_/A vssd vssd vccd vccd _500_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[21\] _613_/Y mprj_logic_high_inst/HI[223] vssd vssd vccd
+ vccd la_oenb_core[21] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[3\] _595_/Y mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd la_oenb_core[3] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[43\] _635_/A la_buf_enable\[43\]/B vssd vssd vccd vccd la_buf\[43\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_431_ _431_/A vssd vssd vccd vccd _431_/Y sky130_fd_sc_hd__inv_8
XFILLER_53_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_362_ _362_/A vssd vssd vccd vccd _362_/Y sky130_fd_sc_hd__inv_2
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input391_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input85_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[29\] _493_/Y la_buf\[29\]/TE vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_13_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_629_ _629_/A vssd vssd vccd vccd _629_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] user_to_mprj_in_gates\[18\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[28\] user_wb_dat_gates\[28\]/Y vssd vssd vccd vccd output612/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput468 output468/A vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_2
XFILLER_25_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput479 output479/A vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_2
XFILLER_9_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[69\] _332_/Y mprj_logic_high_inst/HI[271] vssd vssd vccd
+ vccd la_oenb_core[69] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[17\] _449_/Y mprj_dat_buf\[17\]/TE vssd vssd vccd vccd mprj_dat_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input237_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input404_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_414_ _414_/A vssd vssd vccd vccd _414_/Y sky130_fd_sc_hd__clkinv_8
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _345_/A vssd vssd vccd vccd _345_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[120\] input155/X mprj_logic_high_inst/HI[450] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[120\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[12\] _412_/Y mprj_adr_buf\[12\]/TE vssd vssd vccd vccd mprj_adr_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd vssd vccd vccd
+ output492/A sky130_fd_sc_hd__clkinv_4
XFILLER_29_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd vssd vccd vccd output582/A
+ sky130_fd_sc_hd__inv_2
XFILLER_2_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output623_A output623/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[122\]_B mprj_logic_high_inst/HI[452] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[2\] user_wb_dat_gates\[2\]/Y vssd vssd vccd vccd output614/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_33_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[41\]_B la_buf_enable\[41\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_B mprj_logic_high_inst/HI[443] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[28\] input180/X mprj_logic_high_inst/HI[358] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[28\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input187_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[32\]_B la_buf_enable\[32\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input354_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input48_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[111\] _374_/A la_buf_enable\[111\]/B vssd vssd vccd vccd la_buf\[111\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_ena_buf\[1\] input171/X mprj_logic_high_inst/HI[331] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[1\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[96\] _560_/Y la_buf\[96\]/TE vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__einvp_8
XFILLER_46_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[104\]_B mprj_logic_high_inst/HI[434] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[99\]_B la_buf_enable\[99\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[23\]_B la_buf_enable\[23\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] user_to_mprj_in_gates\[85\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[14\]_B la_buf_enable\[14\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[93\]_B mprj_logic_high_inst/HI[423] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input102_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[7\] _471_/Y la_buf\[7\]/TE vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_49_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[11\] _475_/Y la_buf\[11\]/TE vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__einvp_8
XFILLER_4_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[4\] _404_/Y mprj_adr_buf\[4\]/TE vssd vssd vccd vccd mprj_adr_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[84\]_B mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd vssd vccd vccd output541/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_37_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[13\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[10\] user_wb_dat_gates\[10\]/Y vssd vssd vccd vccd output593/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_48_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] user_to_mprj_in_gates\[111\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[91\]_A_N _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[95\] input254/X mprj_logic_high_inst/HI[425] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[95\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[121\] _384_/Y mprj_logic_high_inst/HI[323] vssd vssd vccd
+ vccd la_oenb_core[121] sky130_fd_sc_hd__einvp_8
XFILLER_1_935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_sel_buf\[2\] _398_/Y mprj_sel_buf\[2\]/TE vssd vssd vccd vccd mprj_sel_o_user[2]
+ sky130_fd_sc_hd__einvp_8
Xinput302 la_oenb_mprj[22] vssd vssd vccd vccd _614_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput335 la_oenb_mprj[52] vssd vssd vccd vccd _644_/A sky130_fd_sc_hd__clkbuf_2
Xinput324 la_oenb_mprj[42] vssd vssd vccd vccd _634_/A sky130_fd_sc_hd__clkbuf_4
Xinput313 la_oenb_mprj[32] vssd vssd vccd vccd _624_/A sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[51\] _643_/Y mprj_logic_high_inst/HI[253] vssd vssd vccd
+ vccd la_oenb_core[51] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[73\] _336_/A la_buf_enable\[73\]/B vssd vssd vccd vccd la_buf\[73\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput357 la_oenb_mprj[72] vssd vssd vccd vccd _335_/A sky130_fd_sc_hd__buf_2
Xinput346 la_oenb_mprj[62] vssd vssd vccd vccd _654_/A sky130_fd_sc_hd__buf_2
Xinput368 la_oenb_mprj[82] vssd vssd vccd vccd _345_/A sky130_fd_sc_hd__clkbuf_4
Xinput379 la_oenb_mprj[92] vssd vssd vccd vccd _355_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input317_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[44\]_A_N _636_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_593_ _593_/A vssd vssd vccd vccd _593_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_16_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[59\] _523_/Y la_buf\[59\]/TE vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_31_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[59\]_A_N _651_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[115\] _579_/Y la_buf\[115\]/TE vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_4_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[57\]_B mprj_logic_high_inst/HI[387] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] user_to_mprj_in_gates\[48\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high_inst/HI[241] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[48\]_B mprj_logic_high_inst/HI[378] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[10\] input143/X mprj_logic_high_inst/HI[340] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[10\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[38\]_A _630_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[99\] _362_/Y mprj_logic_high_inst/HI[301] vssd vssd vccd
+ vccd la_oenb_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input267_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood mprj2_vdd_pwrgood/A vssd vssd vccd vccd output627/A sky130_fd_sc_hd__buf_6
XFILLER_46_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput110 la_data_out_mprj[80] vssd vssd vccd vccd _544_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input434_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput132 la_iena_mprj[0] vssd vssd vccd vccd input132/X sky130_fd_sc_hd__clkbuf_1
Xinput143 la_iena_mprj[10] vssd vssd vccd vccd input143/X sky130_fd_sc_hd__clkbuf_2
Xinput154 la_iena_mprj[11] vssd vssd vccd vccd input154/X sky130_fd_sc_hd__clkbuf_4
Xinput121 la_data_out_mprj[90] vssd vssd vccd vccd _554_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input30_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput165 la_iena_mprj[14] vssd vssd vccd vccd input165/X sky130_fd_sc_hd__clkbuf_1
Xinput176 la_iena_mprj[24] vssd vssd vccd vccd input176/X sky130_fd_sc_hd__clkbuf_1
Xinput187 la_iena_mprj[34] vssd vssd vccd vccd input187/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[39\]_B mprj_logic_high_inst/HI[369] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput198 la_iena_mprj[44] vssd vssd vccd vccd input198/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_645_ _645_/A vssd vssd vccd vccd _645_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_576_ _576_/A vssd vssd vccd vccd _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[29\]_A _621_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd vssd vccd vccd output500/A
+ sky130_fd_sc_hd__inv_2
Xoutput617 output617/A vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_2
Xoutput606 output606/A vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_2
XFILLER_47_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput628 output628/A vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_2
XFILLER_45_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[25\]_A _425_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_A _594_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _416_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[58\] input213/X mprj_logic_high_inst/HI[388] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[58\]/B sky130_fd_sc_hd__and2_1
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _430_/A vssd vssd vccd vccd _430_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_26_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[14\] _606_/Y mprj_logic_high_inst/HI[216] vssd vssd vccd
+ vccd la_oenb_core[14] sky130_fd_sc_hd__einvp_8
X_361_ _361_/A vssd vssd vccd vccd _361_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[36\] _628_/A la_buf_enable\[36\]/B vssd vssd vccd vccd la_buf\[36\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input384_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input78_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_628_ _628_/A vssd vssd vccd vccd _628_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_559_ _559_/A vssd vssd vccd vccd _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput469 output469/A vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_2
XFILLER_47_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__601__A _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__511__A _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input132_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _413_/A vssd vssd vccd vccd _413_/Y sky130_fd_sc_hd__inv_6
XFILLER_53_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _344_/A vssd vssd vccd vccd _344_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[41\] _505_/Y la_buf\[41\]/TE vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__einvp_8
XFILLER_50_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[113\] input147/X mprj_logic_high_inst/HI[443] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[113\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd vssd vccd vccd
+ output484/A sky130_fd_sc_hd__clkinv_4
XFILLER_42_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[29\]_A _461_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output616_A output616/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd vssd vccd vccd output574/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] user_to_mprj_in_gates\[30\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[1\]_A _401_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__331__A _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__506__A _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[81\] _344_/Y mprj_logic_high_inst/HI[283] vssd vssd vccd
+ vccd la_oenb_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input347_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[1\]_B mprj_logic_high_inst/HI[331] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[18\]_A user_wb_dat_gates\[18\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_46_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[89\] _553_/Y la_buf\[89\]/TE vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_21_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[104\] _367_/A la_buf_enable\[104\]/B vssd vssd vccd vccd la_buf\[104\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high_inst/HI[274] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] user_to_mprj_in_gates\[78\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[122\]_B la_buf_enable\[122\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[113\]_B la_buf_enable\[113\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[40\] input194/X mprj_logic_high_inst/HI[370] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[40\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input297_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[4\]_A user_wb_dat_gates\[4\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input60_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[104\]_B la_buf_enable\[104\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd vssd vccd vccd output533/A
+ sky130_fd_sc_hd__inv_2
XFILLER_50_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] user_to_mprj_in_gates\[104\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[88\] input246/X mprj_logic_high_inst/HI[418] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[88\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[114\] _377_/Y mprj_logic_high_inst/HI[316] vssd vssd vccd
+ vccd la_oenb_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_1_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput303 la_oenb_mprj[23] vssd vssd vccd vccd _615_/A sky130_fd_sc_hd__buf_2
Xinput336 la_oenb_mprj[53] vssd vssd vccd vccd _645_/A sky130_fd_sc_hd__buf_2
Xinput325 la_oenb_mprj[43] vssd vssd vccd vccd _635_/A sky130_fd_sc_hd__buf_4
XFILLER_0_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput314 la_oenb_mprj[33] vssd vssd vccd vccd _625_/A sky130_fd_sc_hd__buf_2
XFILLER_40_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput358 la_oenb_mprj[73] vssd vssd vccd vccd _336_/A sky130_fd_sc_hd__clkbuf_4
Xinput347 la_oenb_mprj[63] vssd vssd vccd vccd _655_/A sky130_fd_sc_hd__clkbuf_2
Xinput369 la_oenb_mprj[83] vssd vssd vccd vccd _346_/A sky130_fd_sc_hd__buf_4
Xla_buf_enable\[66\] _329_/A la_buf_enable\[66\]/B vssd vssd vccd vccd la_buf\[66\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[44\] _636_/Y mprj_logic_high_inst/HI[246] vssd vssd vccd
+ vccd la_oenb_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_29_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_irq_buffers\[2\] user_irq_gates\[2\]/Y vssd vssd vccd vccd output630/A sky130_fd_sc_hd__clkinv_4
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_592_ _592_/A vssd vssd vccd vccd _592_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input212_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[108\] _572_/Y la_buf\[108\]/TE vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__einvp_8
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd vssd vccd vccd
+ output465/A sky130_fd_sc_hd__clkinv_4
XFILLER_48_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__604__A _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[0\] _432_/Y mprj_dat_buf\[0\]/TE vssd vssd vccd vccd mprj_dat_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__514__A _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input162_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput100 la_data_out_mprj[71] vssd vssd vccd vccd _535_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput111 la_data_out_mprj[81] vssd vssd vccd vccd _545_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[107\]_TE mprj_logic_high_inst/HI[309] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput122 la_data_out_mprj[91] vssd vssd vccd vccd _555_/A sky130_fd_sc_hd__clkbuf_2
Xinput133 la_iena_mprj[100] vssd vssd vccd vccd input133/X sky130_fd_sc_hd__clkbuf_1
Xinput144 la_iena_mprj[110] vssd vssd vccd vccd input144/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input427_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput166 la_iena_mprj[15] vssd vssd vccd vccd input166/X sky130_fd_sc_hd__clkbuf_1
Xinput177 la_iena_mprj[25] vssd vssd vccd vccd input177/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input23_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput155 la_iena_mprj[120] vssd vssd vccd vccd input155/X sky130_fd_sc_hd__clkbuf_1
X_644_ _644_/A vssd vssd vccd vccd _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput199 la_iena_mprj[45] vssd vssd vccd vccd input199/X sky130_fd_sc_hd__clkbuf_1
Xinput188 la_iena_mprj[35] vssd vssd vccd vccd input188/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[71\] _535_/Y la_buf\[71\]/TE vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__einvp_8
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_575_ _575_/A vssd vssd vccd vccd _575_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xoutput618 output618/A vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_2
Xoutput607 output607/A vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_2
XFILLER_12_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput629 output629/A vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_2
XTAP_147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[90\]_A_N _353_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] user_to_mprj_in_gates\[60\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__334__A _334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_30_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[43\]_A_N _635_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[58\]_A_N _650_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_360_ _360_/A vssd vssd vccd vccd _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[29\] _621_/A la_buf_enable\[29\]/B vssd vssd vccd vccd la_buf\[29\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_42_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input377_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_627_ _627_/A vssd vssd vccd vccd _627_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_53_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_558_ _558_/A vssd vssd vccd vccd _558_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output596_A output596/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_489_ _489_/A vssd vssd vccd vccd _489_/Y sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd vssd vccd vccd output514/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[1\]_B la_buf_enable\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__329__A _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[70\] input227/X mprj_logic_high_inst/HI[400] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[70\]/B sky130_fd_sc_hd__and2_1
XFILLER_47_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input125_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_412_ _412_/A vssd vssd vccd vccd _412_/Y sky130_fd_sc_hd__inv_12
XFILLER_53_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_343_ _343_/A vssd vssd vccd vccd _343_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_42_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[34\] _498_/Y la_buf\[34\]/TE vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__einvp_8
XANTENNA_input90_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[106\] input139/X mprj_logic_high_inst/HI[436] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[106\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd vssd vccd vccd output566/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output609_A output609/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] user_to_mprj_in_gates\[23\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__522__A _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[74\] _337_/Y mprj_logic_high_inst/HI[276] vssd vssd vccd
+ vccd la_oenb_core[74] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[96\] _359_/A la_buf_enable\[96\]/B vssd vssd vccd vccd la_buf\[96\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[22\] _454_/Y mprj_dat_buf\[22\]/TE vssd vssd vccd vccd mprj_dat_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input242_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__432__A _432_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[11\]_A input154/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[2\] _594_/A la_buf_enable\[2\]/B vssd vssd vccd vccd la_buf\[2\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__342__A _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[33\] input186/X mprj_logic_high_inst/HI[363] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[33\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__517__A _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[11\] _603_/A la_buf_enable\[11\]/B vssd vssd vccd vccd la_buf\[11\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input192_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input457_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input53_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] user_to_mprj_in_gates\[90\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__337__A _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high_inst/HI[264] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput326 la_oenb_mprj[44] vssd vssd vccd vccd _636_/A sky130_fd_sc_hd__buf_2
Xinput304 la_oenb_mprj[24] vssd vssd vccd vccd _616_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput315 la_oenb_mprj[34] vssd vssd vccd vccd _626_/A sky130_fd_sc_hd__clkbuf_2
Xuser_to_mprj_oen_buffers\[107\] _370_/Y mprj_logic_high_inst/HI[309] vssd vssd vccd
+ vccd la_oenb_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_40_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput359 la_oenb_mprj[74] vssd vssd vccd vccd _337_/A sky130_fd_sc_hd__buf_2
Xinput348 la_oenb_mprj[64] vssd vssd vccd vccd _656_/A sky130_fd_sc_hd__buf_2
Xinput337 la_oenb_mprj[54] vssd vssd vccd vccd _646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_591_ _591_/A vssd vssd vccd vccd _591_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[59\] _651_/A la_buf_enable\[59\]/B vssd vssd vccd vccd la_buf\[59\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_16_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[37\] _629_/Y mprj_logic_high_inst/HI[239] vssd vssd vccd
+ vccd la_oenb_core[37] sky130_fd_sc_hd__einvp_8
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input205_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd vssd vccd vccd output547/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_1_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[9\]_A _441_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__620__A _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vssd vccd vccd _536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input155_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput112 la_data_out_mprj[82] vssd vssd vccd vccd _546_/A sky130_fd_sc_hd__buf_2
Xinput123 la_data_out_mprj[92] vssd vssd vccd vccd _556_/A sky130_fd_sc_hd__clkbuf_2
Xinput134 la_iena_mprj[101] vssd vssd vccd vccd input134/X sky130_fd_sc_hd__clkbuf_1
Xinput145 la_iena_mprj[111] vssd vssd vccd vccd input145/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input322_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput167 la_iena_mprj[16] vssd vssd vccd vccd input167/X sky130_fd_sc_hd__clkbuf_1
Xinput178 la_iena_mprj[26] vssd vssd vccd vccd input178/X sky130_fd_sc_hd__clkbuf_1
Xinput156 la_iena_mprj[121] vssd vssd vccd vccd input156/X sky130_fd_sc_hd__clkbuf_1
X_643_ _643_/A vssd vssd vccd vccd _643_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput189 la_iena_mprj[36] vssd vssd vccd vccd input189/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input16_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_574_ _574_/A vssd vssd vccd vccd _574_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[64\] _528_/Y la_buf\[64\]/TE vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__einvp_8
XFILLER_17_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_A _589_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[120\] _584_/Y la_buf\[120\]/TE vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[28\] _428_/Y mprj_adr_buf\[28\]/TE vssd vssd vccd vccd mprj_adr_o_user[28]
+ sky130_fd_sc_hd__einvp_8
Xoutput608 output608/A vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_2
XFILLER_49_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[80\]_B la_buf_enable\[80\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput619 output619/A vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_2
XFILLER_45_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__440__A _440_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] user_to_mprj_in_gates\[53\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__615__A _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[116\]_A _580_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[71\]_B la_buf_enable\[71\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__350__A _350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input8_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[12\]_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__525__A _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[62\]_B la_buf_enable\[62\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input272_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[127\] _390_/A la_buf_enable\[127\]/B vssd vssd vccd vccd la_buf\[127\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_626_ _626_/A vssd vssd vccd vccd _626_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_557_ _557_/A vssd vssd vccd vccd _557_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_488_ _488_/A vssd vssd vccd vccd _488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__435__A _435_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd vssd vccd vccd output506/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_B mprj_logic_high_inst/HI[455] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__345__A _345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[63\] input219/X mprj_logic_high_inst/HI[393] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[63\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[116\]_B mprj_logic_high_inst/HI[446] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[41\] _633_/A la_buf_enable\[41\]/B vssd vssd vccd vccd la_buf\[41\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[1\] _593_/Y mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd la_oenb_core[1] sky130_fd_sc_hd__einvp_8
XANTENNA_input118_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_411_ _411_/A vssd vssd vccd vccd _411_/Y sky130_fd_sc_hd__inv_4
XFILLER_42_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ _342_/A vssd vssd vccd vccd _342_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_42_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input83_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[27\] _491_/Y la_buf\[27\]/TE vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__einvp_8
XFILLER_13_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[4\]_A input204/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[107\]_B mprj_logic_high_inst/HI[437] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_609_ _609_/A vssd vssd vccd vccd _609_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[42\]_A_N _634_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[29\]/Y sky130_fd_sc_hd__nand2_2
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] user_to_mprj_in_gates\[16\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[57\]_A_N _649_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[26\] user_wb_dat_gates\[26\]/Y vssd vssd vccd vccd output610/A
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_la_buf_enable\[26\]_B la_buf_enable\[26\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] user_to_mprj_in_gates\[127\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[17\]_B la_buf_enable\[17\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[67\] _330_/Y mprj_logic_high_inst/HI[269] vssd vssd vccd
+ vccd la_oenb_core[67] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[89\] _352_/A la_buf_enable\[89\]/B vssd vssd vccd vccd la_buf\[89\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[96\]_B mprj_logic_high_inst/HI[426] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[15\] _447_/Y mprj_dat_buf\[15\]/TE vssd vssd vccd vccd mprj_dat_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input235_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input402_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[20\]_B mprj_logic_high_inst/HI[350] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[10\] _410_/Y mprj_adr_buf\[10\]/TE vssd vssd vccd vccd mprj_adr_o_user[10]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd vssd vccd vccd
+ output490/A sky130_fd_sc_hd__clkinv_4
XANTENNA_output621_A output621/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[87\]_B mprj_logic_high_inst/HI[417] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd vssd vccd vccd output580/A
+ sky130_fd_sc_hd__inv_2
XFILLER_42_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[0\] user_wb_dat_gates\[0\]/Y vssd vssd vccd vccd output592/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_45_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[11\]_B mprj_logic_high_inst/HI[341] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__623__A _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[4\]_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[26\] input178/X mprj_logic_high_inst/HI[356] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[26\]/B sky130_fd_sc_hd__and2_1
XFILLER_52_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__533__A _533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input352_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input46_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[94\] _558_/Y la_buf\[94\]/TE vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_8_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[59\]_A _651_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__443__A _443_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] user_to_mprj_in_gates\[83\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__353__A _353_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput327 la_oenb_mprj[45] vssd vssd vccd vccd _637_/A sky130_fd_sc_hd__clkbuf_2
Xinput305 la_oenb_mprj[25] vssd vssd vccd vccd _617_/A sky130_fd_sc_hd__buf_2
Xinput316 la_oenb_mprj[35] vssd vssd vccd vccd _627_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput349 la_oenb_mprj[65] vssd vssd vccd vccd _657_/A sky130_fd_sc_hd__clkbuf_2
Xinput338 la_oenb_mprj[55] vssd vssd vccd vccd _647_/A sky130_fd_sc_hd__buf_2
XFILLER_5_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_590_ _590_/A vssd vssd vccd vccd _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input100_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[5\] _469_/Y la_buf\[5\]/TE vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__einvp_8
XFILLER_6_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[2\] _402_/Y mprj_adr_buf\[2\]/TE vssd vssd vccd vccd mprj_adr_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__438__A _438_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd vssd vccd vccd output539/A
+ sky130_fd_sc_hd__inv_2
XFILLER_17_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[10\]_A _442_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[11\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_34_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[28\]_A _428_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__348__A _348_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_A _597_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[93\] input252/X mprj_logic_high_inst/HI[423] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[93\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[19\]_A _419_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_sel_buf\[0\] _396_/Y mprj_sel_buf\[0\]/TE vssd vssd vccd vccd mprj_sel_o_user[0]
+ sky130_fd_sc_hd__einvp_8
Xinput102 la_data_out_mprj[73] vssd vssd vccd vccd _537_/A sky130_fd_sc_hd__buf_2
XFILLER_1_768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput113 la_data_out_mprj[83] vssd vssd vccd vccd _547_/A sky130_fd_sc_hd__clkbuf_4
Xinput124 la_data_out_mprj[93] vssd vssd vccd vccd _557_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput135 la_iena_mprj[102] vssd vssd vccd vccd input135/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input148_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[71\] _334_/A la_buf_enable\[71\]/B vssd vssd vccd vccd la_buf\[71\]/TE
+ sky130_fd_sc_hd__and2b_1
Xinput168 la_iena_mprj[17] vssd vssd vccd vccd input168/X sky130_fd_sc_hd__clkbuf_1
Xinput146 la_iena_mprj[112] vssd vssd vccd vccd input146/X sky130_fd_sc_hd__clkbuf_1
Xinput157 la_iena_mprj[122] vssd vssd vccd vccd input157/X sky130_fd_sc_hd__clkbuf_1
X_642_ _642_/A vssd vssd vccd vccd _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput179 la_iena_mprj[27] vssd vssd vccd vccd input179/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input315_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[30\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_573_ _573_/A vssd vssd vccd vccd _573_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[57\] _521_/Y la_buf\[57\]/TE vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__einvp_8
XFILLER_32_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput609 output609/A vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_2
XFILLER_49_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[113\] _577_/Y la_buf\[113\]/TE vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] user_to_mprj_in_gates\[46\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_23_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] user_to_mprj_in_gates\[8\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[12\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[97\] _360_/Y mprj_logic_high_inst/HI[299] vssd vssd vccd
+ vccd la_oenb_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_5_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__541__A _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input265_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input432_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_625_ _625_/A vssd vssd vccd vccd _625_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_556_ _556_/A vssd vssd vccd vccd _556_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_487_ _487_/A vssd vssd vccd vccd _487_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd vssd vccd vccd output498/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_47_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__451__A _451_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__626__A _626_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_A _404_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__361__A _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[56\] input211/X mprj_logic_high_inst/HI[386] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[56\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _410_/A vssd vssd vccd vccd _410_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_341_ _341_/A vssd vssd vccd vccd _341_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__536__A _536_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[12\] _604_/Y mprj_logic_high_inst/HI[214] vssd vssd vccd
+ vccd la_oenb_core[12] sky130_fd_sc_hd__einvp_8
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[34\] _626_/A la_buf_enable\[34\]/B vssd vssd vccd vccd la_buf\[34\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd vssd vccd vccd output579/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_41_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input382_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input76_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[4\]_B mprj_logic_high_inst/HI[334] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_stb_buf _394_/Y mprj_stb_buf/TE vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__einvp_8
XFILLER_1_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_608_ _608_/A vssd vssd vccd vccd _608_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__446__A _446_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_539_ _539_/A vssd vssd vccd vccd _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[19\] user_wb_dat_gates\[19\]/Y vssd vssd vccd vccd output602/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_29_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[125\]_B la_buf_enable\[125\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__356__A _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[116\]_B la_buf_enable\[116\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input130_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input228_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_buffers\[7\]_A user_wb_dat_gates\[7\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[111\] input145/X mprj_logic_high_inst/HI[441] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[111\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd vssd vccd vccd
+ output482/A sky130_fd_sc_hd__clkinv_4
XFILLER_26_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output614_A output614/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[107\]_B la_buf_enable\[107\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd vssd vccd vccd output572/A
+ sky130_fd_sc_hd__inv_2
XFILLER_0_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[4\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[19\] input170/X mprj_logic_high_inst/HI[349] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[19\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input178_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[41\]_A_N _633_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input345_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input39_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[56\]_A_N _648_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[87\] _551_/Y la_buf\[87\]/TE vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_5_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[102\] _365_/A la_buf_enable\[102\]/B vssd vssd vccd vccd la_buf\[102\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_46_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] user_to_mprj_in_gates\[76\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__634__A _634_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput306 la_oenb_mprj[26] vssd vssd vccd vccd _618_/A sky130_fd_sc_hd__clkbuf_2
Xinput317 la_oenb_mprj[36] vssd vssd vccd vccd _628_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput339 la_oenb_mprj[56] vssd vssd vccd vccd _648_/A sky130_fd_sc_hd__clkbuf_2
Xinput328 la_oenb_mprj[46] vssd vssd vccd vccd _638_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__544__A _544_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input295_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_input462_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_ena_buf\[2\] input462/X user_irq_ena_buf\[2\]/B vssd vssd vccd vccd user_irq_gates\[2\]/B
+ sky130_fd_sc_hd__and2_1
XFILLER_4_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd vssd vccd vccd output531/A
+ sky130_fd_sc_hd__inv_2
XFILLER_34_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__454__A _454_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] user_to_mprj_in_gates\[102\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__364__A _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_33_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[86\] input244/X mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[86\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[112\] _375_/Y mprj_logic_high_inst/HI[314] vssd vssd vccd
+ vccd la_oenb_core[112] sky130_fd_sc_hd__einvp_8
Xinput103 la_data_out_mprj[74] vssd vssd vccd vccd _538_/A sky130_fd_sc_hd__buf_2
Xinput114 la_data_out_mprj[84] vssd vssd vccd vccd _548_/A sky130_fd_sc_hd__buf_4
Xinput125 la_data_out_mprj[94] vssd vssd vccd vccd _558_/A sky130_fd_sc_hd__buf_2
Xinput136 la_iena_mprj[103] vssd vssd vccd vccd input136/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput169 la_iena_mprj[18] vssd vssd vccd vccd input169/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput147 la_iena_mprj[113] vssd vssd vccd vccd input147/X sky130_fd_sc_hd__clkbuf_1
Xinput158 la_iena_mprj[123] vssd vssd vccd vccd input158/X sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[42\] _634_/Y mprj_logic_high_inst/HI[244] vssd vssd vccd
+ vccd la_oenb_core[42] sky130_fd_sc_hd__einvp_8
XANTENNA__539__A _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[64\] _656_/A la_buf_enable\[64\]/B vssd vssd vccd vccd la_buf\[64\]/TE
+ sky130_fd_sc_hd__and2b_1
X_641_ _641_/A vssd vssd vccd vccd _641_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_5_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_buffers\[0\] user_irq_gates\[0\]/Y vssd vssd vccd vccd output628/A sky130_fd_sc_hd__clkinv_4
XFILLER_44_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input210_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_572_ _572_/A vssd vssd vccd vccd _572_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input308_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[106\] _570_/Y la_buf\[106\]/TE vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_45_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__449__A _449_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] user_to_mprj_in_gates\[39\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[4\]_B la_buf_enable\[4\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__359__A _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input258_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input160_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input425_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input21_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_624_ _624_/A vssd vssd vccd vccd _624_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_555_ _555_/A vssd vssd vccd vccd _555_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_486_ _486_/A vssd vssd vccd vccd _486_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_we_buf _395_/Y mprj_we_buf/TE vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__einvp_8
XFILLER_9_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_pwrgood mprj_pwrgood/A vssd vssd vccd vccd output624/A sky130_fd_sc_hd__buf_6
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__642__A _642_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[49\] input203/X mprj_logic_high_inst/HI[379] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[49\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _340_/A vssd vssd vccd vccd _340_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[27\] _619_/A la_buf_enable\[27\]/B vssd vssd vccd vccd la_buf\[27\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__552__A _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input375_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input69_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_607_ _607_/A vssd vssd vccd vccd _607_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_538_ _538_/A vssd vssd vccd vccd _538_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output594_A output594/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_469_ _469_/A vssd vssd vccd vccd _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__462__A _462_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__637__A _637_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__372__A _372_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high_inst/HI[267] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input123_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__A _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[32\] _496_/Y la_buf\[32\]/TE vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__einvp_8
XFILLER_7_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[104\] input137/X mprj_logic_high_inst/HI[434] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[104\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd vssd vccd vccd output564/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output607_A output607/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] user_to_mprj_in_gates\[21\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_buffers\[31\] user_wb_dat_gates\[31\]/Y vssd vssd vccd vccd output616/A
+ sky130_fd_sc_hd__inv_6
Xmprj_dat_buf\[9\] _441_/Y mprj_dat_buf\[9\]/TE vssd vssd vccd vccd mprj_dat_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__367__A _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[72\] _335_/Y mprj_logic_high_inst/HI[274] vssd vssd vccd
+ vccd la_oenb_core[72] sky130_fd_sc_hd__einvp_8
XFILLER_43_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[94\] _357_/A la_buf_enable\[94\]/B vssd vssd vccd vccd la_buf\[94\]/TE
+ sky130_fd_sc_hd__and2b_1
Xoutput590 output590/A vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_2
XFILLER_43_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[20\] _452_/Y mprj_dat_buf\[20\]/TE vssd vssd vccd vccd mprj_dat_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input338_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input240_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] user_to_mprj_in_gates\[69\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_2173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[0\] _592_/A la_buf_enable\[0\]/B vssd vssd vccd vccd la_buf\[0\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__650__A _650_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput318 la_oenb_mprj[37] vssd vssd vccd vccd _629_/A sky130_fd_sc_hd__clkbuf_2
Xinput307 la_oenb_mprj[27] vssd vssd vccd vccd _619_/A sky130_fd_sc_hd__buf_2
XFILLER_44_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput329 la_oenb_mprj[47] vssd vssd vccd vccd _639_/A sky130_fd_sc_hd__buf_4
XFILLER_9_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[31\] input184/X mprj_logic_high_inst/HI[361] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[31\]/B sky130_fd_sc_hd__and2_1
XFILLER_45_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input190_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[92\]_B la_buf_enable\[92\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input288_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input455_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input51_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd vssd vccd vccd output523/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_30_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[83\]_B la_buf_enable\[83\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__470__A _470_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[24\]_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[119\]_A _583_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[40\]_A_N _632_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__645__A _645_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[74\]_B la_buf_enable\[74\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[55\]_A_N _647_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__380__A _380_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[79\] input236/X mprj_logic_high_inst/HI[409] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[79\]/B sky130_fd_sc_hd__and2_1
Xinput104 la_data_out_mprj[75] vssd vssd vccd vccd _539_/A sky130_fd_sc_hd__buf_2
Xinput115 la_data_out_mprj[85] vssd vssd vccd vccd _549_/A sky130_fd_sc_hd__clkbuf_4
Xinput126 la_data_out_mprj[95] vssd vssd vccd vccd _559_/A sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[105\] _368_/Y mprj_logic_high_inst/HI[307] vssd vssd vccd
+ vccd la_oenb_core[105] sky130_fd_sc_hd__einvp_8
Xinput137 la_iena_mprj[104] vssd vssd vccd vccd input137/X sky130_fd_sc_hd__clkbuf_1
Xinput148 la_iena_mprj[114] vssd vssd vccd vccd input148/X sky130_fd_sc_hd__clkbuf_1
Xinput159 la_iena_mprj[124] vssd vssd vccd vccd input159/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_wb_dat_gates\[15\]_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_640_ _640_/A vssd vssd vccd vccd _640_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_5_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_571_ _571_/A vssd vssd vccd vccd _571_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[57\] _649_/A la_buf_enable\[57\]/B vssd vssd vccd vccd la_buf\[57\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[35\] _627_/Y mprj_logic_high_inst/HI[237] vssd vssd vccd
+ vccd la_oenb_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_22_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input203_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__555__A _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input99_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[65\]_B la_buf_enable\[65\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__375__A _375_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[47\]_B la_buf_enable\[47\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input153_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[119\]_B mprj_logic_high_inst/HI[449] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input320_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_623_ _623_/A vssd vssd vccd vccd _623_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_input418_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input14_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[62\] _526_/Y la_buf\[62\]/TE vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_45_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_554_ _554_/A vssd vssd vccd vccd _554_/Y sky130_fd_sc_hd__inv_2
X_485_ _485_/A vssd vssd vccd vccd _485_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[50\]_B mprj_logic_high_inst/HI[380] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[26\] _426_/Y mprj_adr_buf\[26\]/TE vssd vssd vccd vccd mprj_adr_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[7\]_A input237/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] user_to_mprj_in_gates\[51\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[41\]_B mprj_logic_high_inst/HI[371] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_32_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _623_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[32\]_B mprj_logic_high_inst/HI[362] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input368_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input270_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[99\]_B mprj_logic_high_inst/HI[429] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[125\] _388_/A la_buf_enable\[125\]/B vssd vssd vccd vccd la_buf\[125\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_606_ _606_/A vssd vssd vccd vccd _606_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_2_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_537_ _537_/A vssd vssd vccd vccd _537_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[23\]_B mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_468_ _468_/A vssd vssd vccd vccd _468_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_399_ _399_/A vssd vssd vccd vccd _399_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_9_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd vssd vccd vccd output504/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_9_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] user_to_mprj_in_gates\[99\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[14\]_B mprj_logic_high_inst/HI[344] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__653__A _653_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[7\]_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high_inst/HI[312] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[61\] input217/X mprj_logic_high_inst/HI[391] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[61\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_irq_ena_buf\[1\]_B user_irq_ena_buf\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input81_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[25\] _489_/Y la_buf\[25\]/TE vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__einvp_8
XFILLER_6_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd vssd vccd vccd output556/A
+ sky130_fd_sc_hd__inv_2
XFILLER_45_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[27\]/Y sky130_fd_sc_hd__nand2_2
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] user_to_mprj_in_gates\[14\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_31_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[24\] user_wb_dat_gates\[24\]/Y vssd vssd vccd vccd output608/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] user_to_mprj_in_gates\[125\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__648__A _648_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[31\]_A _463_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__383__A _383_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high_inst/HI[234] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput580 output580/A vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[65\] _657_/Y mprj_logic_high_inst/HI[267] vssd vssd vccd
+ vccd la_oenb_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_43_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[87\] _350_/A la_buf_enable\[87\]/B vssd vssd vccd vccd la_buf\[87\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput591 output591/A vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_2
XFILLER_43_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[13\] _445_/Y mprj_dat_buf\[13\]/TE vssd vssd vccd vccd mprj_dat_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input233_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__558__A _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input400_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[22\]_A _454_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd vssd vccd vccd
+ output488/A sky130_fd_sc_hd__clkinv_4
XFILLER_38_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__468__A _468_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_A _445_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput308 la_oenb_mprj[28] vssd vssd vccd vccd _620_/A sky130_fd_sc_hd__clkbuf_4
Xinput319 la_oenb_mprj[38] vssd vssd vccd vccd _630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__378__A _378_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[8\]_A _600_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[11\]_A user_wb_dat_gates\[11\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_12_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[24\] input176/X mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[24\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input183_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input350_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input448_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input44_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[92\] _556_/Y la_buf\[92\]/TE vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_27_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd vssd vccd vccd output625/A sky130_fd_sc_hd__buf_6
XFILLER_21_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] user_to_mprj_in_gates\[81\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_1
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[24\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput105 la_data_out_mprj[76] vssd vssd vccd vccd _540_/A sky130_fd_sc_hd__clkbuf_4
Xinput116 la_data_out_mprj[86] vssd vssd vccd vccd _550_/A sky130_fd_sc_hd__clkbuf_4
Xinput127 la_data_out_mprj[96] vssd vssd vccd vccd _560_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput138 la_iena_mprj[105] vssd vssd vccd vccd input138/X sky130_fd_sc_hd__clkbuf_1
Xinput149 la_iena_mprj[115] vssd vssd vccd vccd input149/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_la_buf_enable\[9\]_A_N _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[15\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_570_ _570_/A vssd vssd vccd vccd _570_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[28\] _620_/Y mprj_logic_high_inst/HI[230] vssd vssd vccd
+ vccd la_oenb_core[28] sky130_fd_sc_hd__einvp_8
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input398_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__571__A _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[3\] _467_/Y la_buf\[3\]/TE vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__einvp_8
XFILLER_10_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[0\] _400_/Y mprj_adr_buf\[0\]/TE vssd vssd vccd vccd mprj_adr_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd vssd vccd vccd output537/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_44_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__481__A _481_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__656__A _656_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[7\]_A _407_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[91\] input250/X mprj_logic_high_inst/HI[421] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[91\]/B sky130_fd_sc_hd__and2_1
XFILLER_46_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input146_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_622_ _622_/A vssd vssd vccd vccd _622_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_24_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input313_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__566__A _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_553_ _553_/A vssd vssd vccd vccd _553_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[55\] _519_/Y la_buf\[55\]/TE vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__einvp_8
XFILLER_44_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_484_ _484_/A vssd vssd vccd vccd _484_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[127\] input162/X mprj_logic_high_inst/HI[457] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[127\]/B sky130_fd_sc_hd__and2_1
XFILLER_18_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[7\]_B mprj_logic_high_inst/HI[337] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[19\] _419_/Y mprj_adr_buf\[19\]/TE vssd vssd vccd vccd mprj_adr_o_user[19]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _575_/Y la_buf\[111\]/TE vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd vssd vccd vccd output589/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_7_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[54\]_A_N _646_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__476__A _476_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[9\] user_wb_dat_gates\[9\]/Y vssd vssd vccd vccd output623/A
+ sky130_fd_sc_hd__clkinv_8
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] user_to_mprj_in_gates\[44\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[69\]_A_N _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] user_to_mprj_in_gates\[6\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__386__A _386_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[95\] _358_/Y mprj_logic_high_inst/HI[297] vssd vssd vccd
+ vccd la_oenb_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_5_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input263_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[119\]_B la_buf_enable\[119\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input430_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[8\] input248/X mprj_logic_high_inst/HI[338] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[8\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[118\] _381_/A la_buf_enable\[118\]/B vssd vssd vccd vccd la_buf\[118\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_605_ _605_/A vssd vssd vccd vccd _605_/Y sky130_fd_sc_hd__clkinv_2
X_536_ _536_/A vssd vssd vccd vccd _536_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_467_ _467_/A vssd vssd vccd vccd _467_/Y sky130_fd_sc_hd__clkinv_2
X_398_ _398_/A vssd vssd vccd vccd _398_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd vssd vccd vccd output496/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_9_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[7\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[54\] input209/X mprj_logic_high_inst/HI[384] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[54\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[10\] _602_/Y mprj_logic_high_inst/HI[212] vssd vssd vccd
+ vccd la_oenb_core[10] sky130_fd_sc_hd__einvp_8
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[32\] _624_/A la_buf_enable\[32\]/B vssd vssd vccd vccd la_buf\[32\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd vssd vccd vccd output557/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_35_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input380_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[18\] _482_/Y la_buf\[18\]/TE vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_6_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input74_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_519_ _519_/A vssd vssd vccd vccd _519_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_21_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[17\] user_wb_dat_gates\[17\]/Y vssd vssd vccd vccd output600/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_25_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] user_to_mprj_in_gates\[118\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput570 output570/A vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_2
Xoutput581 output581/A vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_2
XFILLER_47_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput592 output592/A vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[58\] _650_/Y mprj_logic_high_inst/HI[260] vssd vssd vccd
+ vccd la_oenb_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_8_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input226_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__574__A _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd vssd vccd vccd
+ output480/A sky130_fd_sc_hd__clkinv_4
XFILLER_46_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output612_A output612/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd vssd vccd vccd output570/A
+ sky130_fd_sc_hd__inv_2
XFILLER_37_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_33_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput309 la_oenb_mprj[29] vssd vssd vccd vccd _621_/A sky130_fd_sc_hd__buf_2
XFILLER_44_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__394__A _394_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_24_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[17\] input168/X mprj_logic_high_inst/HI[347] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[17\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input176_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input343_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input37_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[85\] _549_/Y la_buf\[85\]/TE vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_5_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[100\] _363_/A la_buf_enable\[100\]/B vssd vssd vccd vccd la_buf\[100\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] user_to_mprj_in_gates\[74\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_1
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high_inst/HI[224] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[7\]_B la_buf_enable\[7\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__389__A _389_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput106 la_data_out_mprj[77] vssd vssd vccd vccd _541_/A sky130_fd_sc_hd__clkbuf_2
Xinput117 la_data_out_mprj[87] vssd vssd vccd vccd _551_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput128 la_data_out_mprj[97] vssd vssd vccd vccd _561_/A sky130_fd_sc_hd__buf_2
Xinput139 la_iena_mprj[106] vssd vssd vccd vccd input139/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input293_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input460_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[0\] input460/X user_irq_ena_buf\[0\]/B vssd vssd vccd vccd user_irq_gates\[0\]/B
+ sky130_fd_sc_hd__and2_1
XFILLER_10_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd vssd vccd vccd output529/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] user_to_mprj_in_gates\[100\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_2
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[68\]_TE mprj_logic_high_inst/HI[270] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[84\] input242/X mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[84\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[110\] _373_/Y mprj_logic_high_inst/HI[312] vssd vssd vccd
+ vccd la_oenb_core[110] sky130_fd_sc_hd__einvp_8
XFILLER_24_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[40\] _632_/Y mprj_logic_high_inst/HI[242] vssd vssd vccd
+ vccd la_oenb_core[40] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[62\] _654_/A la_buf_enable\[62\]/B vssd vssd vccd vccd la_buf\[62\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_40_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_621_ _621_/A vssd vssd vccd vccd _621_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input139_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_552_ _552_/A vssd vssd vccd vccd _552_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input306_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_483_ _483_/A vssd vssd vccd vccd _483_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[48\] _512_/Y la_buf\[48\]/TE vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_34_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__582__A _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[2\]_A _434_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[104\] _568_/Y la_buf\[104\]/TE vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] user_to_mprj_in_gates\[37\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[88\] _351_/Y mprj_logic_high_inst/HI[290] vssd vssd vccd
+ vccd la_oenb_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_11_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input256_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__577__A _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input423_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_604_ _604_/A vssd vssd vccd vccd _604_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_27_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_535_ _535_/A vssd vssd vccd vccd _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_466_ _466_/A vssd vssd vccd vccd _466_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_43_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_397_ _397_/A vssd vssd vccd vccd _397_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[31\] _431_/Y mprj_adr_buf\[31\]/TE vssd vssd vccd vccd mprj_adr_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__487__A _487_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__397__A _397_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[47\] input201/X mprj_logic_high_inst/HI[377] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[47\]/B sky130_fd_sc_hd__and2_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[25\] _617_/A la_buf_enable\[25\]/B vssd vssd vccd vccd la_buf\[25\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[53\]_A_N _645_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input373_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input67_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[68\]_A_N _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_518_ _518_/A vssd vssd vccd vccd _518_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output592_A output592/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_449_ _449_/A vssd vssd vccd vccd _449_/Y sky130_fd_sc_hd__inv_4
XFILLER_31_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[46\]_A user_to_mprj_in_gates\[46\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput560 output560/A vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_2
Xoutput571 output571/A vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_2
Xoutput582 output582/A vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_2
Xoutput593 output593/A vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_2
XFILLER_8_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input219_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input121_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[100\]_B mprj_logic_high_inst/HI[430] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[95\]_B la_buf_enable\[95\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[30\] _494_/Y la_buf\[30\]/TE vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__einvp_8
XANTENNA__590__A _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[102\] input135/X mprj_logic_high_inst/HI[432] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[102\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[2\]/Y sky130_fd_sc_hd__nand2_8
XFILLER_6_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd vssd vccd vccd
+ output472/A sky130_fd_sc_hd__inv_2
XFILLER_6_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd vssd vccd vccd output562/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_4_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output605_A output605/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_87 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[86\]_B la_buf_enable\[86\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[7\] _439_/Y mprj_dat_buf\[7\]/TE vssd vssd vccd vccd mprj_dat_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[27\]_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[10\]_B la_buf_enable\[10\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[77\]_B la_buf_enable\[77\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input169_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[70\] _333_/Y mprj_logic_high_inst/HI[272] vssd vssd vccd
+ vccd la_oenb_core[70] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[92\] _355_/A la_buf_enable\[92\]/B vssd vssd vccd vccd la_buf\[92\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[18\]_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input336_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[78\] _542_/Y la_buf\[78\]/TE vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__einvp_8
XFILLER_5_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__585__A _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[80\]_B mprj_logic_high_inst/HI[410] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[68\]_B la_buf_enable\[68\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] user_to_mprj_in_gates\[67\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__495__A _495_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput107 la_data_out_mprj[78] vssd vssd vccd vccd _542_/A sky130_fd_sc_hd__buf_2
Xinput118 la_data_out_mprj[88] vssd vssd vccd vccd _552_/A sky130_fd_sc_hd__buf_2
XFILLER_44_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput129 la_data_out_mprj[98] vssd vssd vccd vccd _562_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[62\]_B mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input286_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input453_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[53\]_B mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd vssd vccd vccd output521/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[44\]_B mprj_logic_high_inst/HI[374] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[34\]_A _626_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[77\] input234/X mprj_logic_high_inst/HI[407] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[77\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[103\] _366_/Y mprj_logic_high_inst/HI[305] vssd vssd vccd
+ vccd la_oenb_core[103] sky130_fd_sc_hd__einvp_8
X_620_ _620_/A vssd vssd vccd vccd _620_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_551_ _551_/A vssd vssd vccd vccd _551_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[33\] _625_/Y mprj_logic_high_inst/HI[235] vssd vssd vccd
+ vccd la_oenb_core[33] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[30\]_A _430_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[55\] _647_/A la_buf_enable\[55\]/B vssd vssd vccd vccd la_buf\[55\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[35\]_B mprj_logic_high_inst/HI[365] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_482_ _482_/A vssd vssd vccd vccd _482_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input201_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input97_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput460 user_irq_ena[0] vssd vssd vccd vccd input460/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_A _421_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[26\]_B mprj_logic_high_inst/HI[356] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[16\]_A _608_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[12\]_A _412_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[17\]_B mprj_logic_high_inst/HI[347] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[109\]_A_N _372_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[29\] _461_/Y mprj_dat_buf\[29\]/TE vssd vssd vccd vccd mprj_dat_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input151_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input249_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_603_ _603_/A vssd vssd vccd vccd _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input416_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input12_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[60\] _524_/Y la_buf\[60\]/TE vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__einvp_8
X_534_ _534_/A vssd vssd vccd vccd _534_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__593__A _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_465_ _465_/A vssd vssd vccd vccd _465_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_43_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_396_ _396_/A vssd vssd vccd vccd _396_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_35_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[24\] _424_/Y mprj_adr_buf\[24\]/TE vssd vssd vccd vccd mprj_adr_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput290 la_oenb_mprj[127] vssd vssd vccd vccd _390_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[9\] _601_/A la_buf_enable\[9\]/B vssd vssd vccd vccd la_buf\[9\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input4_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[18\] _610_/A la_buf_enable\[18\]/B vssd vssd vccd vccd la_buf\[18\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_52_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input199_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input366_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[1\] user_irq_core[1] user_irq_gates\[1\]/B vssd vssd vccd vccd user_irq_gates\[1\]/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_46_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__588__A _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[123\] _386_/A la_buf_enable\[123\]/B vssd vssd vccd vccd la_buf\[123\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_A _457_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[7\]_A_N _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_517_ _517_/A vssd vssd vccd vccd _517_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _448_/A vssd vssd vccd vccd _448_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_379_ _379_/A vssd vssd vccd vccd _379_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_35_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] user_to_mprj_in_gates\[97\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__498__A _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput561 output561/A vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_2
Xoutput550 output550/A vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_2
Xoutput572 output572/A vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_2
XFILLER_47_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput583 output583/A vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_2
Xoutput594 output594/A vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_2
XFILLER_47_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_buffers\[14\]_A user_wb_dat_gates\[14\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_1_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input114_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[23\] _487_/Y la_buf\[23\]/TE vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__einvp_8
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd vssd vccd vccd output554/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_45_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[25\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_53_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] user_to_mprj_in_gates\[12\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_53_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_buffers\[22\] user_wb_dat_gates\[22\]/Y vssd vssd vccd vccd output606/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_31_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[27\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] user_to_mprj_in_gates\[123\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[52\]_A_N _644_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[67\]_A_N _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[0\]_A user_wb_dat_gates\[0\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[85\] _348_/A la_buf_enable\[85\]/B vssd vssd vccd vccd la_buf\[85\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[63\] _655_/Y mprj_logic_high_inst/HI[265] vssd vssd vccd
+ vccd la_oenb_core[63] sky130_fd_sc_hd__einvp_8
XFILLER_27_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[18\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[11\] _443_/Y mprj_dat_buf\[11\]/TE vssd vssd vccd vccd mprj_dat_o_user[11]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input231_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input329_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_B la_buf_enable\[100\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[127\] _591_/Y la_buf\[127\]/TE vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__einvp_8
XFILLER_48_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd vssd vccd vccd
+ output486/A sky130_fd_sc_hd__clkinv_4
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput108 la_data_out_mprj[79] vssd vssd vccd vccd _543_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput119 la_data_out_mprj[89] vssd vssd vccd vccd _553_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[22\] input174/X mprj_logic_high_inst/HI[352] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[22\]/B sky130_fd_sc_hd__and2_1
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input181_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input446_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input42_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__596__A _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[90\] _554_/Y la_buf\[90\]/TE vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_35_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput90 la_data_out_mprj[62] vssd vssd vccd vccd _526_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_550_ _550_/A vssd vssd vccd vccd _550_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[48\] _640_/A la_buf_enable\[48\]/B vssd vssd vccd vccd la_buf\[48\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_481_ _481_/A vssd vssd vccd vccd _481_/Y sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_oen_buffers\[8\] _600_/Y mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd la_oenb_core[8] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[26\] _618_/Y mprj_logic_high_inst/HI[228] vssd vssd vccd
+ vccd la_oenb_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_25_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input396_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[1\] _465_/Y la_buf\[1\]/TE vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput461 user_irq_ena[1] vssd vssd vccd vccd input461/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput450 mprj_dat_o_core[7] vssd vssd vccd vccd _439_/A sky130_fd_sc_hd__buf_4
XFILLER_7_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input144_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_602_ _602_/A vssd vssd vccd vccd _602_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input311_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input409_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_533_ _533_/A vssd vssd vccd vccd _533_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_464_ _464_/A vssd vssd vccd vccd _464_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[53\] _517_/Y la_buf\[53\]/TE vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_13_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[125\] input160/X mprj_logic_high_inst/HI[455] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[125\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_395_ _395_/A vssd vssd vccd vccd _395_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[17\] _417_/Y mprj_adr_buf\[17\]/TE vssd vssd vccd vccd mprj_adr_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd vssd vccd vccd output587/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_7_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput280 la_oenb_mprj[118] vssd vssd vccd vccd _381_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xinput291 la_oenb_mprj[12] vssd vssd vccd vccd _604_/A sky130_fd_sc_hd__buf_2
XFILLER_1_1040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] user_to_mprj_in_gates\[42\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[7\] user_wb_dat_gates\[7\]/Y vssd vssd vccd vccd output621/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] user_to_mprj_in_gates\[4\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[93\] _356_/Y mprj_logic_high_inst/HI[295] vssd vssd vccd
+ vccd la_oenb_core[93] sky130_fd_sc_hd__einvp_8
XANTENNA_input261_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input359_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[6\] input226/X mprj_logic_high_inst/HI[336] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[6\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[116\] _379_/A la_buf_enable\[116\]/B vssd vssd vccd vccd la_buf\[116\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_516_ _516_/A vssd vssd vccd vccd _516_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_447_ _447_/A vssd vssd vccd vccd _447_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_378_ _378_/A vssd vssd vccd vccd _378_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_35_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd vssd vccd vccd output494/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_6_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[25\]_TE mprj_logic_high_inst/HI[227] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[108\]_A_N _371_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput562 output562/A vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_2
Xoutput551 output551/A vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_2
Xoutput540 output540/A vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_2
XFILLER_47_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput573 output573/A vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_2
Xoutput584 output584/A vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_2
Xoutput595 output595/A vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_2
XFILLER_25_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[52\] input207/X mprj_logic_high_inst/HI[382] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[52\]/B sky130_fd_sc_hd__and2_1
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[30\] _622_/A la_buf_enable\[30\]/B vssd vssd vccd vccd la_buf\[30\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd vssd vccd vccd output535/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_24_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[16\] _480_/Y la_buf\[16\]/TE vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__einvp_8
XFILLER_32_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input72_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high_inst/HI[250] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__599__A _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[9\] _409_/Y mprj_adr_buf\[9\]/TE vssd vssd vccd vccd mprj_adr_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_43_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[18\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[15\] user_wb_dat_gates\[15\]/Y vssd vssd vccd vccd output598/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] user_to_mprj_in_gates\[116\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[6\]_A_N _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _389_/Y mprj_logic_high_inst/HI[328] vssd vssd vccd
+ vccd la_oenb_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_48_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[56\] _648_/Y mprj_logic_high_inst/HI[258] vssd vssd vccd
+ vccd la_oenb_core[56] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[78\] _341_/A la_buf_enable\[78\]/B vssd vssd vccd vccd la_buf\[78\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_48_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input224_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd vssd vccd vccd
+ output478/A sky130_fd_sc_hd__clkinv_4
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output610_A output610/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput109 la_data_out_mprj[7] vssd vssd vccd vccd _471_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[15\] input166/X mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[15\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input174_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input341_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input439_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input35_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[83\] _547_/Y la_buf\[83\]/TE vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__einvp_8
XFILLER_5_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[5\]_A _437_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[51\]_A_N _643_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] user_to_mprj_in_gates\[72\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_1
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[66\]_A_N _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[19\]_A_N _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput91 la_data_out_mprj[63] vssd vssd vccd vccd _527_/A sky130_fd_sc_hd__clkbuf_2
Xinput80 la_data_out_mprj[53] vssd vssd vccd vccd _517_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_480_ _480_/A vssd vssd vccd vccd _480_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_25_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[19\] _611_/Y mprj_logic_high_inst/HI[221] vssd vssd vccd
+ vccd la_oenb_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_25_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input291_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input389_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[121\]_A _585_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput462 user_irq_ena[2] vssd vssd vccd vccd input462/X sky130_fd_sc_hd__clkbuf_1
Xinput451 mprj_dat_o_core[8] vssd vssd vccd vccd _440_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput440 mprj_dat_o_core[27] vssd vssd vccd vccd _459_/A sky130_fd_sc_hd__buf_2
XANTENNA__400__A _400_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd vssd vccd vccd output527/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[82\] input240/X mprj_logic_high_inst/HI[412] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[82\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[60\] _652_/A la_buf_enable\[60\]/B vssd vssd vccd vccd la_buf\[60\]/TE
+ sky130_fd_sc_hd__and2b_1
X_601_ _601_/A vssd vssd vccd vccd _601_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input137_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_532_ _532_/A vssd vssd vccd vccd _532_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input304_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_463_ _463_/A vssd vssd vccd vccd _463_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_2_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[46\] _510_/Y la_buf\[46\]/TE vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__einvp_8
XFILLER_41_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_394_ _394_/A vssd vssd vccd vccd _394_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[118\] input152/X mprj_logic_high_inst/HI[448] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[118\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[102\] _566_/Y la_buf\[102\]/TE vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_9_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput270 la_oenb_mprj[109] vssd vssd vccd vccd _372_/A sky130_fd_sc_hd__clkbuf_4
Xinput281 la_oenb_mprj[119] vssd vssd vccd vccd _382_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput292 la_oenb_mprj[13] vssd vssd vccd vccd _605_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[121\]_B mprj_logic_high_inst/HI[451] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] user_to_mprj_in_gates\[35\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[40\]_B la_buf_enable\[40\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[89\]_A _553_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[112\]_B mprj_logic_high_inst/HI[442] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[86\] _349_/Y mprj_logic_high_inst/HI[288] vssd vssd vccd
+ vccd la_oenb_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_2_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input254_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[31\]_B la_buf_enable\[31\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input421_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[109\] _372_/A la_buf_enable\[109\]/B vssd vssd vccd vccd la_buf\[109\]/TE
+ sky130_fd_sc_hd__and2b_2
XFILLER_24_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_515_ _515_/A vssd vssd vccd vccd _515_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[103\]_B mprj_logic_high_inst/HI[433] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_446_ _446_/A vssd vssd vccd vccd _446_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[98\]_B la_buf_enable\[98\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_377_ _377_/A vssd vssd vccd vccd _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_B la_buf_enable\[22\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[89\]_B la_buf_enable\[89\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput563 output563/A vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_2
Xoutput552 output552/A vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_2
Xoutput541 output541/A vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_2
Xoutput530 output530/A vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[13\]_B la_buf_enable\[13\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput574 output574/A vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_2
Xoutput585 output585/A vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_2
Xoutput596 output596/A vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_2
XFILLER_25_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[92\]_B mprj_logic_high_inst/HI[422] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[45\] input199/X mprj_logic_high_inst/HI[375] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[45\]/B sky130_fd_sc_hd__and2_1
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[23\] _615_/A la_buf_enable\[23\]/B vssd vssd vccd vccd la_buf\[23\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input371_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input65_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[83\]_B mprj_logic_high_inst/HI[413] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output590_A output590/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ _429_/A vssd vssd vccd vccd _429_/Y sky130_fd_sc_hd__inv_8
XFILLER_37_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[0\]_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput1 caravel_clk vssd vssd vccd vccd _391_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] user_to_mprj_in_gates\[109\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[119\] _382_/Y mprj_logic_high_inst/HI[321] vssd vssd vccd
+ vccd la_oenb_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_0_946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[49\] _641_/Y mprj_logic_high_inst/HI[251] vssd vssd vccd
+ vccd la_oenb_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_19_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input217_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[100\] input133/X mprj_logic_high_inst/HI[430] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[100\]/B sky130_fd_sc_hd__and2_1
XFILLER_7_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[0\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[107\]_A_N _370_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd vssd vccd vccd
+ output470/A sky130_fd_sc_hd__inv_2
XFILLER_43_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd vssd vccd vccd output560/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output603_A output603/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[56\]_B mprj_logic_high_inst/HI[386] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[30\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[5\] _437_/Y mprj_dat_buf\[5\]/TE vssd vssd vccd vccd mprj_dat_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_44_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[47\]_B mprj_logic_high_inst/HI[377] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _629_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input167_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[90\] _353_/A la_buf_enable\[90\]/B vssd vssd vccd vccd la_buf\[90\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_48_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input334_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input28_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[38\]_B mprj_logic_high_inst/HI[368] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[76\] _540_/Y la_buf\[76\]/TE vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_16_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[24\]_A _424_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[29\]_B mprj_logic_high_inst/HI[359] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] user_to_mprj_in_gates\[65\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[5\]_A_N _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _593_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput81 la_data_out_mprj[54] vssd vssd vccd vccd _518_/A sky130_fd_sc_hd__clkbuf_2
Xinput70 la_data_out_mprj[44] vssd vssd vccd vccd _508_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput92 la_data_out_mprj[64] vssd vssd vccd vccd _528_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[15\]_A _415_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input284_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input451_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vssd vccd vccd _450_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput452 mprj_dat_o_core[9] vssd vssd vccd vccd _441_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput441 mprj_dat_o_core[28] vssd vssd vccd vccd _460_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd vssd vccd vccd output519/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[75\] input232/X mprj_logic_high_inst/HI[405] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[75\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _364_/Y mprj_logic_high_inst/HI[303] vssd vssd vccd
+ vccd la_oenb_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_44_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_600_ _600_/A vssd vssd vccd vccd _600_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_27_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_531_ _531_/A vssd vssd vccd vccd _531_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[31\] _623_/Y mprj_logic_high_inst/HI[233] vssd vssd vccd
+ vccd la_oenb_core[31] sky130_fd_sc_hd__einvp_8
XFILLER_2_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[53\] _645_/A la_buf_enable\[53\]/B vssd vssd vccd vccd la_buf\[53\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_33_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_462_ _462_/A vssd vssd vccd vccd _462_/Y sky130_fd_sc_hd__inv_6
XANTENNA_la_buf_enable\[50\]_A_N _642_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_393_ _393_/A vssd vssd vccd vccd _393_/Y sky130_fd_sc_hd__inv_6
XFILLER_13_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[65\]_A_N _657_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input95_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[39\] _503_/Y la_buf\[39\]/TE vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_51_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[28\]_A _460_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput260 la_oenb_mprj[0] vssd vssd vccd vccd _592_/A sky130_fd_sc_hd__clkbuf_2
Xinput271 la_oenb_mprj[10] vssd vssd vccd vccd _602_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput282 la_oenb_mprj[11] vssd vssd vccd vccd _603_/A sky130_fd_sc_hd__clkbuf_2
Xinput293 la_oenb_mprj[14] vssd vssd vccd vccd _606_/A sky130_fd_sc_hd__buf_2
XFILLER_51_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[18\]_A_N _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] user_to_mprj_in_gates\[28\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_2054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[19\]_A _451_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_buffers\[26\]_A user_wb_dat_gates\[26\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_45_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[79\] _342_/Y mprj_logic_high_inst/HI[281] vssd vssd vccd
+ vccd la_oenb_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_2_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[27\] _459_/Y mprj_dat_buf\[27\]/TE vssd vssd vccd vccd mprj_dat_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input247_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[0\]_B mprj_logic_high_inst/HI[330] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input414_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[17\]_A user_wb_dat_gates\[17\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_4_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input10_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_514_ _514_/A vssd vssd vccd vccd _514_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_445_ _445_/A vssd vssd vccd vccd _445_/Y sky130_fd_sc_hd__clkinv_4
X_376_ _376_/A vssd vssd vccd vccd _376_/Y sky130_fd_sc_hd__inv_2
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[22\] _422_/Y mprj_adr_buf\[22\]/TE vssd vssd vccd vccd mprj_adr_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[121\]_B la_buf_enable\[121\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[7\] _599_/A la_buf_enable\[7\]/B vssd vssd vccd vccd la_buf\[7\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput520 output520/A vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_2
Xoutput553 output553/A vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_2
Xoutput542 output542/A vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_2
Xoutput531 output531/A vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_2
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput564 output564/A vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_2
Xoutput575 output575/A vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_2
Xoutput586 output586/A vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_2
Xoutput597 output597/A vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_2
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[112\]_B la_buf_enable\[112\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[38\] input191/X mprj_logic_high_inst/HI[368] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[38\]/B sky130_fd_sc_hd__and2_1
XFILLER_15_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[16\] _608_/A la_buf_enable\[16\]/B vssd vssd vccd vccd la_buf\[16\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input197_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[3\]_A user_wb_dat_gates\[3\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input364_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input58_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[121\] _384_/A la_buf_enable\[121\]/B vssd vssd vccd vccd la_buf\[121\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_4_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[103\]_B la_buf_enable\[103\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ _428_/A vssd vssd vccd vccd _428_/Y sky130_fd_sc_hd__inv_8
XFILLER_50_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_359_ _359_/A vssd vssd vccd vccd _359_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] user_to_mprj_in_gates\[95\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_9_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[0\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput2 caravel_clk2 vssd vssd vccd vccd _392_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input112_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[21\] _485_/Y la_buf\[21\]/TE vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__einvp_8
XFILLER_32_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd vssd vccd vccd output552/A
+ sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_buffers\[4\]_A user_to_mprj_in_gates\[4\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[23\]/Y sky130_fd_sc_hd__nand2_2
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] user_to_mprj_in_gates\[10\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_14_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[20\] user_wb_dat_gates\[20\]/Y vssd vssd vccd vccd output604/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] user_to_mprj_in_gates\[121\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__504__A _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[61\] _653_/Y mprj_logic_high_inst/HI[263] vssd vssd vccd
+ vccd la_oenb_core[61] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[83\] _346_/A la_buf_enable\[83\]/B vssd vssd vccd vccd la_buf\[83\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input327_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[69\] _533_/Y la_buf\[69\]/TE vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__einvp_8
XFILLER_44_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_68 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xla_buf\[125\] _589_/Y la_buf\[125\]/TE vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_10_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] user_to_mprj_in_gates\[58\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput82 la_data_out_mprj[55] vssd vssd vccd vccd _519_/A sky130_fd_sc_hd__clkbuf_2
Xinput71 la_data_out_mprj[45] vssd vssd vccd vccd _509_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput60 la_data_out_mprj[35] vssd vssd vccd vccd _499_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput93 la_data_out_mprj[65] vssd vssd vccd vccd _529_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[20\] input172/X mprj_logic_high_inst/HI[350] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[20\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_A_N _369_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input277_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input40_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input444_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput420 mprj_cyc_o_core vssd vssd vccd vccd _393_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput431 mprj_dat_o_core[19] vssd vssd vccd vccd _451_/A sky130_fd_sc_hd__clkbuf_2
Xinput442 mprj_dat_o_core[29] vssd vssd vccd vccd _461_/A sky130_fd_sc_hd__clkbuf_2
Xinput453 mprj_iena_wb vssd vssd vccd vccd input453/X sky130_fd_sc_hd__buf_2
XFILLER_40_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd vssd vccd vccd output511/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_8_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[0\]_B la_buf_enable\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[68\] input224/X mprj_logic_high_inst/HI[398] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[68\]/B sky130_fd_sc_hd__and2_1
XFILLER_44_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_530_ _530_/A vssd vssd vccd vccd _530_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[46\] _638_/A la_buf_enable\[46\]/B vssd vssd vccd vccd la_buf\[46\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[24\] _616_/Y mprj_logic_high_inst/HI[226] vssd vssd vccd
+ vccd la_oenb_core[24] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[6\] _598_/Y mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd la_oenb_core[6] sky130_fd_sc_hd__einvp_8
XFILLER_32_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_461_ _461_/A vssd vssd vccd vccd _461_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_392_ _392_/A vssd vssd vccd vccd _392_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input394_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input88_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[4\]_A_N _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput250 la_iena_mprj[91] vssd vssd vccd vccd input250/X sky130_fd_sc_hd__clkbuf_1
Xinput261 la_oenb_mprj[100] vssd vssd vccd vccd _363_/A sky130_fd_sc_hd__clkbuf_4
Xinput272 la_oenb_mprj[110] vssd vssd vccd vccd _373_/A sky130_fd_sc_hd__clkbuf_4
Xinput294 la_oenb_mprj[15] vssd vssd vccd vccd _607_/A sky130_fd_sc_hd__clkbuf_2
Xinput283 la_oenb_mprj[120] vssd vssd vccd vccd _383_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__602__A _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__512__A _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input142_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input407_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_513_ _513_/A vssd vssd vccd vccd _513_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_444_ _444_/A vssd vssd vccd vccd _444_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[51\] _515_/Y la_buf\[51\]/TE vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__einvp_8
X_375_ _375_/A vssd vssd vccd vccd _375_/Y sky130_fd_sc_hd__inv_2
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[123\] input158/X mprj_logic_high_inst/HI[453] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[123\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[15\] _415_/Y mprj_adr_buf\[15\]/TE vssd vssd vccd vccd mprj_adr_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output626_A output626/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd vssd vccd vccd output585/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] user_to_mprj_in_gates\[40\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[5\] user_wb_dat_gates\[5\]/Y vssd vssd vccd vccd output619/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_52_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_A input143/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__332__A _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput510 output510/A vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_2
Xoutput554 output554/A vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_2
Xoutput543 output543/A vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_2
Xoutput532 output532/A vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_2
Xoutput521 output521/A vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_2
Xoutput565 output565/A vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_2
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] user_to_mprj_in_gates\[2\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_1
Xoutput576 output576/A vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_2
Xoutput587 output587/A vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_2
XFILLER_8_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput598 output598/A vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_2
XFILLER_46_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[64\]_A_N _656_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[79\]_A_N _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__507__A _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[91\] _354_/Y mprj_logic_high_inst/HI[293] vssd vssd vccd
+ vccd la_oenb_core[91] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[17\]_A_N _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input357_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[99\] _563_/Y la_buf\[99\]/TE vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_4_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[4\] input204/X mprj_logic_high_inst/HI[334] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[4\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[114\] _377_/A la_buf_enable\[114\]/B vssd vssd vccd vccd la_buf\[114\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_46_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_427_ _427_/A vssd vssd vccd vccd _427_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_14_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_358_ _358_/A vssd vssd vccd vccd _358_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd vssd vccd vccd output474/A
+ sky130_fd_sc_hd__inv_6
XFILLER_6_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] user_to_mprj_in_gates\[88\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput3 caravel_rstn vssd vssd vccd vccd input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[50\] input205/X mprj_logic_high_inst/HI[380] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[50\]/B sky130_fd_sc_hd__and2_1
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd vssd vccd vccd output513/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[14\] _478_/Y la_buf\[14\]/TE vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__einvp_8
XANTENNA_input70_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[61\]_TE mprj_logic_high_inst/HI[263] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[7\] _407_/Y mprj_adr_buf\[7\]/TE vssd vssd vccd vccd mprj_adr_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd vssd vccd vccd output544/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[8\]_A _440_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[16\]/Y sky130_fd_sc_hd__nand2_8
XFILLER_50_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[13\] user_wb_dat_gates\[13\]/Y vssd vssd vccd vccd output596/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__610__A _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] user_to_mprj_in_gates\[114\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[98\] input257/X mprj_logic_high_inst/HI[428] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[98\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[124\] _387_/Y mprj_logic_high_inst/HI[326] vssd vssd vccd
+ vccd la_oenb_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_43_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__520__A _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[54\] _646_/Y mprj_logic_high_inst/HI[256] vssd vssd vccd
+ vccd la_oenb_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_0_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[76\] _339_/A la_buf_enable\[76\]/B vssd vssd vccd vccd la_buf\[76\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input222_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[118\] _582_/Y la_buf\[118\]/TE vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_3_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd vssd vccd vccd
+ output476/A sky130_fd_sc_hd__clkinv_4
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__605__A _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput72 la_data_out_mprj[46] vssd vssd vccd vccd _510_/A sky130_fd_sc_hd__clkbuf_2
Xinput50 la_data_out_mprj[26] vssd vssd vccd vccd _490_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 la_data_out_mprj[36] vssd vssd vccd vccd _500_/A sky130_fd_sc_hd__clkbuf_1
Xinput94 la_data_out_mprj[66] vssd vssd vccd vccd _530_/A sky130_fd_sc_hd__clkbuf_2
Xinput83 la_data_out_mprj[56] vssd vssd vccd vccd _520_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_B la_buf_enable\[70\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__340__A _340_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[11\]_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[13\] input164/X mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[13\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__515__A _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input172_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput421 mprj_dat_o_core[0] vssd vssd vccd vccd _432_/A sky130_fd_sc_hd__clkbuf_8
Xinput410 mprj_adr_o_core[2] vssd vssd vccd vccd _402_/A sky130_fd_sc_hd__buf_12
XFILLER_7_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input437_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input33_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput454 mprj_sel_o_core[0] vssd vssd vccd vccd _396_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput432 mprj_dat_o_core[1] vssd vssd vccd vccd _433_/A sky130_fd_sc_hd__clkbuf_4
Xinput443 mprj_dat_o_core[2] vssd vssd vccd vccd _434_/A sky130_fd_sc_hd__buf_4
XFILLER_48_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[81\] _545_/Y la_buf\[81\]/TE vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_5_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] user_to_mprj_in_gates\[70\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_1
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[124\]_B mprj_logic_high_inst/HI[454] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _391_/Y mprj_clk_buf/TE vssd vssd vccd vccd user_clock sky130_fd_sc_hd__einvp_8
XFILLER_22_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__335__A _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[43\]_B la_buf_enable\[43\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[115\]_B mprj_logic_high_inst/HI[445] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_460_ _460_/A vssd vssd vccd vccd _460_/Y sky130_fd_sc_hd__clkinv_4
Xuser_to_mprj_oen_buffers\[17\] _609_/Y mprj_logic_high_inst/HI[219] vssd vssd vccd
+ vccd la_oenb_core[17] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[39\] _631_/A la_buf_enable\[39\]/B vssd vssd vccd vccd la_buf\[39\]/TE
+ sky130_fd_sc_hd__and2b_1
X_391_ _391_/A vssd vssd vccd vccd _391_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_40_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input387_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[3\]_A input193/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput240 la_iena_mprj[82] vssd vssd vccd vccd input240/X sky130_fd_sc_hd__clkbuf_1
Xinput251 la_iena_mprj[92] vssd vssd vccd vccd input251/X sky130_fd_sc_hd__clkbuf_1
Xinput262 la_oenb_mprj[101] vssd vssd vccd vccd _364_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput295 la_oenb_mprj[16] vssd vssd vccd vccd _608_/A sky130_fd_sc_hd__clkbuf_2
Xinput273 la_oenb_mprj[111] vssd vssd vccd vccd _374_/A sky130_fd_sc_hd__buf_4
Xinput284 la_oenb_mprj[121] vssd vssd vccd vccd _384_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_ena_buf\[106\]_B mprj_logic_high_inst/HI[436] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_589_ _589_/A vssd vssd vccd vccd _589_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd vssd vccd vccd output525/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_53_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[25\]_B la_buf_enable\[25\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[105\]_A_N _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[16\]_B la_buf_enable\[16\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[80\] input238/X mprj_logic_high_inst/HI[410] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[80\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[95\]_B mprj_logic_high_inst/HI[425] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input135_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ _512_/A vssd vssd vccd vccd _512_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input302_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_443_ _443_/A vssd vssd vccd vccd _443_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_374_ _374_/A vssd vssd vccd vccd _374_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[44\] _508_/Y la_buf\[44\]/TE vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_13_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[116\] input150/X mprj_logic_high_inst/HI[446] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[116\]/B sky130_fd_sc_hd__and2_1
XFILLER_29_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[100\] _564_/Y la_buf\[100\]/TE vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_9_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output619_A output619/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[86\]_B mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd vssd vccd vccd output577/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] user_to_mprj_in_gates\[33\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_B mprj_logic_high_inst/HI[340] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__613__A _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput500 output500/A vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_2
Xoutput511 output511/A vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_2
XFILLER_47_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput544 output544/A vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_2
Xoutput533 output533/A vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_2
Xoutput522 output522/A vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_2
XANTENNA_user_wb_dat_gates\[3\]_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput566 output566/A vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_2
Xoutput555 output555/A vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_2
Xoutput577 output577/A vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_2
Xoutput588 output588/A vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_2
Xoutput599 output599/A vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_2
XFILLER_45_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[3\]_A_N _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__523__A _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[84\] _347_/Y mprj_logic_high_inst/HI[286] vssd vssd vccd
+ vccd la_oenb_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_2_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input252_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[107\] _370_/A la_buf_enable\[107\]/B vssd vssd vccd vccd la_buf\[107\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_426_ _426_/A vssd vssd vccd vccd _426_/Y sky130_fd_sc_hd__inv_12
XFILLER_53_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_357_ _357_/A vssd vssd vccd vccd _357_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__433__A _433_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[59\]_B mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput4 la_data_out_mprj[0] vssd vssd vccd vccd _464_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__608__A _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__343__A _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[43\] input197/X mprj_logic_high_inst/HI[373] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[43\]/B sky130_fd_sc_hd__and2_1
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__518__A _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[21\] _613_/A la_buf_enable\[21\]/B vssd vssd vccd vccd la_buf\[21\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_23_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input63_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_ack_buffer user_wb_ack_gate/Y vssd vssd vccd vccd output591/A sky130_fd_sc_hd__clkinv_8
XFILLER_19_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_409_ _409_/A vssd vssd vccd vccd _409_/Y sky130_fd_sc_hd__inv_8
XFILLER_14_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[63\]_A_N _655_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[78\]_A_N _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[27\]_A _427_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] user_to_mprj_in_gates\[107\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__338__A _338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[16\]_A_N _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _596_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[18\]_A _418_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[117\] _380_/Y mprj_logic_high_inst/HI[319] vssd vssd vccd
+ vccd la_oenb_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_7_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[47\] _639_/Y mprj_logic_high_inst/HI[249] vssd vssd vccd
+ vccd la_oenb_core[47] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[69\] _332_/A la_buf_enable\[69\]/B vssd vssd vccd vccd la_buf\[69\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input215_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd vssd vccd vccd
+ output468/A sky130_fd_sc_hd__inv_2
XFILLER_43_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd vssd vccd vccd output558/A
+ sky130_fd_sc_hd__inv_2
XANTENNA_output601_A output601/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[20\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput40 la_data_out_mprj[17] vssd vssd vccd vccd _481_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput73 la_data_out_mprj[47] vssd vssd vccd vccd _511_/A sky130_fd_sc_hd__clkbuf_2
Xinput62 la_data_out_mprj[37] vssd vssd vccd vccd _501_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 la_data_out_mprj[27] vssd vssd vccd vccd _491_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__621__A _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput95 la_data_out_mprj[67] vssd vssd vccd vccd _531_/A sky130_fd_sc_hd__clkbuf_2
Xinput84 la_data_out_mprj[57] vssd vssd vccd vccd _521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[3\] _435_/Y mprj_dat_buf\[3\]/TE vssd vssd vccd vccd mprj_dat_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[11\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__531__A _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input165_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput400 mprj_adr_o_core[20] vssd vssd vccd vccd _420_/A sky130_fd_sc_hd__clkbuf_2
Xinput411 mprj_adr_o_core[30] vssd vssd vccd vccd _430_/A sky130_fd_sc_hd__buf_2
XFILLER_48_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input332_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput455 mprj_sel_o_core[1] vssd vssd vccd vccd _397_/A sky130_fd_sc_hd__clkbuf_2
Xinput422 mprj_dat_o_core[10] vssd vssd vccd vccd _442_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput433 mprj_dat_o_core[20] vssd vssd vccd vccd _452_/A sky130_fd_sc_hd__clkbuf_2
Xinput444 mprj_dat_o_core[30] vssd vssd vccd vccd _462_/A sky130_fd_sc_hd__buf_2
XFILLER_48_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input26_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[74\] _538_/Y la_buf\[74\]/TE vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__einvp_8
XFILLER_32_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__441__A _441_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] user_to_mprj_in_gates\[63\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__616__A _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_A _403_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__351__A _351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_390_ _390_/A vssd vssd vccd vccd _390_/Y sky130_fd_sc_hd__inv_2
XANTENNA__526__A _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input282_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[3\]_B mprj_logic_high_inst/HI[333] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput230 la_iena_mprj[73] vssd vssd vccd vccd input230/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput241 la_iena_mprj[83] vssd vssd vccd vccd input241/X sky130_fd_sc_hd__clkbuf_1
Xinput252 la_iena_mprj[93] vssd vssd vccd vccd input252/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput263 la_oenb_mprj[102] vssd vssd vccd vccd _365_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xinput296 la_oenb_mprj[17] vssd vssd vccd vccd _609_/A sky130_fd_sc_hd__buf_2
Xinput274 la_oenb_mprj[112] vssd vssd vccd vccd _375_/A sky130_fd_sc_hd__buf_2
Xinput285 la_oenb_mprj[122] vssd vssd vccd vccd _385_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_657_ _657_/A vssd vssd vccd vccd _657_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_588_ _588_/A vssd vssd vccd vccd _588_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__436__A _436_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd vssd vccd vccd output517/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[124\]_B la_buf_enable\[124\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__346__A _346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[73\] input230/X mprj_logic_high_inst/HI[403] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[73\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[115\]_B la_buf_enable\[115\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input128_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ _511_/A vssd vssd vccd vccd _511_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[51\] _643_/A la_buf_enable\[51\]/B vssd vssd vccd vccd la_buf\[51\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _442_/A vssd vssd vccd vccd _442_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_373_ _373_/A vssd vssd vccd vccd _373_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_wb_dat_buffers\[6\]_A user_wb_dat_gates\[6\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input93_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[37\] _501_/Y la_buf\[37\]/TE vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[109\] input142/X mprj_logic_high_inst/HI[439] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[109\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_B la_buf_enable\[106\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] user_to_mprj_in_gates\[26\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput501 output501/A vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_2
Xoutput545 output545/A vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_2
Xoutput534 output534/A vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_2
Xoutput523 output523/A vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_2
Xoutput512 output512/A vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_2
XANTENNA_user_wb_dat_gates\[3\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput556 output556/A vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_2
XFILLER_5_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput567 output567/A vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_2
Xoutput578 output578/A vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_2
XFILLER_47_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput589 output589/A vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_2
XFILLER_41_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[77\] _340_/Y mprj_logic_high_inst/HI[279] vssd vssd vccd
+ vccd la_oenb_core[77] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[99\] _362_/A la_buf_enable\[99\]/B vssd vssd vccd vccd la_buf\[99\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[25\] _457_/Y mprj_dat_buf\[25\]/TE vssd vssd vccd vccd mprj_dat_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input245_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_17 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input412_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_425_ _425_/A vssd vssd vccd vccd _425_/Y sky130_fd_sc_hd__inv_12
XANTENNA_la_buf_enable\[104\]_A_N _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_356_ _356_/A vssd vssd vccd vccd _356_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[20\] _420_/Y mprj_adr_buf\[20\]/TE vssd vssd vccd vccd mprj_adr_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[119\]_A_N _382_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput5 la_data_out_mprj[100] vssd vssd vccd vccd _564_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__624__A _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[5\] _597_/A la_buf_enable\[5\]/B vssd vssd vccd vccd la_buf\[5\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[36\] input189/X mprj_logic_high_inst/HI[366] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[36\]/B sky130_fd_sc_hd__and2_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__534__A _534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[14\] _606_/A la_buf_enable\[14\]/B vssd vssd vccd vccd la_buf\[14\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input195_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input362_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input56_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _408_/A vssd vssd vccd vccd _408_/Y sky130_fd_sc_hd__clkinv_16
XFILLER_14_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__444__A _444_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_15_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_339_ _339_/A vssd vssd vccd vccd _339_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] user_to_mprj_in_gates\[93\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[2\]_A_N _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__619__A _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__354__A _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__529__A _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input208_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__439__A _439_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd vssd vccd vccd output550/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[21\]/Y sky130_fd_sc_hd__nand2_2
Xinput30 la_data_out_mprj[123] vssd vssd vccd vccd _587_/A sky130_fd_sc_hd__buf_2
XFILLER_15_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput63 la_data_out_mprj[38] vssd vssd vccd vccd _502_/A sky130_fd_sc_hd__clkbuf_1
Xinput41 la_data_out_mprj[18] vssd vssd vccd vccd _482_/A sky130_fd_sc_hd__clkbuf_2
Xinput52 la_data_out_mprj[28] vssd vssd vccd vccd _492_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_la_buf_enable\[3\]_B la_buf_enable\[3\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput96 la_data_out_mprj[68] vssd vssd vccd vccd _532_/A sky130_fd_sc_hd__clkbuf_2
Xinput85 la_data_out_mprj[58] vssd vssd vccd vccd _522_/A sky130_fd_sc_hd__clkbuf_2
Xinput74 la_data_out_mprj[48] vssd vssd vccd vccd _512_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__349__A _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[81\] _344_/A la_buf_enable\[81\]/B vssd vssd vccd vccd la_buf\[81\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input158_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput401 mprj_adr_o_core[21] vssd vssd vccd vccd _421_/A sky130_fd_sc_hd__buf_2
Xinput412 mprj_adr_o_core[31] vssd vssd vccd vccd _431_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput423 mprj_dat_o_core[11] vssd vssd vccd vccd _443_/A sky130_fd_sc_hd__clkbuf_4
Xinput434 mprj_dat_o_core[21] vssd vssd vccd vccd _453_/A sky130_fd_sc_hd__clkbuf_2
Xinput445 mprj_dat_o_core[31] vssd vssd vccd vccd _463_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input325_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput456 mprj_sel_o_core[2] vssd vssd vccd vccd _398_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_la_buf_enable\[62\]_A_N _654_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input19_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[67\] _531_/Y la_buf\[67\]/TE vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[77\]_A_N _340_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[123\] _587_/Y la_buf\[123\]/TE vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__einvp_8
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] user_to_mprj_in_gates\[56\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__632__A _632_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__542__A _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input442_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_iena_mprj[64] vssd vssd vccd vccd input220/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput231 la_iena_mprj[74] vssd vssd vccd vccd input231/X sky130_fd_sc_hd__clkbuf_1
Xinput242 la_iena_mprj[84] vssd vssd vccd vccd input242/X sky130_fd_sc_hd__clkbuf_1
Xinput253 la_iena_mprj[94] vssd vssd vccd vccd input253/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput297 la_oenb_mprj[18] vssd vssd vccd vccd _610_/A sky130_fd_sc_hd__clkbuf_2
Xinput264 la_oenb_mprj[103] vssd vssd vccd vccd _366_/A sky130_fd_sc_hd__clkbuf_4
Xinput275 la_oenb_mprj[113] vssd vssd vccd vccd _376_/A sky130_fd_sc_hd__clkbuf_4
Xinput286 la_oenb_mprj[123] vssd vssd vccd vccd _386_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_656_ _656_/A vssd vssd vccd vccd _656_/Y sky130_fd_sc_hd__inv_2
X_587_ _587_/A vssd vssd vccd vccd _587_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output494_A output494/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd vssd vccd vccd output509/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__362__A _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[66\] input222/X mprj_logic_high_inst/HI[396] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[66\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_510_ _510_/A vssd vssd vccd vccd _510_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[4\] _596_/Y mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd la_oenb_core[4] sky130_fd_sc_hd__einvp_8
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__537__A _537_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[22\] _614_/Y mprj_logic_high_inst/HI[224] vssd vssd vccd
+ vccd la_oenb_core[22] sky130_fd_sc_hd__einvp_8
X_441_ _441_/A vssd vssd vccd vccd _441_/Y sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[44\] _636_/A la_buf_enable\[44\]/B vssd vssd vccd vccd la_buf\[44\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _372_/A vssd vssd vccd vccd _372_/Y sky130_fd_sc_hd__inv_2
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input392_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input86_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_639_ _639_/A vssd vssd vccd vccd _639_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__447__A _447_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] user_to_mprj_in_gates\[19\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_53_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput502 output502/A vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_2
Xuser_wb_dat_buffers\[29\] user_wb_dat_gates\[29\]/Y vssd vssd vccd vccd output613/A
+ sky130_fd_sc_hd__clkinv_8
Xoutput535 output535/A vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_2
Xoutput524 output524/A vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_2
Xoutput513 output513/A vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_2
XFILLER_47_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput568 output568/A vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_2
Xoutput557 output557/A vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_2
Xoutput546 output546/A vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_2
XFILLER_5_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput579 output579/A vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_2
XFILLER_8_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__A _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[18\] _450_/Y mprj_dat_buf\[18\]/TE vssd vssd vccd vccd mprj_dat_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input238_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input140_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input405_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_424_ _424_/A vssd vssd vccd vccd _424_/Y sky130_fd_sc_hd__clkinv_16
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_355_ _355_/A vssd vssd vccd vccd _355_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_31_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[121\] input156/X mprj_logic_high_inst/HI[451] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[121\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[91\]_A _555_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[13\] _413_/Y mprj_adr_buf\[13\]/TE vssd vssd vccd vccd mprj_adr_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd vssd vccd vccd
+ output493/A sky130_fd_sc_hd__clkinv_4
XFILLER_46_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd vssd vccd vccd output583/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output624_A output624/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput6 la_data_out_mprj[101] vssd vssd vccd vccd _565_/A sky130_fd_sc_hd__clkbuf_4
Xuser_wb_dat_buffers\[3\] user_wb_dat_gates\[3\]/Y vssd vssd vccd vccd output617/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_51_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__640__A _640_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] user_to_mprj_in_gates\[0\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[29\] input181/X mprj_logic_high_inst/HI[359] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[29\]/B sky130_fd_sc_hd__and2_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input188_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[91\]_B la_buf_enable\[91\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__550__A _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input355_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input49_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[112\] _375_/A la_buf_enable\[112\]/B vssd vssd vccd vccd la_buf\[112\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_43_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[97\] _561_/Y la_buf\[97\]/TE vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[2\] input182/X mprj_logic_high_inst/HI[332] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[2\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_407_ _407_/A vssd vssd vccd vccd _407_/Y sky130_fd_sc_hd__inv_8
X_338_ _338_/A vssd vssd vccd vccd _338_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_B la_buf_enable\[82\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] user_to_mprj_in_gates\[86\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[23\]_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__635__A _635_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_B la_buf_enable\[73\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__370__A _370_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[103\]_A_N _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[14\]_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[118\]_A_N _381_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input103_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__545__A _545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd vssd vccd vccd output463/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_36_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[64\]_B la_buf_enable\[64\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[12\] _476_/Y la_buf\[12\]/TE vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__einvp_8
Xla_buf\[8\] _472_/Y la_buf\[8\]/TE vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__einvp_8
XFILLER_49_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[5\] _405_/Y mprj_adr_buf\[5\]/TE vssd vssd vccd vccd mprj_adr_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_43_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd vssd vccd vccd output542/A
+ sky130_fd_sc_hd__inv_2
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__455__A _455_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[14\]/Y sky130_fd_sc_hd__nand2_4
Xinput20 la_data_out_mprj[114] vssd vssd vccd vccd _578_/A sky130_fd_sc_hd__clkbuf_1
Xinput31 la_data_out_mprj[124] vssd vssd vccd vccd _588_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput64 la_data_out_mprj[39] vssd vssd vccd vccd _503_/A sky130_fd_sc_hd__clkbuf_1
Xinput42 la_data_out_mprj[19] vssd vssd vccd vccd _483_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 la_data_out_mprj[29] vssd vssd vccd vccd _493_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput97 la_data_out_mprj[69] vssd vssd vccd vccd _533_/A sky130_fd_sc_hd__clkbuf_2
Xinput86 la_data_out_mprj[59] vssd vssd vccd vccd _523_/A sky130_fd_sc_hd__clkbuf_2
Xinput75 la_data_out_mprj[49] vssd vssd vccd vccd _513_/A sky130_fd_sc_hd__clkbuf_2
Xuser_wb_dat_buffers\[11\] user_wb_dat_gates\[11\]/Y vssd vssd vccd vccd output594/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[127\]_B mprj_logic_high_inst/HI[457] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] user_to_mprj_in_gates\[112\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__365__A _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[28\]_A _492_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[96\] input255/X mprj_logic_high_inst/HI[426] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[96\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[122\] _385_/Y mprj_logic_high_inst/HI[324] vssd vssd vccd
+ vccd la_oenb_core[122] sky130_fd_sc_hd__einvp_8
XFILLER_27_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[3\] _399_/Y mprj_sel_buf\[3\]/TE vssd vssd vccd vccd mprj_sel_o_user[3]
+ sky130_fd_sc_hd__einvp_8
Xinput402 mprj_adr_o_core[22] vssd vssd vccd vccd _422_/A sky130_fd_sc_hd__clkbuf_2
Xuser_to_mprj_oen_buffers\[52\] _644_/Y mprj_logic_high_inst/HI[254] vssd vssd vccd
+ vccd la_oenb_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput413 mprj_adr_o_core[3] vssd vssd vccd vccd _403_/A sky130_fd_sc_hd__buf_2
Xinput446 mprj_dat_o_core[3] vssd vssd vccd vccd _435_/A sky130_fd_sc_hd__buf_2
Xinput424 mprj_dat_o_core[12] vssd vssd vccd vccd _444_/A sky130_fd_sc_hd__clkbuf_4
Xinput435 mprj_dat_o_core[22] vssd vssd vccd vccd _454_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[118\]_B mprj_logic_high_inst/HI[448] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[74\] _337_/A la_buf_enable\[74\]/B vssd vssd vccd vccd la_buf\[74\]/TE
+ sky130_fd_sc_hd__and2b_1
Xinput457 mprj_sel_o_core[3] vssd vssd vccd vccd _399_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input220_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input318_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[1\]_A_N _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[116\] _580_/Y la_buf\[116\]/TE vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_4_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[6\]_A input226/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk2_buf_A _392_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[109\]_B mprj_logic_high_inst/HI[439] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] user_to_mprj_in_gates\[49\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[40\]_B mprj_logic_high_inst/HI[370] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_A _622_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[11\] input154/X mprj_logic_high_inst/HI[341] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[11\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_B mprj_logic_high_inst/HI[361] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[19\]_B la_buf_enable\[19\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input170_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input268_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[98\]_B mprj_logic_high_inst/HI[428] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput210 la_iena_mprj[55] vssd vssd vccd vccd input210/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input435_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput232 la_iena_mprj[75] vssd vssd vccd vccd input232/X sky130_fd_sc_hd__clkbuf_1
Xinput221 la_iena_mprj[65] vssd vssd vccd vccd input221/X sky130_fd_sc_hd__clkbuf_1
Xinput243 la_iena_mprj[85] vssd vssd vccd vccd input243/X sky130_fd_sc_hd__clkbuf_1
Xinput254 la_iena_mprj[95] vssd vssd vccd vccd input254/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input31_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput265 la_oenb_mprj[104] vssd vssd vccd vccd _367_/A sky130_fd_sc_hd__buf_2
Xinput276 la_oenb_mprj[114] vssd vssd vccd vccd _377_/A sky130_fd_sc_hd__clkbuf_4
Xinput287 la_oenb_mprj[124] vssd vssd vccd vccd _387_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput298 la_oenb_mprj[19] vssd vssd vccd vccd _611_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_655_ _655_/A vssd vssd vccd vccd _655_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_586_ _586_/A vssd vssd vccd vccd _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[22\]_B mprj_logic_high_inst/HI[352] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd vssd vccd vccd output501/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_32_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _604_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[89\]_B mprj_logic_high_inst/HI[419] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[13\]_B mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__643__A _643_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[6\]_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[61\]_A_N _653_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[76\]_A_N _339_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[59\] input214/X mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[59\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[0\]_B user_irq_ena_buf\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ _440_/A vssd vssd vccd vccd _440_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ _371_/A vssd vssd vccd vccd _371_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[15\] _607_/Y mprj_logic_high_inst/HI[217] vssd vssd vccd
+ vccd la_oenb_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_14_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[37\] _629_/A la_buf_enable\[37\]/B vssd vssd vccd vccd la_buf\[37\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[14\]_A_N _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input385_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[29\]_A_N _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input79_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_638_ _638_/A vssd vssd vccd vccd _638_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_569_ _569_/A vssd vssd vccd vccd _569_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__463__A _463_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput536 output536/A vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_2
Xoutput525 output525/A vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_2
Xoutput503 output503/A vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_2
Xoutput514 output514/A vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_2
Xoutput558 output558/A vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_2
Xoutput547 output547/A vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_2
Xoutput569 output569/A vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_2
XFILLER_47_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__638__A _638_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_A _462_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__373__A _373_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input133_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__548__A _548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input300_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_423_ _423_/A vssd vssd vccd vccd _423_/Y sky130_fd_sc_hd__inv_8
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[21\]_A _453_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[42\] _506_/Y la_buf\[42\]/TE vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__einvp_8
X_354_ _354_/A vssd vssd vccd vccd _354_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[114\] input148/X mprj_logic_high_inst/HI[444] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[114\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high_inst/HI[233] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output617_A output617/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd vssd vccd vccd output575/A
+ sky130_fd_sc_hd__clkinv_4
Xinput7 la_data_out_mprj[102] vssd vssd vccd vccd _566_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] user_to_mprj_in_gates\[31\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_37 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__368__A _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[7\]_A _599_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_buffers\[10\]_A user_wb_dat_gates\[10\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[82\] _345_/Y mprj_logic_high_inst/HI[284] vssd vssd vccd
+ vccd la_oenb_core[82] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[30\] _462_/Y mprj_dat_buf\[30\]/TE vssd vssd vccd vccd mprj_dat_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input348_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input250_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[105\] _368_/A la_buf_enable\[105\]/B vssd vssd vccd vccd la_buf\[105\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_406_ _406_/A vssd vssd vccd vccd _406_/Y sky130_fd_sc_hd__clkinv_8
X_337_ _337_/A vssd vssd vccd vccd _337_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_41_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] user_to_mprj_in_gates\[79\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[23\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__651__A _651_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[41\] input195/X mprj_logic_high_inst/HI[371] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[41\]/B sky130_fd_sc_hd__and2_1
XFILLER_44_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input298_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__561__A _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd vssd vccd vccd output534/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_50_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 la_data_out_mprj[105] vssd vssd vccd vccd _569_/A sky130_fd_sc_hd__clkbuf_1
Xinput21 la_data_out_mprj[115] vssd vssd vccd vccd _579_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__471__A _471_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput54 la_data_out_mprj[2] vssd vssd vccd vccd _466_/A sky130_fd_sc_hd__clkbuf_2
Xinput43 la_data_out_mprj[1] vssd vssd vccd vccd _465_/A sky130_fd_sc_hd__clkbuf_2
Xinput32 la_data_out_mprj[125] vssd vssd vccd vccd _589_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput98 la_data_out_mprj[6] vssd vssd vccd vccd _470_/A sky130_fd_sc_hd__clkbuf_2
Xinput87 la_data_out_mprj[5] vssd vssd vccd vccd _469_/A sky130_fd_sc_hd__clkbuf_2
Xinput76 la_data_out_mprj[4] vssd vssd vccd vccd _468_/A sky130_fd_sc_hd__clkbuf_2
Xinput65 la_data_out_mprj[3] vssd vssd vccd vccd _467_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] user_to_mprj_in_gates\[105\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__646__A _646_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2_uq6 vssd2_uq5 mprj2_logic_high
XANTENNA_mprj_adr_buf\[6\]_A _406_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__A _381_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[89\] input247/X mprj_logic_high_inst/HI[419] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[89\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[115\] _378_/Y mprj_logic_high_inst/HI[317] vssd vssd vccd
+ vccd la_oenb_core[115] sky130_fd_sc_hd__einvp_8
Xinput403 mprj_adr_o_core[23] vssd vssd vccd vccd _423_/A sky130_fd_sc_hd__clkbuf_2
Xinput414 mprj_adr_o_core[4] vssd vssd vccd vccd _404_/A sky130_fd_sc_hd__buf_12
Xinput425 mprj_dat_o_core[13] vssd vssd vccd vccd _445_/A sky130_fd_sc_hd__clkbuf_4
Xinput436 mprj_dat_o_core[23] vssd vssd vccd vccd _455_/A sky130_fd_sc_hd__buf_2
Xinput458 mprj_stb_o_core vssd vssd vccd vccd _394_/A sky130_fd_sc_hd__buf_4
Xinput447 mprj_dat_o_core[4] vssd vssd vccd vccd _436_/A sky130_fd_sc_hd__buf_4
Xuser_to_mprj_oen_buffers\[45\] _637_/Y mprj_logic_high_inst/HI[247] vssd vssd vccd
+ vccd la_oenb_core[45] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[67\] _330_/A la_buf_enable\[67\]/B vssd vssd vccd vccd la_buf\[67\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_1207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input213_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__556__A _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[6\]_B mprj_logic_high_inst/HI[336] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[109\] _573_/Y la_buf\[109\]/TE vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__einvp_8
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd vssd vccd vccd
+ output466/A sky130_fd_sc_hd__inv_2
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__466__A _466_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[102\]_A_N _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_A_N _380_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[127\]_B la_buf_enable\[127\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[1\] _433_/Y mprj_dat_buf\[1\]/TE vssd vssd vccd vccd mprj_dat_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf_enable\[26\]/B la_buf_enable\[27\]/B
+ la_buf_enable\[28\]/B la_buf_enable\[29\]/B la_buf_enable\[30\]/B la_buf_enable\[31\]/B
+ la_buf_enable\[32\]/B la_buf_enable\[33\]/B la_buf_enable\[34\]/B la_buf_enable\[35\]/B
+ mprj_adr_buf\[0\]/TE la_buf_enable\[36\]/B la_buf_enable\[37\]/B la_buf_enable\[38\]/B
+ la_buf_enable\[39\]/B la_buf_enable\[40\]/B la_buf_enable\[41\]/B la_buf_enable\[42\]/B
+ la_buf_enable\[43\]/B la_buf_enable\[44\]/B la_buf_enable\[45\]/B mprj_adr_buf\[1\]/TE
+ la_buf_enable\[46\]/B la_buf_enable\[47\]/B la_buf_enable\[48\]/B la_buf_enable\[49\]/B
+ la_buf_enable\[50\]/B la_buf_enable\[51\]/B la_buf_enable\[52\]/B la_buf_enable\[53\]/B
+ la_buf_enable\[54\]/B la_buf_enable\[55\]/B mprj_adr_buf\[2\]/TE la_buf_enable\[56\]/B
+ la_buf_enable\[57\]/B la_buf_enable\[58\]/B la_buf_enable\[59\]/B la_buf_enable\[60\]/B
+ la_buf_enable\[61\]/B la_buf_enable\[62\]/B la_buf_enable\[63\]/B la_buf_enable\[64\]/B
+ la_buf_enable\[65\]/B mprj_adr_buf\[3\]/TE la_buf_enable\[66\]/B la_buf_enable\[67\]/B
+ la_buf_enable\[68\]/B la_buf_enable\[69\]/B la_buf_enable\[70\]/B la_buf_enable\[71\]/B
+ la_buf_enable\[72\]/B la_buf_enable\[73\]/B la_buf_enable\[74\]/B la_buf_enable\[75\]/B
+ mprj_adr_buf\[4\]/TE la_buf_enable\[76\]/B la_buf_enable\[77\]/B la_buf_enable\[78\]/B
+ la_buf_enable\[79\]/B la_buf_enable\[80\]/B la_buf_enable\[81\]/B la_buf_enable\[82\]/B
+ la_buf_enable\[83\]/B la_buf_enable\[84\]/B la_buf_enable\[85\]/B mprj_adr_buf\[5\]/TE
+ la_buf_enable\[86\]/B la_buf_enable\[87\]/B la_buf_enable\[88\]/B la_buf_enable\[89\]/B
+ la_buf_enable\[90\]/B la_buf_enable\[91\]/B la_buf_enable\[92\]/B la_buf_enable\[93\]/B
+ la_buf_enable\[94\]/B la_buf_enable\[95\]/B mprj_adr_buf\[6\]/TE la_buf_enable\[96\]/B
+ la_buf_enable\[97\]/B la_buf_enable\[98\]/B la_buf_enable\[99\]/B la_buf_enable\[100\]/B
+ la_buf_enable\[101\]/B la_buf_enable\[102\]/B la_buf_enable\[103\]/B la_buf_enable\[104\]/B
+ la_buf_enable\[105\]/B mprj_adr_buf\[7\]/TE la_buf_enable\[106\]/B la_buf_enable\[107\]/B
+ la_buf_enable\[108\]/B la_buf_enable\[109\]/B la_buf_enable\[110\]/B la_buf_enable\[111\]/B
+ la_buf_enable\[112\]/B la_buf_enable\[113\]/B la_buf_enable\[114\]/B la_buf_enable\[115\]/B
+ mprj_adr_buf\[8\]/TE la_buf_enable\[116\]/B la_buf_enable\[117\]/B la_buf_enable\[118\]/B
+ la_buf_enable\[119\]/B la_buf_enable\[120\]/B la_buf_enable\[121\]/B la_buf_enable\[122\]/B
+ la_buf_enable\[123\]/B la_buf_enable\[124\]/B la_buf_enable\[125\]/B mprj_adr_buf\[9\]/TE
+ mprj_clk_buf/TE la_buf_enable\[126\]/B la_buf_enable\[127\]/B mprj_logic_high_inst/HI[202]
+ mprj_logic_high_inst/HI[203] mprj_logic_high_inst/HI[204] mprj_logic_high_inst/HI[205]
+ mprj_logic_high_inst/HI[206] mprj_logic_high_inst/HI[207] mprj_logic_high_inst/HI[208]
+ mprj_logic_high_inst/HI[209] mprj_adr_buf\[10\]/TE mprj_logic_high_inst/HI[210]
+ mprj_logic_high_inst/HI[211] mprj_logic_high_inst/HI[212] mprj_logic_high_inst/HI[213]
+ mprj_logic_high_inst/HI[214] mprj_logic_high_inst/HI[215] mprj_logic_high_inst/HI[216]
+ mprj_logic_high_inst/HI[217] mprj_logic_high_inst/HI[218] mprj_logic_high_inst/HI[219]
+ mprj_adr_buf\[11\]/TE mprj_logic_high_inst/HI[220] mprj_logic_high_inst/HI[221]
+ mprj_logic_high_inst/HI[222] mprj_logic_high_inst/HI[223] mprj_logic_high_inst/HI[224]
+ mprj_logic_high_inst/HI[225] mprj_logic_high_inst/HI[226] mprj_logic_high_inst/HI[227]
+ mprj_logic_high_inst/HI[228] mprj_logic_high_inst/HI[229] mprj_adr_buf\[12\]/TE
+ mprj_logic_high_inst/HI[230] mprj_logic_high_inst/HI[231] mprj_logic_high_inst/HI[232]
+ mprj_logic_high_inst/HI[233] mprj_logic_high_inst/HI[234] mprj_logic_high_inst/HI[235]
+ mprj_logic_high_inst/HI[236] mprj_logic_high_inst/HI[237] mprj_logic_high_inst/HI[238]
+ mprj_logic_high_inst/HI[239] mprj_adr_buf\[13\]/TE mprj_logic_high_inst/HI[240]
+ mprj_logic_high_inst/HI[241] mprj_logic_high_inst/HI[242] mprj_logic_high_inst/HI[243]
+ mprj_logic_high_inst/HI[244] mprj_logic_high_inst/HI[245] mprj_logic_high_inst/HI[246]
+ mprj_logic_high_inst/HI[247] mprj_logic_high_inst/HI[248] mprj_logic_high_inst/HI[249]
+ mprj_adr_buf\[14\]/TE mprj_logic_high_inst/HI[250] mprj_logic_high_inst/HI[251]
+ mprj_logic_high_inst/HI[252] mprj_logic_high_inst/HI[253] mprj_logic_high_inst/HI[254]
+ mprj_logic_high_inst/HI[255] mprj_logic_high_inst/HI[256] mprj_logic_high_inst/HI[257]
+ mprj_logic_high_inst/HI[258] mprj_logic_high_inst/HI[259] mprj_adr_buf\[15\]/TE
+ mprj_logic_high_inst/HI[260] mprj_logic_high_inst/HI[261] mprj_logic_high_inst/HI[262]
+ mprj_logic_high_inst/HI[263] mprj_logic_high_inst/HI[264] mprj_logic_high_inst/HI[265]
+ mprj_logic_high_inst/HI[266] mprj_logic_high_inst/HI[267] mprj_logic_high_inst/HI[268]
+ mprj_logic_high_inst/HI[269] mprj_adr_buf\[16\]/TE mprj_logic_high_inst/HI[270]
+ mprj_logic_high_inst/HI[271] mprj_logic_high_inst/HI[272] mprj_logic_high_inst/HI[273]
+ mprj_logic_high_inst/HI[274] mprj_logic_high_inst/HI[275] mprj_logic_high_inst/HI[276]
+ mprj_logic_high_inst/HI[277] mprj_logic_high_inst/HI[278] mprj_logic_high_inst/HI[279]
+ mprj_adr_buf\[17\]/TE mprj_logic_high_inst/HI[280] mprj_logic_high_inst/HI[281]
+ mprj_logic_high_inst/HI[282] mprj_logic_high_inst/HI[283] mprj_logic_high_inst/HI[284]
+ mprj_logic_high_inst/HI[285] mprj_logic_high_inst/HI[286] mprj_logic_high_inst/HI[287]
+ mprj_logic_high_inst/HI[288] mprj_logic_high_inst/HI[289] mprj_adr_buf\[18\]/TE
+ mprj_logic_high_inst/HI[290] mprj_logic_high_inst/HI[291] mprj_logic_high_inst/HI[292]
+ mprj_logic_high_inst/HI[293] mprj_logic_high_inst/HI[294] mprj_logic_high_inst/HI[295]
+ mprj_logic_high_inst/HI[296] mprj_logic_high_inst/HI[297] mprj_logic_high_inst/HI[298]
+ mprj_logic_high_inst/HI[299] mprj_adr_buf\[19\]/TE mprj_clk2_buf/TE mprj_logic_high_inst/HI[300]
+ mprj_logic_high_inst/HI[301] mprj_logic_high_inst/HI[302] mprj_logic_high_inst/HI[303]
+ mprj_logic_high_inst/HI[304] mprj_logic_high_inst/HI[305] mprj_logic_high_inst/HI[306]
+ mprj_logic_high_inst/HI[307] mprj_logic_high_inst/HI[308] mprj_logic_high_inst/HI[309]
+ mprj_adr_buf\[20\]/TE mprj_logic_high_inst/HI[310] mprj_logic_high_inst/HI[311]
+ mprj_logic_high_inst/HI[312] mprj_logic_high_inst/HI[313] mprj_logic_high_inst/HI[314]
+ mprj_logic_high_inst/HI[315] mprj_logic_high_inst/HI[316] mprj_logic_high_inst/HI[317]
+ mprj_logic_high_inst/HI[318] mprj_logic_high_inst/HI[319] mprj_adr_buf\[21\]/TE
+ mprj_logic_high_inst/HI[320] mprj_logic_high_inst/HI[321] mprj_logic_high_inst/HI[322]
+ mprj_logic_high_inst/HI[323] mprj_logic_high_inst/HI[324] mprj_logic_high_inst/HI[325]
+ mprj_logic_high_inst/HI[326] mprj_logic_high_inst/HI[327] mprj_logic_high_inst/HI[328]
+ mprj_logic_high_inst/HI[329] mprj_adr_buf\[22\]/TE mprj_logic_high_inst/HI[330]
+ mprj_logic_high_inst/HI[331] mprj_logic_high_inst/HI[332] mprj_logic_high_inst/HI[333]
+ mprj_logic_high_inst/HI[334] mprj_logic_high_inst/HI[335] mprj_logic_high_inst/HI[336]
+ mprj_logic_high_inst/HI[337] mprj_logic_high_inst/HI[338] mprj_logic_high_inst/HI[339]
+ mprj_adr_buf\[23\]/TE mprj_logic_high_inst/HI[340] mprj_logic_high_inst/HI[341]
+ mprj_logic_high_inst/HI[342] mprj_logic_high_inst/HI[343] mprj_logic_high_inst/HI[344]
+ mprj_logic_high_inst/HI[345] mprj_logic_high_inst/HI[346] mprj_logic_high_inst/HI[347]
+ mprj_logic_high_inst/HI[348] mprj_logic_high_inst/HI[349] mprj_adr_buf\[24\]/TE
+ mprj_logic_high_inst/HI[350] mprj_logic_high_inst/HI[351] mprj_logic_high_inst/HI[352]
+ mprj_logic_high_inst/HI[353] mprj_logic_high_inst/HI[354] mprj_logic_high_inst/HI[355]
+ mprj_logic_high_inst/HI[356] mprj_logic_high_inst/HI[357] mprj_logic_high_inst/HI[358]
+ mprj_logic_high_inst/HI[359] mprj_adr_buf\[25\]/TE mprj_logic_high_inst/HI[360]
+ mprj_logic_high_inst/HI[361] mprj_logic_high_inst/HI[362] mprj_logic_high_inst/HI[363]
+ mprj_logic_high_inst/HI[364] mprj_logic_high_inst/HI[365] mprj_logic_high_inst/HI[366]
+ mprj_logic_high_inst/HI[367] mprj_logic_high_inst/HI[368] mprj_logic_high_inst/HI[369]
+ mprj_adr_buf\[26\]/TE mprj_logic_high_inst/HI[370] mprj_logic_high_inst/HI[371]
+ mprj_logic_high_inst/HI[372] mprj_logic_high_inst/HI[373] mprj_logic_high_inst/HI[374]
+ mprj_logic_high_inst/HI[375] mprj_logic_high_inst/HI[376] mprj_logic_high_inst/HI[377]
+ mprj_logic_high_inst/HI[378] mprj_logic_high_inst/HI[379] mprj_adr_buf\[27\]/TE
+ mprj_logic_high_inst/HI[380] mprj_logic_high_inst/HI[381] mprj_logic_high_inst/HI[382]
+ mprj_logic_high_inst/HI[383] mprj_logic_high_inst/HI[384] mprj_logic_high_inst/HI[385]
+ mprj_logic_high_inst/HI[386] mprj_logic_high_inst/HI[387] mprj_logic_high_inst/HI[388]
+ mprj_logic_high_inst/HI[389] mprj_adr_buf\[28\]/TE mprj_logic_high_inst/HI[390]
+ mprj_logic_high_inst/HI[391] mprj_logic_high_inst/HI[392] mprj_logic_high_inst/HI[393]
+ mprj_logic_high_inst/HI[394] mprj_logic_high_inst/HI[395] mprj_logic_high_inst/HI[396]
+ mprj_logic_high_inst/HI[397] mprj_logic_high_inst/HI[398] mprj_logic_high_inst/HI[399]
+ mprj_adr_buf\[29\]/TE mprj_cyc_buf/TE mprj_logic_high_inst/HI[400] mprj_logic_high_inst/HI[401]
+ mprj_logic_high_inst/HI[402] mprj_logic_high_inst/HI[403] mprj_logic_high_inst/HI[404]
+ mprj_logic_high_inst/HI[405] mprj_logic_high_inst/HI[406] mprj_logic_high_inst/HI[407]
+ mprj_logic_high_inst/HI[408] mprj_logic_high_inst/HI[409] mprj_adr_buf\[30\]/TE
+ mprj_logic_high_inst/HI[410] mprj_logic_high_inst/HI[411] mprj_logic_high_inst/HI[412]
+ mprj_logic_high_inst/HI[413] mprj_logic_high_inst/HI[414] mprj_logic_high_inst/HI[415]
+ mprj_logic_high_inst/HI[416] mprj_logic_high_inst/HI[417] mprj_logic_high_inst/HI[418]
+ mprj_logic_high_inst/HI[419] mprj_adr_buf\[31\]/TE mprj_logic_high_inst/HI[420]
+ mprj_logic_high_inst/HI[421] mprj_logic_high_inst/HI[422] mprj_logic_high_inst/HI[423]
+ mprj_logic_high_inst/HI[424] mprj_logic_high_inst/HI[425] mprj_logic_high_inst/HI[426]
+ mprj_logic_high_inst/HI[427] mprj_logic_high_inst/HI[428] mprj_logic_high_inst/HI[429]
+ mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430] mprj_logic_high_inst/HI[431] mprj_logic_high_inst/HI[432]
+ mprj_logic_high_inst/HI[433] mprj_logic_high_inst/HI[434] mprj_logic_high_inst/HI[435]
+ mprj_logic_high_inst/HI[436] mprj_logic_high_inst/HI[437] mprj_logic_high_inst/HI[438]
+ mprj_logic_high_inst/HI[439] mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440] mprj_logic_high_inst/HI[441]
+ mprj_logic_high_inst/HI[442] mprj_logic_high_inst/HI[443] mprj_logic_high_inst/HI[444]
+ mprj_logic_high_inst/HI[445] mprj_logic_high_inst/HI[446] mprj_logic_high_inst/HI[447]
+ mprj_logic_high_inst/HI[448] mprj_logic_high_inst/HI[449] mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450]
+ mprj_logic_high_inst/HI[451] mprj_logic_high_inst/HI[452] mprj_logic_high_inst/HI[453]
+ mprj_logic_high_inst/HI[454] mprj_logic_high_inst/HI[455] mprj_logic_high_inst/HI[456]
+ mprj_logic_high_inst/HI[457] user_irq_ena_buf\[0\]/B user_irq_ena_buf\[1\]/B mprj_dat_buf\[3\]/TE
+ user_irq_ena_buf\[2\]/B mprj_pwrgood/A user_to_mprj_wb_ena_buf/B mprj_dat_buf\[4\]/TE
+ mprj_dat_buf\[5\]/TE mprj_dat_buf\[6\]/TE mprj_dat_buf\[7\]/TE mprj_stb_buf/TE mprj_dat_buf\[8\]/TE
+ mprj_dat_buf\[9\]/TE mprj_dat_buf\[10\]/TE mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE
+ mprj_dat_buf\[13\]/TE mprj_dat_buf\[14\]/TE mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE
+ mprj_dat_buf\[17\]/TE mprj_we_buf/TE mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE
+ mprj_dat_buf\[20\]/TE mprj_dat_buf\[21\]/TE mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE
+ mprj_dat_buf\[24\]/TE mprj_dat_buf\[25\]/TE mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE
+ mprj_sel_buf\[0\]/TE mprj_dat_buf\[28\]/TE mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE
+ mprj_dat_buf\[31\]/TE la_buf_enable\[0\]/B la_buf_enable\[1\]/B la_buf_enable\[2\]/B
+ la_buf_enable\[3\]/B la_buf_enable\[4\]/B la_buf_enable\[5\]/B mprj_sel_buf\[1\]/TE
+ la_buf_enable\[6\]/B la_buf_enable\[7\]/B la_buf_enable\[8\]/B la_buf_enable\[9\]/B
+ la_buf_enable\[10\]/B la_buf_enable\[11\]/B la_buf_enable\[12\]/B la_buf_enable\[13\]/B
+ la_buf_enable\[14\]/B la_buf_enable\[15\]/B mprj_sel_buf\[2\]/TE la_buf_enable\[16\]/B
+ la_buf_enable\[17\]/B la_buf_enable\[18\]/B la_buf_enable\[19\]/B la_buf_enable\[20\]/B
+ la_buf_enable\[21\]/B la_buf_enable\[22\]/B la_buf_enable\[23\]/B la_buf_enable\[24\]/B
+ la_buf_enable\[25\]/B mprj_sel_buf\[3\]/TE vccd1_uq5 vssd1_uq4 mprj_logic_high
XFILLER_26_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__376__A _376_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input163_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[118\]_B la_buf_enable\[118\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput211 la_iena_mprj[56] vssd vssd vccd vccd input211/X sky130_fd_sc_hd__clkbuf_1
Xinput200 la_iena_mprj[46] vssd vssd vccd vccd input200/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput233 la_iena_mprj[76] vssd vssd vccd vccd input233/X sky130_fd_sc_hd__clkbuf_1
Xinput222 la_iena_mprj[66] vssd vssd vccd vccd input222/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input330_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput244 la_iena_mprj[86] vssd vssd vccd vccd input244/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input428_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput255 la_iena_mprj[96] vssd vssd vccd vccd input255/X sky130_fd_sc_hd__clkbuf_1
Xinput266 la_oenb_mprj[105] vssd vssd vccd vccd _368_/A sky130_fd_sc_hd__buf_4
Xinput277 la_oenb_mprj[115] vssd vssd vccd vccd _378_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input24_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput288 la_oenb_mprj[125] vssd vssd vccd vccd _388_/A sky130_fd_sc_hd__clkbuf_4
X_654_ _654_/A vssd vssd vccd vccd _654_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput299 la_oenb_mprj[1] vssd vssd vccd vccd _593_/A sky130_fd_sc_hd__buf_2
XFILLER_5_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[72\] _536_/Y la_buf\[72\]/TE vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__einvp_8
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_585_ _585_/A vssd vssd vccd vccd _585_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[9\]_A user_wb_dat_gates\[9\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[109\]_B la_buf_enable\[109\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] user_to_mprj_in_gates\[61\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[6\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[0\]_A_N _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_370_ _370_/A vssd vssd vccd vccd _370_/Y sky130_fd_sc_hd__inv_2
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input280_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input378_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_637_ _637_/A vssd vssd vccd vccd _637_/Y sky130_fd_sc_hd__inv_2
X_568_ _568_/A vssd vssd vccd vccd _568_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output597_A output597/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd vssd vccd vccd output515/A
+ sky130_fd_sc_hd__clkinv_4
X_499_ _499_/A vssd vssd vccd vccd _499_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput526 output526/A vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_2
Xoutput504 output504/A vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_2
Xoutput515 output515/A vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_2
Xoutput559 output559/A vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_2
Xoutput548 output548/A vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_2
Xoutput537 output537/A vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_2
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__654__A _654_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[71\] input228/X mprj_logic_high_inst/HI[401] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[71\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input126_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_422_ _422_/A vssd vssd vccd vccd _422_/Y sky130_fd_sc_hd__inv_6
XFILLER_14_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__564__A _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/A vssd vssd vccd vccd _353_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input91_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[35\] _499_/Y la_buf\[35\]/TE vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_10_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[107\] input140/X mprj_logic_high_inst/HI[437] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[107\]/B sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[7\]/Y sky130_fd_sc_hd__nand2_8
XFILLER_10_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput8 la_data_out_mprj[103] vssd vssd vccd vccd _567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd vssd vccd vccd output567/A
+ sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[60\]_A_N _652_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__474__A _474_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_36_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] user_to_mprj_in_gates\[24\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[75\]_A_N _338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_A_N _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__649__A _649_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_A_N _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__384__A _384_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[75\] _338_/Y mprj_logic_high_inst/HI[277] vssd vssd vccd
+ vccd la_oenb_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_3_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[97\] _360_/A la_buf_enable\[97\]/B vssd vssd vccd vccd la_buf\[97\]/TE
+ sky130_fd_sc_hd__and2b_2
XFILLER_47_1892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[23\] _455_/Y mprj_dat_buf\[23\]/TE vssd vssd vccd vccd mprj_dat_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input243_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__559__A _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input410_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_405_ _405_/A vssd vssd vccd vccd _405_/Y sky130_fd_sc_hd__inv_16
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _336_/A vssd vssd vccd vccd _336_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__469__A _469_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[6\]_B la_buf_enable\[6\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[3\] _595_/A la_buf_enable\[3\]/B vssd vssd vccd vccd la_buf\[3\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_21_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__379__A _379_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high_inst/HI[223] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[34\] input187/X mprj_logic_high_inst/HI[364] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[34\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[12\] _604_/A la_buf_enable\[12\]/B vssd vssd vccd vccd la_buf\[12\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input193_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input360_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input458_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input54_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xpowergood_check mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A vccd vssd vccd vssd vccd vssd
+ mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput11 la_data_out_mprj[106] vssd vssd vccd vccd _570_/A sky130_fd_sc_hd__buf_2
Xinput22 la_data_out_mprj[116] vssd vssd vccd vccd _580_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput44 la_data_out_mprj[20] vssd vssd vccd vccd _484_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 la_data_out_mprj[30] vssd vssd vccd vccd _494_/A sky130_fd_sc_hd__clkbuf_2
Xinput33 la_data_out_mprj[126] vssd vssd vccd vccd _590_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput88 la_data_out_mprj[60] vssd vssd vccd vccd _524_/A sky130_fd_sc_hd__clkbuf_2
Xinput77 la_data_out_mprj[50] vssd vssd vccd vccd _514_/A sky130_fd_sc_hd__clkbuf_2
Xinput66 la_data_out_mprj[40] vssd vssd vccd vccd _504_/A sky130_fd_sc_hd__clkbuf_2
Xinput99 la_data_out_mprj[70] vssd vssd vccd vccd _534_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] user_to_mprj_in_gates\[91\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[43\]_A input197/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput415 mprj_adr_o_core[5] vssd vssd vccd vccd _405_/A sky130_fd_sc_hd__clkbuf_4
Xinput426 mprj_dat_o_core[14] vssd vssd vccd vccd _446_/A sky130_fd_sc_hd__buf_4
Xinput404 mprj_adr_o_core[24] vssd vssd vccd vccd _424_/A sky130_fd_sc_hd__buf_4
Xinput437 mprj_dat_o_core[24] vssd vssd vccd vccd _456_/A sky130_fd_sc_hd__clkbuf_2
Xuser_to_mprj_oen_buffers\[108\] _371_/Y mprj_logic_high_inst/HI[310] vssd vssd vccd
+ vccd la_oenb_core[108] sky130_fd_sc_hd__einvp_8
Xinput459 mprj_we_o_core vssd vssd vccd vccd _395_/A sky130_fd_sc_hd__clkbuf_2
Xinput448 mprj_dat_o_core[5] vssd vssd vccd vccd _437_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[38\] _630_/Y mprj_logic_high_inst/HI[240] vssd vssd vccd
+ vccd la_oenb_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_44_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input206_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__572__A _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[1\]_A _433_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high_inst/HI[269] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd vssd vccd vccd output548/A
+ sky130_fd_sc_hd__clkinv_2
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__482__A _482_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A _657_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput201 la_iena_mprj[47] vssd vssd vccd vccd input201/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input156_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput234 la_iena_mprj[77] vssd vssd vccd vccd input234/X sky130_fd_sc_hd__clkbuf_1
Xinput223 la_iena_mprj[67] vssd vssd vccd vccd input223/X sky130_fd_sc_hd__clkbuf_1
Xinput212 la_iena_mprj[57] vssd vssd vccd vccd input212/X sky130_fd_sc_hd__clkbuf_1
Xinput245 la_iena_mprj[87] vssd vssd vccd vccd input245/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input323_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput256 la_iena_mprj[97] vssd vssd vccd vccd input256/X sky130_fd_sc_hd__clkbuf_1
Xinput267 la_oenb_mprj[106] vssd vssd vccd vccd _369_/A sky130_fd_sc_hd__buf_2
Xinput278 la_oenb_mprj[116] vssd vssd vccd vccd _379_/A sky130_fd_sc_hd__clkbuf_4
X_653_ _653_/A vssd vssd vccd vccd _653_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input17_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput289 la_oenb_mprj[126] vssd vssd vccd vccd _389_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__567__A _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_584_ _584_/A vssd vssd vccd vccd _584_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf\[65\] _529_/Y la_buf\[65\]/TE vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_44_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[121\] _585_/Y la_buf\[121\]/TE vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[29\] _429_/Y mprj_adr_buf\[29\]/TE vssd vssd vccd vccd mprj_adr_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_45_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__477__A _477_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] user_to_mprj_in_gates\[54\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input9_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__387__A _387_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input273_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input440_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[101\]_A_N _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_636_ _636_/A vssd vssd vccd vccd _636_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_44_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[116\]_A_N _379_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_567_ _567_/A vssd vssd vccd vccd _567_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[94\]_A _558_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_498_ _498_/A vssd vssd vccd vccd _498_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd vssd vccd vccd output507/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_16_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput527 output527/A vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_2
Xoutput505 output505/A vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_2
Xoutput516 output516/A vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_2
Xoutput549 output549/A vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_2
Xoutput538 output538/A vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_2
XFILLER_29_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[64\] input220/X mprj_logic_high_inst/HI[394] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[64\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[42\] _634_/A la_buf_enable\[42\]/B vssd vssd vccd vccd la_buf\[42\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[2\] _594_/Y mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd la_oenb_core[2] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[20\] _612_/Y mprj_logic_high_inst/HI[222] vssd vssd vccd
+ vccd la_oenb_core[20] sky130_fd_sc_hd__einvp_8
XFILLER_26_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input119_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_421_ _421_/A vssd vssd vccd vccd _421_/Y sky130_fd_sc_hd__inv_12
XFILLER_53_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_352_ _352_/A vssd vssd vccd vccd _352_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input390_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[94\]_B la_buf_enable\[94\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input84_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[28\] _492_/Y la_buf\[28\]/TE vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__einvp_8
XFILLER_13_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput9 la_data_out_mprj[104] vssd vssd vccd vccd _568_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_619_ _619_/A vssd vssd vccd vccd _619_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] user_to_mprj_in_gates\[17\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[85\]_B la_buf_enable\[85\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[27\] user_wb_dat_gates\[27\]/Y vssd vssd vccd vccd output611/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_25_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[76\]_B la_buf_enable\[76\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[68\] _331_/Y mprj_logic_high_inst/HI[270] vssd vssd vccd
+ vccd la_oenb_core[68] sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[17\]_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[16\] _448_/Y mprj_dat_buf\[16\]/TE vssd vssd vccd vccd mprj_dat_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input236_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input403_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__575__A _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_404_ _404_/A vssd vssd vccd vccd _404_/Y sky130_fd_sc_hd__inv_2
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_335_ _335_/A vssd vssd vccd vccd _335_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_B la_buf_enable\[67\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[11\] _411_/Y mprj_adr_buf\[11\]/TE vssd vssd vccd vccd mprj_adr_o_user[11]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd vssd vccd vccd
+ output491/A sky130_fd_sc_hd__clkinv_4
XFILLER_2_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output622_A output622/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd vssd vccd vccd output581/A
+ sky130_fd_sc_hd__inv_2
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__485__A _485_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[1\] user_wb_dat_gates\[1\]/Y vssd vssd vccd vccd output603/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_0_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[61\]_B mprj_logic_high_inst/HI[391] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[27\] input179/X mprj_logic_high_inst/HI[357] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[27\]/B sky130_fd_sc_hd__and2_1
XFILLER_52_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[51\]_A _643_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input186_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input353_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input47_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[110\] _373_/A la_buf_enable\[110\]/B vssd vssd vccd vccd la_buf\[110\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[74\]_A_N _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[95\] _559_/Y la_buf\[95\]/TE vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[0\] input132/X mprj_logic_high_inst/HI[330] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[0\]/B sky130_fd_sc_hd__and2_1
XFILLER_19_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[89\]_A_N _352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[52\]_B mprj_logic_high_inst/HI[382] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[12\]_A_N _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput12 la_data_out_mprj[107] vssd vssd vccd vccd _571_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[9\]_A input259/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput45 la_data_out_mprj[21] vssd vssd vccd vccd _485_/A sky130_fd_sc_hd__clkbuf_2
Xinput23 la_data_out_mprj[117] vssd vssd vccd vccd _581_/A sky130_fd_sc_hd__clkbuf_4
Xinput34 la_data_out_mprj[127] vssd vssd vccd vccd _591_/A sky130_fd_sc_hd__buf_2
XFILLER_11_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput89 la_data_out_mprj[61] vssd vssd vccd vccd _525_/A sky130_fd_sc_hd__clkbuf_2
Xinput78 la_data_out_mprj[51] vssd vssd vccd vccd _515_/A sky130_fd_sc_hd__clkbuf_2
Xinput67 la_data_out_mprj[41] vssd vssd vccd vccd _505_/A sky130_fd_sc_hd__clkbuf_2
Xinput56 la_data_out_mprj[31] vssd vssd vccd vccd _495_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[27\]_A_N _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] user_to_mprj_in_gates\[84\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[43\]_B mprj_logic_high_inst/HI[373] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[33\]_A _625_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput416 mprj_adr_o_core[6] vssd vssd vccd vccd _406_/A sky130_fd_sc_hd__clkbuf_2
Xinput427 mprj_dat_o_core[15] vssd vssd vccd vccd _447_/A sky130_fd_sc_hd__buf_4
Xinput405 mprj_adr_o_core[25] vssd vssd vccd vccd _425_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput449 mprj_dat_o_core[6] vssd vssd vccd vccd _438_/A sky130_fd_sc_hd__clkbuf_4
Xinput438 mprj_dat_o_core[25] vssd vssd vccd vccd _457_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input101_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[34\]_B mprj_logic_high_inst/HI[364] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[112\]_TE mprj_logic_high_inst/HI[314] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[6\] _470_/Y la_buf\[6\]/TE vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__einvp_8
XFILLER_7_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[10\] _474_/Y la_buf\[10\]/TE vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_4_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[3\] _403_/Y mprj_adr_buf\[3\]/TE vssd vssd vccd vccd mprj_adr_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_47_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[20\]_A _420_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd vssd vccd vccd output540/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_1_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[25\]_B mprj_logic_high_inst/HI[355] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[12\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[15\]_A _607_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] user_to_mprj_in_gates\[110\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_mprj_adr_buf\[11\]_A _411_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[16\]_B mprj_logic_high_inst/HI[346] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[9\]_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[94\] input253/X mprj_logic_high_inst/HI[424] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[94\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[120\] _383_/Y mprj_logic_high_inst/HI[322] vssd vssd vccd
+ vccd la_oenb_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_44_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _397_/Y mprj_sel_buf\[1\]/TE vssd vssd vccd vccd mprj_sel_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput202 la_iena_mprj[48] vssd vssd vccd vccd input202/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput235 la_iena_mprj[78] vssd vssd vccd vccd input235/X sky130_fd_sc_hd__clkbuf_1
Xinput224 la_iena_mprj[68] vssd vssd vccd vccd input224/X sky130_fd_sc_hd__clkbuf_1
Xinput213 la_iena_mprj[58] vssd vssd vccd vccd input213/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input149_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[72\] _335_/A la_buf_enable\[72\]/B vssd vssd vccd vccd la_buf\[72\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_40_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[50\] _642_/Y mprj_logic_high_inst/HI[252] vssd vssd vccd
+ vccd la_oenb_core[50] sky130_fd_sc_hd__einvp_8
Xinput246 la_iena_mprj[88] vssd vssd vccd vccd input246/X sky130_fd_sc_hd__clkbuf_1
Xinput257 la_iena_mprj[98] vssd vssd vccd vccd input257/X sky130_fd_sc_hd__clkbuf_1
Xinput268 la_oenb_mprj[107] vssd vssd vccd vccd _370_/A sky130_fd_sc_hd__clkbuf_4
Xinput279 la_oenb_mprj[117] vssd vssd vccd vccd _380_/A sky130_fd_sc_hd__clkbuf_4
X_652_ _652_/A vssd vssd vccd vccd _652_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input316_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_583_ _583_/A vssd vssd vccd vccd _583_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[58\] _522_/Y la_buf\[58\]/TE vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__einvp_8
XANTENNA__583__A _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[114\] _578_/Y la_buf\[114\]/TE vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__einvp_8
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] user_to_mprj_in_gates\[47\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] user_to_mprj_in_gates\[9\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[98\] _361_/Y mprj_logic_high_inst/HI[300] vssd vssd vccd
+ vccd la_oenb_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_6_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input266_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input433_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_635_ _635_/A vssd vssd vccd vccd _635_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_dat_buf\[24\]_A _456_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_566_ _566_/A vssd vssd vccd vccd _566_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_497_ _497_/A vssd vssd vccd vccd _497_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output485_A output485/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd vssd vccd vccd output499/A
+ sky130_fd_sc_hd__inv_2
XFILLER_47_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput506 output506/A vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_2
Xoutput517 output517/A vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_2
XFILLER_47_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput539 output539/A vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_2
Xoutput528 output528/A vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_2
XFILLER_25_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__488__A _488_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[15\]_A _447_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__398__A _398_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[57\] input212/X mprj_logic_high_inst/HI[387] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[57\]/B sky130_fd_sc_hd__and2_1
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[13\]_A user_wb_dat_gates\[13\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ _420_/A vssd vssd vccd vccd _420_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_14_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[13\] _605_/Y mprj_logic_high_inst/HI[215] vssd vssd vccd
+ vccd la_oenb_core[13] sky130_fd_sc_hd__einvp_8
X_351_ _351_/A vssd vssd vccd vccd _351_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[35\] _627_/A la_buf_enable\[35\]/B vssd vssd vccd vccd la_buf\[35\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd vssd vccd vccd output590/A
+ sky130_fd_sc_hd__inv_6
XANTENNA_input383_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input77_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_618_ _618_/A vssd vssd vccd vccd _618_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_549_ _549_/A vssd vssd vccd vccd _549_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[26\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_A_N _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[115\]_A_N _378_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[17\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input131_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input229_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _403_/A vssd vssd vccd vccd _403_/Y sky130_fd_sc_hd__inv_12
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[40\] _504_/Y la_buf\[40\]/TE vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__einvp_8
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_334_ _334_/A vssd vssd vccd vccd _334_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__591__A _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[112\] input146/X mprj_logic_high_inst/HI[442] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[112\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd vssd vccd vccd
+ output483/A sky130_fd_sc_hd__clkinv_4
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output615_A output615/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd vssd vccd vccd output573/A
+ sky130_fd_sc_hd__inv_2
XFILLER_37_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_A _409_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _343_/Y mprj_logic_high_inst/HI[282] vssd vssd vccd
+ vccd la_oenb_core[80] sky130_fd_sc_hd__einvp_8
XANTENNA_input179_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input346_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[88\] _552_/Y la_buf\[88\]/TE vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__einvp_8
XANTENNA__586__A _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[103\] _366_/A la_buf_enable\[103\]/B vssd vssd vccd vccd la_buf\[103\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput13 la_data_out_mprj[108] vssd vssd vccd vccd _572_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[9\]_B mprj_logic_high_inst/HI[339] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput35 la_data_out_mprj[12] vssd vssd vccd vccd _476_/A sky130_fd_sc_hd__clkbuf_2
Xinput46 la_data_out_mprj[22] vssd vssd vccd vccd _486_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput24 la_data_out_mprj[118] vssd vssd vccd vccd _582_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput79 la_data_out_mprj[52] vssd vssd vccd vccd _516_/A sky130_fd_sc_hd__clkbuf_2
Xinput68 la_data_out_mprj[42] vssd vssd vccd vccd _506_/A sky130_fd_sc_hd__clkbuf_2
Xinput57 la_data_out_mprj[32] vssd vssd vccd vccd _496_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] user_to_mprj_in_gates\[77\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__496__A _496_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput417 mprj_adr_o_core[7] vssd vssd vccd vccd _407_/A sky130_fd_sc_hd__clkbuf_2
Xinput428 mprj_dat_o_core[16] vssd vssd vccd vccd _448_/A sky130_fd_sc_hd__clkbuf_4
Xinput406 mprj_adr_o_core[26] vssd vssd vccd vccd _426_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput439 mprj_dat_o_core[26] vssd vssd vccd vccd _458_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input296_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd vssd vccd vccd output532/A
+ sky130_fd_sc_hd__inv_2
XFILLER_15_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] user_to_mprj_in_gates\[103\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[73\]_A_N _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[88\]_A_N _351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[87\] input245/X mprj_logic_high_inst/HI[417] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[87\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[113\] _376_/Y mprj_logic_high_inst/HI[315] vssd vssd vccd
+ vccd la_oenb_core[113] sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _392_/Y mprj_clk2_buf/TE vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__einvp_8
XFILLER_1_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput225 la_iena_mprj[69] vssd vssd vccd vccd input225/X sky130_fd_sc_hd__clkbuf_1
Xinput214 la_iena_mprj[59] vssd vssd vccd vccd input214/X sky130_fd_sc_hd__clkbuf_1
Xinput203 la_iena_mprj[49] vssd vssd vccd vccd input203/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput236 la_iena_mprj[79] vssd vssd vccd vccd input236/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_A_N _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput247 la_iena_mprj[89] vssd vssd vccd vccd input247/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput258 la_iena_mprj[99] vssd vssd vccd vccd input258/X sky130_fd_sc_hd__clkbuf_1
Xinput269 la_oenb_mprj[108] vssd vssd vccd vccd _371_/A sky130_fd_sc_hd__buf_4
Xuser_to_mprj_oen_buffers\[43\] _635_/Y mprj_logic_high_inst/HI[245] vssd vssd vccd
+ vccd la_oenb_core[43] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[65\] _657_/A la_buf_enable\[65\]/B vssd vssd vccd vccd la_buf\[65\]/TE
+ sky130_fd_sc_hd__and2b_1
X_651_ _651_/A vssd vssd vccd vccd _651_/Y sky130_fd_sc_hd__inv_2
Xuser_irq_buffers\[1\] user_irq_gates\[1\]/Y vssd vssd vccd vccd output629/A sky130_fd_sc_hd__clkinv_4
XFILLER_44_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_582_ _582_/A vssd vssd vccd vccd _582_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input211_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input309_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[107\] _571_/Y la_buf\[107\]/TE vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_45_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd vssd vccd vccd
+ output464/A sky130_fd_sc_hd__clkinv_4
XFILLER_47_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input259_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input161_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input426_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input22_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_634_ _634_/A vssd vssd vccd vccd _634_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[70\] _534_/Y la_buf\[70\]/TE vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_45_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__594__A _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_565_ _565_/A vssd vssd vccd vccd _565_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_496_ _496_/A vssd vssd vccd vccd _496_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput507 output507/A vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_2
Xoutput518 output518/A vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_2
Xoutput529 output529/A vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_2
XFILLER_45_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high_inst/HI[226] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _350_/A vssd vssd vccd vccd _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[28\] _620_/A la_buf_enable\[28\]/B vssd vssd vccd vccd la_buf\[28\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input376_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__589__A _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_617_ _617_/A vssd vssd vccd vccd _617_/Y sky130_fd_sc_hd__clkinv_2
X_548_ _548_/A vssd vssd vccd vccd _548_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output595_A output595/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_479_ _479_/A vssd vssd vccd vccd _479_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[9\]_B la_buf_enable\[9\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input124_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_402_ _402_/A vssd vssd vccd vccd _402_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_333_ _333_/A vssd vssd vccd vccd _333_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[33\] _497_/Y la_buf\[33\]/TE vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[105\] input138/X mprj_logic_high_inst/HI[435] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[105\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd vssd vccd vccd output565/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_4_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output608_A output608/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] user_to_mprj_in_gates\[22\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[46\]_A input200/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[73\] _336_/Y mprj_logic_high_inst/HI[275] vssd vssd vccd
+ vccd la_oenb_core[73] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[95\] _358_/A la_buf_enable\[95\]/B vssd vssd vccd vccd la_buf\[95\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[21\] _453_/Y mprj_dat_buf\[21\]/TE vssd vssd vccd vccd mprj_dat_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input339_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input241_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput36 la_data_out_mprj[13] vssd vssd vccd vccd _477_/A sky130_fd_sc_hd__clkbuf_2
Xinput14 la_data_out_mprj[109] vssd vssd vccd vccd _573_/A sky130_fd_sc_hd__clkbuf_4
Xinput25 la_data_out_mprj[119] vssd vssd vccd vccd _583_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput69 la_data_out_mprj[43] vssd vssd vccd vccd _507_/A sky130_fd_sc_hd__clkbuf_2
Xinput47 la_data_out_mprj[23] vssd vssd vccd vccd _487_/A sky130_fd_sc_hd__clkbuf_2
Xinput58 la_data_out_mprj[33] vssd vssd vccd vccd _497_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[114\]_A_N _377_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[1\] _593_/A la_buf_enable\[1\]/B vssd vssd vccd vccd la_buf\[1\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput418 mprj_adr_o_core[8] vssd vssd vccd vccd _408_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput407 mprj_adr_o_core[27] vssd vssd vccd vccd _427_/A sky130_fd_sc_hd__buf_2
Xinput429 mprj_dat_o_core[17] vssd vssd vccd vccd _449_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[32\] input185/X mprj_logic_high_inst/HI[362] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[32\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[10\] _602_/A la_buf_enable\[10\]/B vssd vssd vccd vccd la_buf\[10\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_input191_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input289_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input456_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input52_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__597__A _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[102\]_A _566_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput226 la_iena_mprj[6] vssd vssd vccd vccd input226/X sky130_fd_sc_hd__clkbuf_2
Xinput215 la_iena_mprj[5] vssd vssd vccd vccd input215/X sky130_fd_sc_hd__buf_2
Xinput204 la_iena_mprj[4] vssd vssd vccd vccd input204/X sky130_fd_sc_hd__buf_2
XFILLER_40_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _369_/Y mprj_logic_high_inst/HI[308] vssd vssd vccd
+ vccd la_oenb_core[106] sky130_fd_sc_hd__einvp_8
Xinput259 la_iena_mprj[9] vssd vssd vccd vccd input259/X sky130_fd_sc_hd__buf_2
Xinput248 la_iena_mprj[8] vssd vssd vccd vccd input248/X sky130_fd_sc_hd__clkbuf_4
Xinput237 la_iena_mprj[7] vssd vssd vccd vccd input237/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_650_ _650_/A vssd vssd vccd vccd _650_/Y sky130_fd_sc_hd__clkinv_2
X_581_ _581_/A vssd vssd vccd vccd _581_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[58\] _650_/A la_buf_enable\[58\]/B vssd vssd vccd vccd la_buf\[58\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[36\] _628_/Y mprj_logic_high_inst/HI[238] vssd vssd vccd
+ vccd la_oenb_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_22_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input204_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[97\]_A _561_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[120\]_B mprj_logic_high_inst/HI[450] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[111\]_B mprj_logic_high_inst/HI[441] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input154_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[30\]_B la_buf_enable\[30\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input321_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_633_ _633_/A vssd vssd vccd vccd _633_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input15_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input419_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_564_ _564_/A vssd vssd vccd vccd _564_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[63\] _527_/Y la_buf\[63\]/TE vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__einvp_8
XFILLER_38_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_495_ _495_/A vssd vssd vccd vccd _495_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[102\]_B mprj_logic_high_inst/HI[432] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[97\]_B la_buf_enable\[97\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[27\] _427_/Y mprj_adr_buf\[27\]/TE vssd vssd vccd vccd mprj_adr_o_user[27]
+ sky130_fd_sc_hd__einvp_8
Xoutput508 output508/A vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_2
XFILLER_5_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput519 output519/A vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_2
XFILLER_10_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_ack_gate mprj_ack_i_user user_wb_ack_gate/B vssd vssd vccd vccd user_wb_ack_gate/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_49_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[21\]_B la_buf_enable\[21\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[72\]_A_N _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] user_to_mprj_in_gates\[52\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[87\]_A_N _350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[88\]_B la_buf_enable\[88\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[10\]_A_N _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[25\]_A_N _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[29\]_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[12\]_B la_buf_enable\[12\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[91\]_B mprj_logic_high_inst/HI[421] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[79\]_B la_buf_enable\[79\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input271_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input369_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[126\] _389_/A la_buf_enable\[126\]/B vssd vssd vccd vccd la_buf\[126\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_616_ _616_/A vssd vssd vccd vccd _616_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_547_ _547_/A vssd vssd vccd vccd _547_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_17_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_478_ _478_/A vssd vssd vccd vccd _478_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd vssd vccd vccd output505/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[63\]_A _655_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[62\] input218/X mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[62\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[40\] _632_/A la_buf_enable\[40\]/B vssd vssd vccd vccd la_buf\[40\]/TE
+ sky130_fd_sc_hd__and2b_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[0\] _592_/Y mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd la_oenb_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_27_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_401_ _401_/A vssd vssd vccd vccd _401_/Y sky130_fd_sc_hd__inv_12
XANTENNA_input117_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_332_ _332_/A vssd vssd vccd vccd _332_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_A _646_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input82_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[26\] _490_/Y la_buf\[26\]/TE vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_6_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[55\]_B mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[28\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_33_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] user_to_mprj_in_gates\[15\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_oen_buffers\[45\]_A _637_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[25\] user_wb_dat_gates\[25\]/Y vssd vssd vccd vccd output609/A
+ sky130_fd_sc_hd__inv_6
XFILLER_29_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] user_to_mprj_in_gates\[126\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[46\]_B mprj_logic_high_inst/HI[376] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_A _628_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[66\] _329_/Y mprj_logic_high_inst/HI[268] vssd vssd vccd
+ vccd la_oenb_core[66] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[88\] _351_/A la_buf_enable\[88\]/B vssd vssd vccd vccd la_buf\[88\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[14\] _446_/Y mprj_dat_buf\[14\]/TE vssd vssd vccd vccd mprj_dat_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input234_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[37\]_B mprj_logic_high_inst/HI[367] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input401_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high_inst/HI[239] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput15 la_data_out_mprj[10] vssd vssd vccd vccd _474_/A sky130_fd_sc_hd__clkbuf_2
Xinput26 la_data_out_mprj[11] vssd vssd vccd vccd _475_/A sky130_fd_sc_hd__clkbuf_2
Xinput37 la_data_out_mprj[14] vssd vssd vccd vccd _478_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 la_data_out_mprj[24] vssd vssd vccd vccd _488_/A sky130_fd_sc_hd__clkbuf_2
Xinput59 la_data_out_mprj[34] vssd vssd vccd vccd _498_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd vssd vccd vccd
+ output489/A sky130_fd_sc_hd__clkinv_4
XFILLER_2_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output620_A output620/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[23\]_A _423_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[28\]_B mprj_logic_high_inst/HI[358] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vssd vccd vccd _409_/A sky130_fd_sc_hd__clkbuf_2
Xinput408 mprj_adr_o_core[28] vssd vssd vccd vccd _428_/A sky130_fd_sc_hd__buf_2
XFILLER_9_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_A _414_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[19\]_B mprj_logic_high_inst/HI[349] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[25\] input177/X mprj_logic_high_inst/HI[355] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[25\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input184_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input351_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input449_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input45_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[93\] _557_/Y la_buf\[93\]/TE vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] user_to_mprj_in_gates\[82\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_1
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput227 la_iena_mprj[70] vssd vssd vccd vccd input227/X sky130_fd_sc_hd__clkbuf_1
Xinput216 la_iena_mprj[60] vssd vssd vccd vccd input216/X sky130_fd_sc_hd__clkbuf_1
Xinput205 la_iena_mprj[50] vssd vssd vccd vccd input205/X sky130_fd_sc_hd__clkbuf_1
Xinput238 la_iena_mprj[80] vssd vssd vccd vccd input238/X sky130_fd_sc_hd__clkbuf_1
Xinput249 la_iena_mprj[90] vssd vssd vccd vccd input249/X sky130_fd_sc_hd__clkbuf_1
X_580_ _580_/A vssd vssd vccd vccd _580_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[29\] _621_/Y mprj_logic_high_inst/HI[231] vssd vssd vccd
+ vccd la_oenb_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_51_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input399_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[4\] _468_/Y la_buf\[4\]/TE vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__einvp_8
XFILLER_49_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[113\]_A_N _376_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[1\] _401_/Y mprj_adr_buf\[1\]/TE vssd vssd vccd vccd mprj_adr_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[27\]_A _459_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd vssd vccd vccd output538/A
+ sky130_fd_sc_hd__inv_2
XFILLER_1_1554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[10\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[18\]_A _450_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[92\] input251/X mprj_logic_high_inst/HI[422] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[92\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input147_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[70\] _333_/A la_buf_enable\[70\]/B vssd vssd vccd vccd la_buf\[70\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_632_ _632_/A vssd vssd vccd vccd _632_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_wb_dat_buffers\[16\]_A user_wb_dat_gates\[16\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input314_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_563_ _563_/A vssd vssd vccd vccd _563_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf\[56\] _520_/Y la_buf\[56\]/TE vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_44_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_494_ _494_/A vssd vssd vccd vccd _494_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_wb_ena_buf input453/X user_to_mprj_wb_ena_buf/B vssd vssd vccd vccd
+ user_wb_ack_gate/B sky130_fd_sc_hd__and2_4
XFILLER_9_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput509 output509/A vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_2
Xla_buf\[112\] _576_/Y la_buf\[112\]/TE vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__einvp_8
XFILLER_10_1172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[120\]_B la_buf_enable\[120\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] user_to_mprj_in_gates\[45\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_23_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] user_to_mprj_in_gates\[7\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_wb_dat_gates\[29\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[111\]_B la_buf_enable\[111\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high_inst/HI[272] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_buffers\[2\]_A user_wb_dat_gates\[2\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[96\] _359_/Y mprj_logic_high_inst/HI[298] vssd vssd vccd
+ vccd la_oenb_core[96] sky130_fd_sc_hd__einvp_8
XFILLER_30_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input264_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[9\] input259/X mprj_logic_high_inst/HI[339] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[9\]/B sky130_fd_sc_hd__and2_1
XFILLER_7_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[119\] _382_/A la_buf_enable\[119\]/B vssd vssd vccd vccd la_buf\[119\]/TE
+ sky130_fd_sc_hd__and2b_2
XFILLER_37_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_615_ _615_/A vssd vssd vccd vccd _615_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_546_ _546_/A vssd vssd vccd vccd _546_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[102\]_B la_buf_enable\[102\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_477_ _477_/A vssd vssd vccd vccd _477_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd vssd vccd vccd output497/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj2_pwrgood mprj2_pwrgood/A vssd vssd vccd vccd output626/A sky130_fd_sc_hd__buf_12
XFILLER_8_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[55\] input210/X mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[55\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_400_ _400_/A vssd vssd vccd vccd _400_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_42_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[11\] _603_/Y mprj_logic_high_inst/HI[213] vssd vssd vccd
+ vccd la_oenb_core[11] sky130_fd_sc_hd__einvp_8
XFILLER_39_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _331_/A vssd vssd vccd vccd _331_/Y sky130_fd_sc_hd__inv_2
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[33\] _625_/A la_buf_enable\[33\]/B vssd vssd vccd vccd la_buf\[33\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd vssd vccd vccd output568/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_35_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input381_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[71\]_A_N _334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[19\] _483_/Y la_buf\[19\]/TE vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__einvp_8
XANTENNA_input75_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_A_N _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[24\]_A_N _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[3\]_A user_to_mprj_in_gates\[3\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_529_ _529_/A vssd vssd vccd vccd _529_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[18\] user_wb_dat_gates\[18\]/Y vssd vssd vccd vccd output601/A
+ sky130_fd_sc_hd__inv_6
XFILLER_29_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] user_to_mprj_in_gates\[119\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[59\] _651_/Y mprj_logic_high_inst/HI[261] vssd vssd vccd
+ vccd la_oenb_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_8_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input227_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[110\] input144/X mprj_logic_high_inst/HI[440] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[110\]/B sky130_fd_sc_hd__and2_1
XFILLER_50_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput16 la_data_out_mprj[110] vssd vssd vccd vccd _574_/A sky130_fd_sc_hd__clkbuf_4
Xinput27 la_data_out_mprj[120] vssd vssd vccd vccd _584_/A sky130_fd_sc_hd__buf_2
XFILLER_11_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput38 la_data_out_mprj[15] vssd vssd vccd vccd _479_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput49 la_data_out_mprj[25] vssd vssd vccd vccd _489_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__404__A _404_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd vssd vccd vccd
+ output481/A sky130_fd_sc_hd__clkinv_4
XFILLER_42_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output613_A output613/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd vssd vccd vccd output571/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_0_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_0_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput409 mprj_adr_o_core[29] vssd vssd vccd vccd _429_/A sky130_fd_sc_hd__buf_2
XFILLER_44_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high_inst/HI[307] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[18\] input169/X mprj_logic_high_inst/HI[348] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[18\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input177_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input344_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input38_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[86\] _550_/Y la_buf\[86\]/TE vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_21_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[101\] _364_/A la_buf_enable\[101\]/B vssd vssd vccd vccd la_buf\[101\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] user_to_mprj_in_gates\[75\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput217 la_iena_mprj[61] vssd vssd vccd vccd input217/X sky130_fd_sc_hd__clkbuf_1
Xinput206 la_iena_mprj[51] vssd vssd vccd vccd input206/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput228 la_iena_mprj[71] vssd vssd vccd vccd input228/X sky130_fd_sc_hd__clkbuf_1
Xinput239 la_iena_mprj[81] vssd vssd vccd vccd input239/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input294_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input461_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_ena_buf\[1\] input461/X user_irq_ena_buf\[1\]/B vssd vssd vccd vccd user_irq_gates\[1\]/B
+ sky130_fd_sc_hd__and2_1
XFILLER_45_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd vssd vccd vccd output530/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] user_to_mprj_in_gates\[101\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_1
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[85\] input243/X mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[85\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[111\] _374_/Y mprj_logic_high_inst/HI[313] vssd vssd vccd
+ vccd la_oenb_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_44_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[41\] _633_/Y mprj_logic_high_inst/HI[243] vssd vssd vccd
+ vccd la_oenb_core[41] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[63\] _655_/A la_buf_enable\[63\]/B vssd vssd vccd vccd la_buf\[63\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_631_ _631_/A vssd vssd vccd vccd _631_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_562_ _562_/A vssd vssd vccd vccd _562_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input307_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_493_ _493_/A vssd vssd vccd vccd _493_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_44_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[49\] _513_/Y la_buf\[49\]/TE vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[105\] _569_/Y la_buf\[105\]/TE vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_45_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] user_to_mprj_in_gates\[38\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[112\]_A_N _375_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[127\]_A_N _390_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[89\] _352_/Y mprj_logic_high_inst/HI[291] vssd vssd vccd
+ vccd la_oenb_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_2_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input257_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input20_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input424_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_614_ _614_/A vssd vssd vccd vccd _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_545_ _545_/A vssd vssd vccd vccd _545_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_476_ _476_/A vssd vssd vccd vccd _476_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[48\] input202/X mprj_logic_high_inst/HI[378] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[48\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ _330_/A vssd vssd vccd vccd _330_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[26\] _618_/A la_buf_enable\[26\]/B vssd vssd vccd vccd la_buf\[26\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input374_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input68_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_528_ _528_/A vssd vssd vccd vccd _528_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output593_A output593/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_459_ _459_/A vssd vssd vccd vccd _459_/Y sky130_fd_sc_hd__inv_6
XFILLER_31_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high_inst/HI[262] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__510__A _510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input122_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_41 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[31\] _495_/Y la_buf\[31\]/TE vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__einvp_8
Xinput17 la_data_out_mprj[111] vssd vssd vccd vccd _575_/A sky130_fd_sc_hd__buf_4
Xinput28 la_data_out_mprj[121] vssd vssd vccd vccd _585_/A sky130_fd_sc_hd__clkbuf_2
Xuser_to_mprj_in_ena_buf\[103\] input136/X mprj_logic_high_inst/HI[433] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[103\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[3\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput39 la_data_out_mprj[16] vssd vssd vccd vccd _480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd vssd vccd vccd
+ output473/A sky130_fd_sc_hd__clkinv_4
XFILLER_38_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd vssd vccd vccd output563/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output606_A output606/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] user_to_mprj_in_gates\[20\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[114\]_A _578_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_buffers\[30\] user_wb_dat_gates\[30\]/Y vssd vssd vccd vccd output615/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__330__A _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[8\] _440_/Y mprj_dat_buf\[8\]/TE vssd vssd vccd vccd mprj_dat_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_44_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[70\]_A_N _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[10\]_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[85\]_A_N _348_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__505__A _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[71\] _334_/Y mprj_logic_high_inst/HI[273] vssd vssd vccd
+ vccd la_oenb_core[71] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[23\]_A_N _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[93\] _356_/A la_buf_enable\[93\]/B vssd vssd vccd vccd la_buf\[93\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_43_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput490 output490/A vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_2
XFILLER_43_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input337_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[79\] _543_/Y la_buf\[79\]/TE vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_21_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] user_to_mprj_in_gates\[68\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[123\]_B mprj_logic_high_inst/HI[453] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_A _488_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[42\]_B la_buf_enable\[42\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput218 la_iena_mprj[62] vssd vssd vccd vccd input218/X sky130_fd_sc_hd__clkbuf_1
Xinput207 la_iena_mprj[52] vssd vssd vccd vccd input207/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vssd vccd vccd input229/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[114\]_B mprj_logic_high_inst/HI[444] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[30\] input183/X mprj_logic_high_inst/HI[360] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[30\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input287_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input454_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[33\]_B la_buf_enable\[33\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input50_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[105\]_B mprj_logic_high_inst/HI[435] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd vssd vccd vccd output522/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_30_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[24\]_B la_buf_enable\[24\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[15\]_B la_buf_enable\[15\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[78\] input235/X mprj_logic_high_inst/HI[408] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[78\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[104\] _367_/Y mprj_logic_high_inst/HI[306] vssd vssd vccd
+ vccd la_oenb_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[94\]_B mprj_logic_high_inst/HI[424] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_630_ _630_/A vssd vssd vccd vccd _630_/Y sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[56\] _648_/A la_buf_enable\[56\]/B vssd vssd vccd vccd la_buf\[56\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[34\] _626_/Y mprj_logic_high_inst/HI[236] vssd vssd vccd
+ vccd la_oenb_core[34] sky130_fd_sc_hd__einvp_8
XFILLER_22_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_561_ _561_/A vssd vssd vccd vccd _561_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_44_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_492_ _492_/A vssd vssd vccd vccd _492_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input202_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input98_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[85\]_B mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high_inst/HI[219] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__603__A _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input152_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_613_ _613_/A vssd vssd vccd vccd _613_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input417_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input13_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[61\] _525_/Y la_buf\[61\]/TE vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_44_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_544_ _544_/A vssd vssd vccd vccd _544_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_475_ _475_/A vssd vssd vccd vccd _475_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[57\]_A _649_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[25\] _425_/Y mprj_adr_buf\[25\]/TE vssd vssd vccd vccd mprj_adr_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[58\]_B mprj_logic_high_inst/HI[388] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] user_to_mprj_in_gates\[50\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_1
Xinput390 mprj_adr_o_core[11] vssd vssd vccd vccd _411_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_A _640_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__333__A _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[49\]_B mprj_logic_high_inst/HI[379] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[19\] _611_/A la_buf_enable\[19\]/B vssd vssd vccd vccd la_buf\[19\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_52_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input367_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[2\] user_irq_core[2] user_irq_gates\[2\]/B vssd vssd vccd vccd user_irq_gates\[2\]/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_46_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[124\] _387_/A la_buf_enable\[124\]/B vssd vssd vccd vccd la_buf\[124\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_527_ _527_/A vssd vssd vccd vccd _527_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_458_ _458_/A vssd vssd vccd vccd _458_/Y sky130_fd_sc_hd__inv_4
XFILLER_53_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_389_ _389_/A vssd vssd vccd vccd _389_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd vssd vccd vccd output503/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_9_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] user_to_mprj_in_gates\[98\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[26\]_A _426_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[111\]_A_N _374_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[126\]_A_N _389_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[17\]_A _417_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[60\] input216/X mprj_logic_high_inst/HI[390] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[60\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input115_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input80_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput18 la_data_out_mprj[112] vssd vssd vccd vccd _576_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[24\] _488_/Y la_buf\[24\]/TE vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__einvp_8
XFILLER_32_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput29 la_data_out_mprj[122] vssd vssd vccd vccd _586_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd vssd vccd vccd output555/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_45_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[26\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_53_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] user_to_mprj_in_gates\[13\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[23\] user_wb_dat_gates\[23\]/Y vssd vssd vccd vccd output607/A
+ sky130_fd_sc_hd__inv_6
XANTENNA__611__A _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] user_to_mprj_in_gates\[124\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__521__A _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput480 output480/A vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_2
XFILLER_43_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[64\] _656_/Y mprj_logic_high_inst/HI[266] vssd vssd vccd
+ vccd la_oenb_core[64] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[86\] _349_/A la_buf_enable\[86\]/B vssd vssd vccd vccd la_buf\[86\]/TE
+ sky130_fd_sc_hd__and2b_1
Xoutput491 output491/A vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_2
XFILLER_43_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[12\] _444_/Y mprj_dat_buf\[12\]/TE vssd vssd vccd vccd mprj_dat_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input232_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_cyc_buf_A _393_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd vssd vccd vccd
+ output487/A sky130_fd_sc_hd__clkinv_4
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__606__A _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[2\]_A _402_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__341__A _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput208 la_iena_mprj[53] vssd vssd vccd vccd input208/X sky130_fd_sc_hd__clkbuf_1
Xinput219 la_iena_mprj[63] vssd vssd vccd vccd input219/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high_inst/HI[275] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[23\] input175/X mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[23\]/B sky130_fd_sc_hd__and2_1
XANTENNA__516__A _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input182_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input447_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input43_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[2\]_B mprj_logic_high_inst/HI[332] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[91\] _555_/Y la_buf\[91\]/TE vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_23_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] user_to_mprj_in_gates\[80\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[84\]_A_N _347_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[123\]_B la_buf_enable\[123\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[99\]_A_N _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_A_N _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__336__A _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[114\]_B la_buf_enable\[114\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_560_ _560_/A vssd vssd vccd vccd _560_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[27\] _619_/Y mprj_logic_high_inst/HI[229] vssd vssd vccd
+ vccd la_oenb_core[27] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[49\] _641_/A la_buf_enable\[49\]/B vssd vssd vccd vccd la_buf\[49\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[9\] _601_/Y mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd la_oenb_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_491_ _491_/A vssd vssd vccd vccd _491_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input397_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[2\] _466_/Y la_buf\[2\]/TE vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_49_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[105\]_B la_buf_enable\[105\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd vssd vccd vccd output536/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[2\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[90\] input249/X mprj_logic_high_inst/HI[420] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[90\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input145_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_612_ _612_/A vssd vssd vccd vccd _612_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_24_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input312_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/A vssd vssd vccd vccd _543_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_44_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_474_ _474_/A vssd vssd vccd vccd _474_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_41_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[54\] _518_/Y la_buf\[54\]/TE vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_25_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[126\] input161/X mprj_logic_high_inst/HI[456] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[126\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[110\] _574_/Y la_buf\[110\]/TE vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__einvp_8
XFILLER_29_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[18\] _418_/Y mprj_adr_buf\[18\]/TE vssd vssd vccd vccd mprj_adr_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd vssd vccd vccd output588/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_49_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput380 la_oenb_mprj[93] vssd vssd vccd vccd _356_/A sky130_fd_sc_hd__buf_2
XFILLER_36_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xinput391 mprj_adr_o_core[12] vssd vssd vccd vccd _412_/A sky130_fd_sc_hd__buf_2
XFILLER_1_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] user_to_mprj_in_gates\[43\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_buffers\[8\] user_wb_dat_gates\[8\]/Y vssd vssd vccd vccd output622/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_51_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] user_to_mprj_in_gates\[5\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high_inst/HI[310] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__524__A _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[94\] _357_/Y mprj_logic_high_inst/HI[296] vssd vssd vccd
+ vccd la_oenb_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_46_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input262_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[7\] input237/X mprj_logic_high_inst/HI[337] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[7\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[117\] _380_/A la_buf_enable\[117\]/B vssd vssd vccd vccd la_buf\[117\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_526_ _526_/A vssd vssd vccd vccd _526_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_457_ _457_/A vssd vssd vccd vccd _457_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_388_ _388_/A vssd vssd vccd vccd _388_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__434__A _434_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd vssd vccd vccd output495/A
+ sky130_fd_sc_hd__inv_2
XFILLER_9_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__609__A _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__344__A _344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_49_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[53\] input208/X mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[53\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__519__A _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input108_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[31\] _623_/A la_buf_enable\[31\]/B vssd vssd vccd vccd la_buf\[31\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd vssd vccd vccd output546/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_19_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput19 la_data_out_mprj[113] vssd vssd vccd vccd _577_/A sky130_fd_sc_hd__clkbuf_4
Xla_buf\[17\] _481_/Y la_buf\[17\]/TE vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input73_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_509_ _509_/A vssd vssd vccd vccd _509_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[19\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_53_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[2\]_B la_buf_enable\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[16\] user_wb_dat_gates\[16\]/Y vssd vssd vccd vccd output599/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_5_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] user_to_mprj_in_gates\[117\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__339__A _339_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[127\] _390_/Y mprj_logic_high_inst/HI[329] vssd vssd vccd
+ vccd la_oenb_core[127] sky130_fd_sc_hd__einvp_8
Xoutput470 output470/A vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_2
XFILLER_43_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput481 output481/A vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_2
Xoutput492 output492/A vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_2
XFILLER_47_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[79\] _342_/A la_buf_enable\[79\]/B vssd vssd vccd vccd la_buf\[79\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[57\] _649_/Y mprj_logic_high_inst/HI[259] vssd vssd vccd
+ vccd la_oenb_core[57] sky130_fd_sc_hd__einvp_8
XFILLER_43_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input225_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_A_N _373_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[125\]_A_N _388_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd vssd vccd vccd
+ output479/A sky130_fd_sc_hd__inv_2
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output611_A output611/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd vssd vccd vccd output569/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__622__A _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput209 la_iena_mprj[54] vssd vssd vccd vccd input209/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[16\] input167/X mprj_logic_high_inst/HI[346] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[16\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__532__A _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input175_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input342_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input36_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[84\] _548_/Y la_buf\[84\]/TE vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_1_2237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__442__A _442_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] user_to_mprj_in_gates\[73\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__617__A _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[12\]_A input163/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__352__A _352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__527__A _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_490_ _490_/A vssd vssd vccd vccd _490_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input292_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A _437_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd vssd vccd vccd output528/A
+ sky130_fd_sc_hd__inv_2
XFILLER_34_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__347__A _347_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[83\] input241/X mprj_logic_high_inst/HI[413] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[83\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[61\] _653_/A la_buf_enable\[61\]/B vssd vssd vccd vccd la_buf\[61\]/TE
+ sky130_fd_sc_hd__and2b_1
X_611_ _611_/A vssd vssd vccd vccd _611_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_24_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input138_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_542_ _542_/A vssd vssd vccd vccd _542_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input305_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_473_ _473_/A vssd vssd vccd vccd _473_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[47\] _511_/Y la_buf\[47\]/TE vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__einvp_8
XFILLER_35_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[83\]_A_N _346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[119\] input153/X mprj_logic_high_inst/HI[449] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[119\]/B sky130_fd_sc_hd__and2_1
XFILLER_9_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[90\]_A _554_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[98\]_A_N _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[103\] _567_/Y la_buf\[103\]/TE vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_42_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[21\]_A_N _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput370 la_oenb_mprj[84] vssd vssd vccd vccd _347_/A sky130_fd_sc_hd__buf_4
Xinput381 la_oenb_mprj[94] vssd vssd vccd vccd _357_/A sky130_fd_sc_hd__buf_4
XFILLER_36_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput392 mprj_adr_o_core[13] vssd vssd vccd vccd _413_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[36\]_A_N _628_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] user_to_mprj_in_gates\[36\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[90\]_B la_buf_enable\[90\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__540__A _540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[87\] _350_/Y mprj_logic_high_inst/HI[289] vssd vssd vccd
+ vccd la_oenb_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_29_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input255_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input422_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[31\]_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_525_ _525_/A vssd vssd vccd vccd _525_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[126\]_A _590_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_456_ _456_/A vssd vssd vccd vccd _456_/Y sky130_fd_sc_hd__inv_4
X_387_ _387_/A vssd vssd vccd vccd _387_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[30\] _430_/Y mprj_adr_buf\[30\]/TE vssd vssd vccd vccd mprj_adr_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_output474_A output474/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[81\]_B la_buf_enable\[81\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__450__A _450_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[22\]_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__625__A _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[72\]_B la_buf_enable\[72\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput630 output630/A vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_wb_ena_buf_A input453/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__360__A _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[46\] input200/X mprj_logic_high_inst/HI[376] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[46\]/B sky130_fd_sc_hd__and2_1
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[24\] _616_/A la_buf_enable\[24\]/B vssd vssd vccd vccd la_buf\[24\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__535__A _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input372_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[63\]_B la_buf_enable\[63\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_508_ _508_/A vssd vssd vccd vccd _508_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_output591_A output591/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__445__A _445_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_439_ _439_/A vssd vssd vccd vccd _439_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_6_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[126\]_B mprj_logic_high_inst/HI[456] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__355__A _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[45\]_B la_buf_enable\[45\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput471 output471/A vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_2
Xoutput482 output482/A vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_2
Xoutput493 output493/A vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_2
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[117\]_B mprj_logic_high_inst/HI[447] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input218_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input120_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[1\]/Y sky130_fd_sc_hd__nand2_8
XFILLER_7_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[101\] input134/X mprj_logic_high_inst/HI[431] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[101\]/B sky130_fd_sc_hd__and2_1
XFILLER_32_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[36\]_B la_buf_enable\[36\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[5\]_A input215/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd vssd vccd vccd
+ output471/A sky130_fd_sc_hd__clkinv_4
XFILLER_26_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[108\]_B mprj_logic_high_inst/HI[438] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd vssd vccd vccd output561/A
+ sky130_fd_sc_hd__inv_2
XFILLER_4_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output604_A output604/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[31\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_21_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[27\]_B la_buf_enable\[27\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _438_/Y mprj_dat_buf\[6\]/TE vssd vssd vccd vccd mprj_dat_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[30\]_B mprj_logic_high_inst/HI[360] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[18\]_B la_buf_enable\[18\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input168_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[20\]_A _612_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[91\] _354_/A la_buf_enable\[91\]/B vssd vssd vccd vccd la_buf\[91\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[97\]_B mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input335_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input29_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[77\] _541_/Y la_buf\[77\]/TE vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_35_519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_B mprj_logic_high_inst/HI[351] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[11\]_A _603_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[88\]_B mprj_logic_high_inst/HI[418] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] user_to_mprj_in_gates\[66\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[12\]_B mprj_logic_high_inst/HI[342] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__633__A _633_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[124\]_A_N _387_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__543__A _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input285_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input452_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd vssd vccd vccd output520/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__628__A _628_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[76\] input233/X mprj_logic_high_inst/HI[406] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[76\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[102\] _365_/Y mprj_logic_high_inst/HI[304] vssd vssd vccd
+ vccd la_oenb_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_29_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_610_ _610_/A vssd vssd vccd vccd _610_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__538__A _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ _541_/A vssd vssd vccd vccd _541_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[32\] _624_/Y mprj_logic_high_inst/HI[234] vssd vssd vccd
+ vccd la_oenb_core[32] sky130_fd_sc_hd__einvp_8
XFILLER_2_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[54\] _646_/A la_buf_enable\[54\]/B vssd vssd vccd vccd la_buf\[54\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_472_ _472_/A vssd vssd vccd vccd _472_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input200_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[20\]_A _452_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input96_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput360 la_oenb_mprj[75] vssd vssd vccd vccd _338_/A sky130_fd_sc_hd__buf_2
Xinput371 la_oenb_mprj[85] vssd vssd vccd vccd _348_/A sky130_fd_sc_hd__buf_4
XFILLER_7_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__448__A _448_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput382 la_oenb_mprj[95] vssd vssd vccd vccd _358_/A sky130_fd_sc_hd__clkbuf_4
Xinput393 mprj_adr_o_core[14] vssd vssd vccd vccd _414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] user_to_mprj_in_gates\[29\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_A _429_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__358__A _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[28\] _460_/Y mprj_dat_buf\[28\]/TE vssd vssd vccd vccd mprj_dat_o_user[28]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input150_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input248_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input415_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input11_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[31\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_524_ _524_/A vssd vssd vccd vccd _524_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_455_ _455_/A vssd vssd vccd vccd _455_/Y sky130_fd_sc_hd__inv_6
XFILLER_53_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_386_ _386_/A vssd vssd vccd vccd _386_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[23\] _423_/Y mprj_adr_buf\[23\]/TE vssd vssd vccd vccd mprj_adr_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput190 la_iena_mprj[37] vssd vssd vccd vccd input190/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[8\] _600_/A la_buf_enable\[8\]/B vssd vssd vccd vccd la_buf\[8\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__641__A _641_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput620 output620/A vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_2
XFILLER_43_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_wb_ena_buf_B user_to_mprj_wb_ena_buf/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_A_N _345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[13\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high_inst/HI[278] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[39\] input192/X mprj_logic_high_inst/HI[369] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[39\]/B sky130_fd_sc_hd__and2_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[97\]_A_N _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[17\] _609_/A la_buf_enable\[17\]/B vssd vssd vccd vccd la_buf\[17\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input198_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__551__A _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input365_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[0\] user_irq_core[0] user_irq_gates\[0\]/B vssd vssd vccd vccd user_irq_gates\[0\]/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_input59_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[122\] _385_/A la_buf_enable\[122\]/B vssd vssd vccd vccd la_buf\[122\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_4_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_507_ _507_/A vssd vssd vccd vccd _507_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ _438_/A vssd vssd vccd vccd _438_/Y sky130_fd_sc_hd__inv_2
X_369_ _369_/A vssd vssd vccd vccd _369_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_35_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] user_to_mprj_in_gates\[96\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__636__A _636_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[5\]_A _405_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__371__A _371_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput494 output494/A vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_2
Xoutput472 output472/A vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_2
Xoutput483 output483/A vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_2
XFILLER_47_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input113_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__546__A _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[22\] _486_/Y la_buf\[22\]/TE vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__einvp_8
XFILLER_7_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[5\]_B mprj_logic_high_inst/HI[335] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd vssd vccd vccd output553/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_37_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[24\]/Y sky130_fd_sc_hd__nand2_2
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] user_to_mprj_in_gates\[11\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_2
XFILLER_50_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[21\] user_wb_dat_gates\[21\]/Y vssd vssd vccd vccd output605/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_B la_buf_enable\[126\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] user_to_mprj_in_gates\[122\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__366__A _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[62\] _654_/Y mprj_logic_high_inst/HI[264] vssd vssd vccd
+ vccd la_oenb_core[62] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[84\] _347_/A la_buf_enable\[84\]/B vssd vssd vccd vccd la_buf\[84\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_B la_buf_enable\[117\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[10\] _442_/Y mprj_dat_buf\[10\]/TE vssd vssd vccd vccd mprj_dat_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_input230_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input328_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_buffers\[8\]_A user_wb_dat_gates\[8\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[126\] _590_/Y la_buf\[126\]/TE vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[108\]_B la_buf_enable\[108\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] user_to_mprj_in_gates\[59\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[21\] input173/X mprj_logic_high_inst/HI[351] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[21\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input180_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input41_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input445_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd vssd vccd vccd output512/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_32_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__644__A _644_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[69\] input225/X mprj_logic_high_inst/HI[399] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[69\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_540_ _540_/A vssd vssd vccd vccd _540_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[47\] _639_/A la_buf_enable\[47\]/B vssd vssd vccd vccd la_buf\[47\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[25\] _617_/Y mprj_logic_high_inst/HI[227] vssd vssd vccd
+ vccd la_oenb_core[25] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[7\] _599_/Y mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd la_oenb_core[7] sky130_fd_sc_hd__einvp_8
X_471_ _471_/A vssd vssd vccd vccd _471_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_25_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input395_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input89_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[0\] _464_/Y la_buf\[0\]/TE vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_4_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput361 la_oenb_mprj[76] vssd vssd vccd vccd _339_/A sky130_fd_sc_hd__clkbuf_4
Xinput350 la_oenb_mprj[66] vssd vssd vccd vccd _329_/A sky130_fd_sc_hd__buf_4
Xinput372 la_oenb_mprj[86] vssd vssd vccd vccd _349_/A sky130_fd_sc_hd__buf_4
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput383 la_oenb_mprj[96] vssd vssd vccd vccd _359_/A sky130_fd_sc_hd__clkbuf_2
Xinput394 mprj_adr_o_core[15] vssd vssd vccd vccd _415_/A sky130_fd_sc_hd__buf_2
XFILLER_35_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__464__A _464_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[123\]_A_N _386_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__639__A _639_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__374__A _374_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_1521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input143_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__549__A _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input310_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input408_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_523_ _523_/A vssd vssd vccd vccd _523_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_454_ _454_/A vssd vssd vccd vccd _454_/Y sky130_fd_sc_hd__inv_4
XFILLER_26_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[52\] _516_/Y la_buf\[52\]/TE vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[124\] input159/X mprj_logic_high_inst/HI[454] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[124\]/B sky130_fd_sc_hd__and2_1
XFILLER_53_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_385_ _385_/A vssd vssd vccd vccd _385_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[16\] _416_/Y mprj_adr_buf\[16\]/TE vssd vssd vccd vccd mprj_adr_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output627_A output627/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd vssd vccd vccd output586/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A _459_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_rstn_buf input3/X mprj_rstn_buf/TE vssd vssd vccd vccd user_reset sky130_fd_sc_hd__einvp_8
Xinput180 la_iena_mprj[28] vssd vssd vccd vccd input180/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput191 la_iena_mprj[38] vssd vssd vccd vccd input191/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] user_to_mprj_in_gates\[41\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_buffers\[6\] user_wb_dat_gates\[6\]/Y vssd vssd vccd vccd output620/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_52_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[5\]_B la_buf_enable\[5\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput610 output610/A vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_2
Xoutput621 output621/A vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_2
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] user_to_mprj_in_gates\[3\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_2
XTAP_150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__369__A _369_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high_inst/HI[323] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[92\] _355_/Y mprj_logic_high_inst/HI[294] vssd vssd vccd
+ vccd la_oenb_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input260_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input358_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[5\] input215/X mprj_logic_high_inst/HI[335] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[5\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[115\] _378_/A la_buf_enable\[115\]/B vssd vssd vccd vccd la_buf\[115\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_34_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_506_ _506_/A vssd vssd vccd vccd _506_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_437_ _437_/A vssd vssd vccd vccd _437_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_368_ _368_/A vssd vssd vccd vccd _368_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd vssd vccd vccd output485/A
+ sky130_fd_sc_hd__inv_6
XFILLER_6_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] user_to_mprj_in_gates\[89\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__652__A _652_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput495 output495/A vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_2
Xoutput473 output473/A vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_2
Xoutput484 output484/A vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_2
XFILLER_47_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[51\] input206/X mprj_logic_high_inst/HI[381] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[51\]/B sky130_fd_sc_hd__and2_1
XFILLER_19_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_cyc_buf _393_/Y mprj_cyc_buf/TE vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd vssd vccd vccd output524/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_42_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__562__A _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[119\]_TE la_buf\[119\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[15\] _479_/Y la_buf\[15\]/TE vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_7_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input71_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[8\] _408_/Y mprj_adr_buf\[8\]/TE vssd vssd vccd vccd mprj_adr_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_43_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd vssd vccd vccd output545/A
+ sky130_fd_sc_hd__inv_2
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[17\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[81\]_A_N _344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_buffers\[14\] user_wb_dat_gates\[14\]/Y vssd vssd vccd vccd output597/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high_inst/HI[268] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[96\]_A_N _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] user_to_mprj_in_gates\[115\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA__647__A _647_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[34\]_A_N _626_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__382__A _382_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[49\]_A_N _641_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[99\] input258/X mprj_logic_high_inst/HI[429] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[99\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[125\] _388_/Y mprj_logic_high_inst/HI[327] vssd vssd vccd
+ vccd la_oenb_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_0_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[55\] _647_/Y mprj_logic_high_inst/HI[257] vssd vssd vccd
+ vccd la_oenb_core[55] sky130_fd_sc_hd__einvp_8
XFILLER_25_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[77\] _340_/A la_buf_enable\[77\]/B vssd vssd vccd vccd la_buf\[77\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_input223_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__557__A _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[119\] _583_/Y la_buf\[119\]/TE vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__einvp_8
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd vssd vccd vccd
+ output477/A sky130_fd_sc_hd__clkinv_4
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__467__A _467_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__377__A _377_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[14\] input165/X mprj_logic_high_inst/HI[344] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[14\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input173_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input340_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input438_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input34_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[82\] _546_/Y la_buf\[82\]/TE vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_48_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] user_to_mprj_in_gates\[71\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_1
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_470_ _470_/A vssd vssd vccd vccd _470_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[18\] _610_/Y mprj_logic_high_inst/HI[220] vssd vssd vccd
+ vccd la_oenb_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_25_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input290_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input388_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_B la_buf_enable\[93\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__570__A _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput362 la_oenb_mprj[77] vssd vssd vccd vccd _340_/A sky130_fd_sc_hd__clkbuf_4
Xinput351 la_oenb_mprj[67] vssd vssd vccd vccd _330_/A sky130_fd_sc_hd__buf_4
Xinput340 la_oenb_mprj[57] vssd vssd vccd vccd _649_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput373 la_oenb_mprj[87] vssd vssd vccd vccd _350_/A sky130_fd_sc_hd__clkbuf_4
Xinput384 la_oenb_mprj[97] vssd vssd vccd vccd _360_/A sky130_fd_sc_hd__clkbuf_4
Xinput395 mprj_adr_o_core[16] vssd vssd vccd vccd _416_/A sky130_fd_sc_hd__buf_2
XFILLER_35_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_599_ _599_/A vssd vssd vccd vccd _599_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_43_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd vssd vccd vccd output526/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_34_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[84\]_B la_buf_enable\[84\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__480__A _480_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[25\]_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A _655_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[75\]_B la_buf_enable\[75\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__390__A _390_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[81\] input239/X mprj_logic_high_inst/HI[411] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[81\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[16\]_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input136_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_522_ _522_/A vssd vssd vccd vccd _522_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input303_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__565__A _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_453_ _453_/A vssd vssd vccd vccd _453_/Y sky130_fd_sc_hd__inv_4
XFILLER_26_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_384_ _384_/A vssd vssd vccd vccd _384_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf\[45\] _509_/Y la_buf\[45\]/TE vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__einvp_8
XFILLER_51_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[117\] input151/X mprj_logic_high_inst/HI[447] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[117\]/B sky130_fd_sc_hd__and2_1
XFILLER_51_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[66\]_B la_buf_enable\[66\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[101\] _565_/Y la_buf\[101\]/TE vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_9_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput170 la_iena_mprj[19] vssd vssd vccd vccd input170/X sky130_fd_sc_hd__clkbuf_1
Xinput181 la_iena_mprj[29] vssd vssd vccd vccd input181/X sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd vssd vccd vccd output578/A
+ sky130_fd_sc_hd__clkinv_4
Xinput192 la_iena_mprj[39] vssd vssd vccd vccd input192/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__475__A _475_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] user_to_mprj_in_gates\[34\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput600 output600/A vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_2
Xoutput611 output611/A vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_2
Xoutput622 output622/A vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_2
XFILLER_47_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__385__A _385_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[85\] _348_/Y mprj_logic_high_inst/HI[287] vssd vssd vccd
+ vccd la_oenb_core[85] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[50\]_A _642_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input253_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input420_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[108\] _371_/A la_buf_enable\[108\]/B vssd vssd vccd vccd la_buf\[108\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_505_ _505_/A vssd vssd vccd vccd _505_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[51\]_B mprj_logic_high_inst/HI[381] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[122\]_A_N _385_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_436_ _436_/A vssd vssd vccd vccd _436_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_367_ _367_/A vssd vssd vccd vccd _367_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[8\]_A input248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[41\]_A _633_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[42\]_B mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_A _624_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput463 output463/A vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_2
Xoutput474 output474/A vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_2
Xoutput485 output485/A vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_2
Xoutput496 output496/A vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_2
XFILLER_47_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[44\] input198/X mprj_logic_high_inst/HI[374] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[44\]/B sky130_fd_sc_hd__and2_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[33\]_B mprj_logic_high_inst/HI[363] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[22\] _614_/A la_buf_enable\[22\]/B vssd vssd vccd vccd la_buf\[22\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_23_460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input370_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_A _615_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input64_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[24\]_B mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_419_ _419_/A vssd vssd vccd vccd _419_/Y sky130_fd_sc_hd__inv_16
XFILLER_14_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _606_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] user_to_mprj_in_gates\[108\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_A _410_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[15\]_B mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[8\]_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _381_/Y mprj_logic_high_inst/HI[320] vssd vssd vccd
+ vccd la_oenb_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_25_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[48\] _640_/Y mprj_logic_high_inst/HI[250] vssd vssd vccd
+ vccd la_oenb_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_47_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[2\]_B user_irq_ena_buf\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input216_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__573__A _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd vssd vccd vccd
+ output469/A sky130_fd_sc_hd__inv_2
XFILLER_43_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd vssd vccd vccd output559/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output602_A output602/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[4\] _436_/Y mprj_dat_buf\[4\]/TE vssd vssd vccd vccd mprj_dat_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input166_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__568__A _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input333_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[80\]_A_N _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input27_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[75\] _539_/Y la_buf\[75\]/TE vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[23\]_A _455_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[56\]_TE mprj_logic_high_inst/HI[258] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[95\]_A_N _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[33\]_A_N _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[48\]_A_N _640_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] user_to_mprj_in_gates\[64\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[14\]_A _446_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__388__A _388_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high_inst/HI[281] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[9\]_A _601_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[12\]_A user_wb_dat_gates\[12\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input283_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput330 la_oenb_mprj[48] vssd vssd vccd vccd _640_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput352 la_oenb_mprj[68] vssd vssd vccd vccd _331_/A sky130_fd_sc_hd__clkbuf_2
Xinput341 la_oenb_mprj[58] vssd vssd vccd vccd _650_/A sky130_fd_sc_hd__buf_2
Xinput363 la_oenb_mprj[78] vssd vssd vccd vccd _341_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput374 la_oenb_mprj[88] vssd vssd vccd vccd _351_/A sky130_fd_sc_hd__buf_4
Xinput385 la_oenb_mprj[98] vssd vssd vccd vccd _361_/A sky130_fd_sc_hd__clkbuf_4
Xinput396 mprj_adr_o_core[17] vssd vssd vccd vccd _417_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_598_ _598_/A vssd vssd vccd vccd _598_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd vssd vccd vccd output518/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_8_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[25\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[74\] input231/X mprj_logic_high_inst/HI[404] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[74\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[100\] _363_/Y mprj_logic_high_inst/HI[302] vssd vssd vccd
+ vccd la_oenb_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_24_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[16\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[30\] _622_/Y mprj_logic_high_inst/HI[232] vssd vssd vccd
+ vccd la_oenb_core[30] sky130_fd_sc_hd__einvp_8
XFILLER_2_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input129_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[52\] _644_/A la_buf_enable\[52\]/B vssd vssd vccd vccd la_buf\[52\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_521_ _521_/A vssd vssd vccd vccd _521_/Y sky130_fd_sc_hd__inv_2
X_452_ _452_/A vssd vssd vccd vccd _452_/Y sky130_fd_sc_hd__inv_4
X_383_ _383_/A vssd vssd vccd vccd _383_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__581__A _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input94_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[38\] _502_/Y la_buf\[38\]/TE vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_51_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput171 la_iena_mprj[1] vssd vssd vccd vccd input171/X sky130_fd_sc_hd__clkbuf_1
Xinput160 la_iena_mprj[125] vssd vssd vccd vccd input160/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput193 la_iena_mprj[3] vssd vssd vccd vccd input193/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput182 la_iena_mprj[2] vssd vssd vccd vccd input182/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] user_to_mprj_in_gates\[27\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput601 output601/A vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_2
Xoutput623 output623/A vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_2
Xoutput612 output612/A vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_2
XFILLER_47_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[8\]_A _408_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[78\] _341_/Y mprj_logic_high_inst/HI[280] vssd vssd vccd
+ vccd la_oenb_core[78] sky130_fd_sc_hd__einvp_8
XFILLER_2_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[26\] _458_/Y mprj_dat_buf\[26\]/TE vssd vssd vccd vccd mprj_dat_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input246_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input413_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__576__A _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_504_ _504_/A vssd vssd vccd vccd _504_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_435_ _435_/A vssd vssd vccd vccd _435_/Y sky130_fd_sc_hd__inv_2
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_366_ _366_/A vssd vssd vccd vccd _366_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[8\]_B mprj_logic_high_inst/HI[338] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[21\] _421_/Y mprj_adr_buf\[21\]/TE vssd vssd vccd vccd mprj_adr_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__486__A _486_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[6\] _598_/A la_buf_enable\[6\]/B vssd vssd vccd vccd la_buf\[6\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput464 output464/A vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_2
Xoutput475 output475/A vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_2
Xoutput486 output486/A vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_2
Xoutput497 output497/A vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_2
XFILLER_25_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[37\] input190/X mprj_logic_high_inst/HI[367] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[37\]/B sky130_fd_sc_hd__and2_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[15\] _607_/A la_buf_enable\[15\]/B vssd vssd vccd vccd la_buf\[15\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input196_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input363_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input57_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[120\] _383_/A la_buf_enable\[120\]/B vssd vssd vccd vccd la_buf\[120\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_418_ _418_/A vssd vssd vccd vccd _418_/Y sky130_fd_sc_hd__inv_12
XFILLER_14_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_349_ _349_/A vssd vssd vccd vccd _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] user_to_mprj_in_gates\[94\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[8\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[121\]_A_N _384_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input209_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input111_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[20\] _484_/Y la_buf\[20\]/TE vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__einvp_8
XFILLER_11_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd vssd vccd vccd output551/A
+ sky130_fd_sc_hd__inv_2
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[22\]/Y sky130_fd_sc_hd__nand2_2
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] user_to_mprj_in_gates\[120\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[60\] _652_/Y mprj_logic_high_inst/HI[262] vssd vssd vccd
+ vccd la_oenb_core[60] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[82\] _345_/A la_buf_enable\[82\]/B vssd vssd vccd vccd la_buf\[82\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_input159_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input326_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__584__A _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[68\] _532_/Y la_buf\[68\]/TE vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__einvp_8
XFILLER_51_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[124\] _588_/Y la_buf\[124\]/TE vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_12_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] user_to_mprj_in_gates\[57\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__494__A _494_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_50_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input276_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__579__A _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input443_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput320 la_oenb_mprj[39] vssd vssd vccd vccd _631_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high_inst/HI[225] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xinput353 la_oenb_mprj[69] vssd vssd vccd vccd _332_/A sky130_fd_sc_hd__clkbuf_2
Xinput342 la_oenb_mprj[59] vssd vssd vccd vccd _651_/A sky130_fd_sc_hd__clkbuf_2
Xinput331 la_oenb_mprj[49] vssd vssd vccd vccd _641_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput364 la_oenb_mprj[79] vssd vssd vccd vccd _342_/A sky130_fd_sc_hd__clkbuf_4
Xinput375 la_oenb_mprj[89] vssd vssd vccd vccd _352_/A sky130_fd_sc_hd__buf_4
Xinput386 la_oenb_mprj[99] vssd vssd vccd vccd _362_/A sky130_fd_sc_hd__clkbuf_4
Xinput397 mprj_adr_o_core[18] vssd vssd vccd vccd _418_/A sky130_fd_sc_hd__buf_2
XFILLER_48_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_597_ _597_/A vssd vssd vccd vccd _597_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd vssd vccd vccd output510/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_51_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__489__A _489_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[8\]_B la_buf_enable\[8\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[94\]_A_N _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[67\] input223/X mprj_logic_high_inst/HI[397] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[67\]/B sky130_fd_sc_hd__and2_1
XFILLER_46_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_520_ _520_/A vssd vssd vccd vccd _520_/Y sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_oen_buffers\[5\] _597_/Y mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd la_oenb_core[5] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[23\] _615_/Y mprj_logic_high_inst/HI[225] vssd vssd vccd
+ vccd la_oenb_core[23] sky130_fd_sc_hd__einvp_8
X_451_ _451_/A vssd vssd vccd vccd _451_/Y sky130_fd_sc_hd__inv_4
XFILLER_32_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[45\] _637_/A la_buf_enable\[45\]/B vssd vssd vccd vccd la_buf\[45\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_382_ _382_/A vssd vssd vccd vccd _382_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[32\]_A_N _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input393_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[47\]_A_N _639_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input87_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput172 la_iena_mprj[20] vssd vssd vccd vccd input172/X sky130_fd_sc_hd__clkbuf_1
Xinput150 la_iena_mprj[116] vssd vssd vccd vccd input150/X sky130_fd_sc_hd__clkbuf_1
Xinput161 la_iena_mprj[126] vssd vssd vccd vccd input161/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput194 la_iena_mprj[40] vssd vssd vccd vccd input194/X sky130_fd_sc_hd__clkbuf_1
Xinput183 la_iena_mprj[30] vssd vssd vccd vccd input183/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_649_ _649_/A vssd vssd vccd vccd _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high_inst/HI[271] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput602 output602/A vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_2
Xoutput613 output613/A vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_2
Xoutput624 output624/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_2
XFILLER_47_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[19\] _451_/Y mprj_dat_buf\[19\]/TE vssd vssd vccd vccd mprj_dat_o_user[19]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input239_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input141_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input406_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_503_ _503_/A vssd vssd vccd vccd _503_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_434_ _434_/A vssd vssd vccd vccd _434_/Y sky130_fd_sc_hd__inv_2
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[50\] _514_/Y la_buf\[50\]/TE vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__einvp_8
XANTENNA__592__A _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_365_ _365_/A vssd vssd vccd vccd _365_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[122\] input157/X mprj_logic_high_inst/HI[452] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[122\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[3\]_A _435_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[14\] _414_/Y mprj_adr_buf\[14\]/TE vssd vssd vccd vccd mprj_adr_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_42_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd vssd vccd vccd output584/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_output625_A output625/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[4\] user_wb_dat_gates\[4\]/Y vssd vssd vccd vccd output618/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_51_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] user_to_mprj_in_gates\[1\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_1
Xoutput465 output465/A vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_2
Xoutput476 output476/A vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_2
Xoutput487 output487/A vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_2
Xoutput498 output498/A vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_2
XFILLER_25_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input189_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[90\] _353_/Y mprj_logic_high_inst/HI[292] vssd vssd vccd
+ vccd la_oenb_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_2_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input356_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[98\] _562_/Y la_buf\[98\]/TE vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[3\] input193/X mprj_logic_high_inst/HI[333] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[3\]/B sky130_fd_sc_hd__and2_1
XANTENNA__587__A _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[113\] _376_/A la_buf_enable\[113\]/B vssd vssd vccd vccd la_buf\[113\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_417_ _417_/A vssd vssd vccd vccd _417_/Y sky130_fd_sc_hd__inv_6
X_348_ _348_/A vssd vssd vccd vccd _348_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] user_to_mprj_in_gates\[87\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__497__A _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input104_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd vssd vccd vccd output502/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_23_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[13\] _477_/Y la_buf\[13\]/TE vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__einvp_8
XFILLER_32_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[9\] _473_/Y la_buf\[9\]/TE vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_48_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[6\] _406_/Y mprj_adr_buf\[6\]/TE vssd vssd vccd vccd mprj_adr_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_47_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd vssd vccd vccd output543/A
+ sky130_fd_sc_hd__clkinv_4
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] user_wb_ack_gate/B vssd vssd vccd vccd
+ user_wb_dat_gates\[15\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[12\] user_wb_dat_gates\[12\]/Y vssd vssd vccd vccd output595/A
+ sky130_fd_sc_hd__clkinv_8
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] user_to_mprj_in_gates\[113\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[110\]_B mprj_logic_high_inst/HI[440] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[97\] input256/X mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[97\]/B sky130_fd_sc_hd__and2_1
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[123\] _386_/Y mprj_logic_high_inst/HI[325] vssd vssd vccd
+ vccd la_oenb_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_27_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[53\] _645_/Y mprj_logic_high_inst/HI[255] vssd vssd vccd
+ vccd la_oenb_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_0_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[75\] _338_/A la_buf_enable\[75\]/B vssd vssd vccd vccd la_buf\[75\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input221_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input319_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[101\]_B mprj_logic_high_inst/HI[431] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[96\]_B la_buf_enable\[96\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[117\] _581_/Y la_buf\[117\]/TE vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_4_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd vssd vccd vccd
+ output475/A sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[20\]_B la_buf_enable\[20\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[120\]_A_N _383_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[87\]_B la_buf_enable\[87\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[28\]_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_B la_buf_enable\[11\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[90\]_B mprj_logic_high_inst/HI[420] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_53_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[12\] input163/X mprj_logic_high_inst/HI[342] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[12\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[78\]_B la_buf_enable\[78\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input171_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input269_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[19\]_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput321 la_oenb_mprj[3] vssd vssd vccd vccd _595_/A sky130_fd_sc_hd__clkbuf_2
Xinput310 la_oenb_mprj[2] vssd vssd vccd vccd _594_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input436_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput354 la_oenb_mprj[6] vssd vssd vccd vccd _598_/A sky130_fd_sc_hd__clkbuf_2
Xinput343 la_oenb_mprj[5] vssd vssd vccd vccd _597_/A sky130_fd_sc_hd__buf_2
Xinput332 la_oenb_mprj[4] vssd vssd vccd vccd _596_/A sky130_fd_sc_hd__buf_2
XANTENNA_input32_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[80\] _544_/Y la_buf\[80\]/TE vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__einvp_8
Xinput387 la_oenb_mprj[9] vssd vssd vccd vccd _601_/A sky130_fd_sc_hd__clkbuf_2
Xinput376 la_oenb_mprj[8] vssd vssd vccd vccd _600_/A sky130_fd_sc_hd__buf_2
Xinput365 la_oenb_mprj[7] vssd vssd vccd vccd _599_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__595__A _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput398 mprj_adr_o_core[19] vssd vssd vccd vccd _419_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_596_ _596_/A vssd vssd vccd vccd _596_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[69\]_B la_buf_enable\[69\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_450_ _450_/A vssd vssd vccd vccd _450_/Y sky130_fd_sc_hd__inv_4
Xuser_to_mprj_oen_buffers\[16\] _608_/Y mprj_logic_high_inst/HI[218] vssd vssd vccd
+ vccd la_oenb_core[16] sky130_fd_sc_hd__einvp_8
X_381_ _381_/A vssd vssd vccd vccd _381_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[38\] _630_/A la_buf_enable\[38\]/B vssd vssd vccd vccd la_buf\[38\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_40_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input386_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput140 la_iena_mprj[107] vssd vssd vccd vccd input140/X sky130_fd_sc_hd__clkbuf_1
Xinput151 la_iena_mprj[117] vssd vssd vccd vccd input151/X sky130_fd_sc_hd__clkbuf_1
Xinput162 la_iena_mprj[127] vssd vssd vccd vccd input162/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput195 la_iena_mprj[41] vssd vssd vccd vccd input195/X sky130_fd_sc_hd__clkbuf_1
Xinput173 la_iena_mprj[21] vssd vssd vccd vccd input173/X sky130_fd_sc_hd__clkbuf_1
Xinput184 la_iena_mprj[31] vssd vssd vccd vccd input184/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_user_to_mprj_in_ena_buf\[54\]_B mprj_logic_high_inst/HI[384] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_648_ _648_/A vssd vssd vccd vccd _648_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_36_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_579_ _579_/A vssd vssd vccd vccd _579_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_53_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high_inst/HI[316] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[44\]_A _636_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput614 output614/A vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_2
Xoutput603 output603/A vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_2
Xoutput625 output625/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_2
XFILLER_47_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[45\]_B mprj_logic_high_inst/HI[375] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_A _627_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_A _431_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input134_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[36\]_B mprj_logic_high_inst/HI[366] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_input301_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_502_ _502_/A vssd vssd vccd vccd _502_/Y sky130_fd_sc_hd__inv_2
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _433_/A vssd vssd vccd vccd _433_/Y sky130_fd_sc_hd__inv_2
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_364_ _364_/A vssd vssd vccd vccd _364_/Y sky130_fd_sc_hd__clkinv_2
Xla_buf\[43\] _507_/Y la_buf\[43\]/TE vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[115\] input149/X mprj_logic_high_inst/HI[445] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[115\]/B sky130_fd_sc_hd__and2_1
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[26\]_A _618_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output618_A output618/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd vssd vccd vccd output576/A
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_adr_buf\[22\]_A _422_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[27\]_B mprj_logic_high_inst/HI[357] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_51_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] user_to_mprj_in_gates\[32\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_A_N _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[17\]_A _609_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_A_N _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput466 output466/A vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_2
Xoutput477 output477/A vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_2
Xoutput499 output499/A vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_2
Xoutput488 output488/A vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_2
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_A _413_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[46\]_A_N _638_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_B mprj_logic_high_inst/HI[348] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[83\] _346_/Y mprj_logic_high_inst/HI[285] vssd vssd vccd
+ vccd la_oenb_core[83] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[31\] _463_/Y mprj_dat_buf\[31\]/TE vssd vssd vccd vccd mprj_dat_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input349_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input251_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[106\] _369_/A la_buf_enable\[106\]/B vssd vssd vccd vccd la_buf\[106\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_416_ _416_/A vssd vssd vccd vccd _416_/Y sky130_fd_sc_hd__inv_12
X_347_ _347_/A vssd vssd vccd vccd _347_/Y sky130_fd_sc_hd__inv_2
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[97\]_TE la_buf\[97\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[42\] input196/X mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd user_to_mprj_in_gates\[42\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[20\] _612_/A la_buf_enable\[20\]/B vssd vssd vccd vccd la_buf\[20\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_input299_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input62_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__598__A _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[26\]_A _458_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[17\]_A _449_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] user_to_mprj_in_gates\[106\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[116\] _379_/Y mprj_logic_high_inst/HI[318] vssd vssd vccd
+ vccd la_oenb_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_5_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _638_/Y mprj_logic_high_inst/HI[248] vssd vssd vccd
+ vccd la_oenb_core[46] sky130_fd_sc_hd__einvp_8
XFILLER_47_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[68\] _331_/A la_buf_enable\[68\]/B vssd vssd vccd vccd la_buf\[68\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input214_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[15\]_A user_wb_dat_gates\[15\]/Y vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_5_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd vssd vccd vccd
+ output467/A sky130_fd_sc_hd__inv_2
XFILLER_43_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[28\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[2\] _434_/Y mprj_dat_buf\[2\]/TE vssd vssd vccd vccd mprj_dat_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_26_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_B la_buf_enable\[110\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_buffers\[1\]_A user_wb_dat_gates\[1\]/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input164_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[19\]_B user_wb_ack_gate/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput300 la_oenb_mprj[20] vssd vssd vccd vccd _612_/A sky130_fd_sc_hd__clkbuf_2
Xinput311 la_oenb_mprj[30] vssd vssd vccd vccd _622_/A sky130_fd_sc_hd__buf_2
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput344 la_oenb_mprj[60] vssd vssd vccd vccd _652_/A sky130_fd_sc_hd__buf_2
Xinput333 la_oenb_mprj[50] vssd vssd vccd vccd _642_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input331_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput322 la_oenb_mprj[40] vssd vssd vccd vccd _632_/A sky130_fd_sc_hd__buf_4
XANTENNA_input429_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput355 la_oenb_mprj[70] vssd vssd vccd vccd _333_/A sky130_fd_sc_hd__buf_2
Xinput366 la_oenb_mprj[80] vssd vssd vccd vccd _343_/A sky130_fd_sc_hd__clkbuf_4
Xinput377 la_oenb_mprj[90] vssd vssd vccd vccd _353_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input25_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput388 mprj_adr_o_core[0] vssd vssd vccd vccd _400_/A sky130_fd_sc_hd__buf_12
Xinput399 mprj_adr_o_core[1] vssd vssd vccd vccd _401_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[73\] _537_/Y la_buf\[73\]/TE vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__einvp_8
XFILLER_28_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[101\]_B la_buf_enable\[101\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_595_ _595_/A vssd vssd vccd vccd _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] user_to_mprj_in_gates\[62\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_380_ _380_/A vssd vssd vccd vccd _380_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input281_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_74 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input379_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput163 la_iena_mprj[12] vssd vssd vccd vccd input163/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput130 la_data_out_mprj[99] vssd vssd vccd vccd _563_/A sky130_fd_sc_hd__clkbuf_2
Xinput141 la_iena_mprj[108] vssd vssd vccd vccd input141/X sky130_fd_sc_hd__clkbuf_1
Xinput152 la_iena_mprj[118] vssd vssd vccd vccd input152/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xinput196 la_iena_mprj[42] vssd vssd vccd vccd input196/X sky130_fd_sc_hd__clkbuf_1
Xinput174 la_iena_mprj[22] vssd vssd vccd vccd input174/X sky130_fd_sc_hd__clkbuf_1
Xinput185 la_iena_mprj[32] vssd vssd vccd vccd input185/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_647_ _647_/A vssd vssd vccd vccd _647_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_578_ _578_/A vssd vssd vccd vccd _578_/Y sky130_fd_sc_hd__inv_4
XFILLER_17_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd vssd vccd vccd output516/A
+ sky130_fd_sc_hd__clkinv_4
XFILLER_12_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xoutput604 output604/A vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_2
Xoutput615 output615/A vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_2
Xoutput626 output626/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

