magic
tech sky130A
magscale 1 2
timestamp 1677512548
<< obsli1 >>
rect 1012 1071 7912 8721
<< obsm1 >>
rect 290 960 8634 9444
<< metal2 >>
rect 754 9200 810 10000
rect 1030 9200 1086 10000
rect 1306 9200 1362 10000
rect 1582 9200 1638 10000
rect 1858 9200 1914 10000
rect 2134 9200 2190 10000
rect 2410 9200 2466 10000
rect 2686 9200 2742 10000
rect 2962 9200 3018 10000
rect 3238 9200 3294 10000
rect 3514 9200 3570 10000
rect 3790 9200 3846 10000
rect 4066 9200 4122 10000
rect 4342 9200 4398 10000
rect 4618 9200 4674 10000
rect 4894 9200 4950 10000
rect 5170 9200 5226 10000
rect 5446 9200 5502 10000
rect 5722 9200 5778 10000
rect 5998 9200 6054 10000
rect 6274 9200 6330 10000
rect 6550 9200 6606 10000
rect 6826 9200 6882 10000
rect 7102 9200 7158 10000
rect 7378 9200 7434 10000
rect 7654 9200 7710 10000
rect 7930 9200 7986 10000
rect 8206 9200 8262 10000
rect 294 0 350 800
rect 754 0 810 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
<< obsm2 >>
rect 296 9144 698 9466
rect 866 9144 974 9466
rect 1142 9144 1250 9466
rect 1418 9144 1526 9466
rect 1694 9144 1802 9466
rect 1970 9144 2078 9466
rect 2246 9144 2354 9466
rect 2522 9144 2630 9466
rect 2798 9144 2906 9466
rect 3074 9144 3182 9466
rect 3350 9144 3458 9466
rect 3626 9144 3734 9466
rect 3902 9144 4010 9466
rect 4178 9144 4286 9466
rect 4454 9144 4562 9466
rect 4730 9144 4838 9466
rect 5006 9144 5114 9466
rect 5282 9144 5390 9466
rect 5558 9144 5666 9466
rect 5834 9144 5942 9466
rect 6110 9144 6218 9466
rect 6386 9144 6494 9466
rect 6662 9144 6770 9466
rect 6938 9144 7046 9466
rect 7214 9144 7322 9466
rect 7490 9144 7598 9466
rect 7766 9144 7874 9466
rect 8042 9144 8150 9466
rect 8318 9144 8628 9466
rect 296 856 8628 9144
rect 406 575 698 856
rect 866 575 1158 856
rect 1326 575 1618 856
rect 1786 575 2078 856
rect 2246 575 2538 856
rect 2706 575 2998 856
rect 3166 575 3458 856
rect 3626 575 3918 856
rect 4086 575 4378 856
rect 4546 575 4838 856
rect 5006 575 5298 856
rect 5466 575 5758 856
rect 5926 575 6218 856
rect 6386 575 6678 856
rect 6846 575 7138 856
rect 7306 575 7598 856
rect 7766 575 8058 856
rect 8226 575 8518 856
<< metal3 >>
rect 0 8984 800 9104
rect 8200 9120 9000 9240
rect 8200 8712 9000 8832
rect 0 8304 800 8424
rect 8200 8304 9000 8424
rect 8200 7896 9000 8016
rect 0 7624 800 7744
rect 8200 7488 9000 7608
rect 0 6944 800 7064
rect 8200 7080 9000 7200
rect 8200 6672 9000 6792
rect 0 6264 800 6384
rect 8200 6264 9000 6384
rect 8200 5856 9000 5976
rect 0 5584 800 5704
rect 8200 5448 9000 5568
rect 0 4904 800 5024
rect 8200 5040 9000 5160
rect 8200 4632 9000 4752
rect 0 4224 800 4344
rect 8200 4224 9000 4344
rect 8200 3816 9000 3936
rect 0 3544 800 3664
rect 8200 3408 9000 3528
rect 0 2864 800 2984
rect 8200 3000 9000 3120
rect 8200 2592 9000 2712
rect 0 2184 800 2304
rect 8200 2184 9000 2304
rect 8200 1776 9000 1896
rect 0 1504 800 1624
rect 8200 1368 9000 1488
rect 0 824 800 944
rect 8200 960 9000 1080
rect 8200 552 9000 672
<< obsm3 >>
rect 800 9184 8120 9212
rect 880 9040 8120 9184
rect 880 8912 8218 9040
rect 880 8904 8120 8912
rect 800 8632 8120 8904
rect 800 8504 8218 8632
rect 880 8224 8120 8504
rect 800 8096 8218 8224
rect 800 7824 8120 8096
rect 880 7816 8120 7824
rect 880 7688 8218 7816
rect 880 7544 8120 7688
rect 800 7408 8120 7544
rect 800 7280 8218 7408
rect 800 7144 8120 7280
rect 880 7000 8120 7144
rect 880 6872 8218 7000
rect 880 6864 8120 6872
rect 800 6592 8120 6864
rect 800 6464 8218 6592
rect 880 6184 8120 6464
rect 800 6056 8218 6184
rect 800 5784 8120 6056
rect 880 5776 8120 5784
rect 880 5648 8218 5776
rect 880 5504 8120 5648
rect 800 5368 8120 5504
rect 800 5240 8218 5368
rect 800 5104 8120 5240
rect 880 4960 8120 5104
rect 880 4832 8218 4960
rect 880 4824 8120 4832
rect 800 4552 8120 4824
rect 800 4424 8218 4552
rect 880 4144 8120 4424
rect 800 4016 8218 4144
rect 800 3744 8120 4016
rect 880 3736 8120 3744
rect 880 3608 8218 3736
rect 880 3464 8120 3608
rect 800 3328 8120 3464
rect 800 3200 8218 3328
rect 800 3064 8120 3200
rect 880 2920 8120 3064
rect 880 2792 8218 2920
rect 880 2784 8120 2792
rect 800 2512 8120 2784
rect 800 2384 8218 2512
rect 880 2104 8120 2384
rect 800 1976 8218 2104
rect 800 1704 8120 1976
rect 880 1696 8120 1704
rect 880 1568 8218 1696
rect 880 1424 8120 1568
rect 800 1288 8120 1424
rect 800 1160 8218 1288
rect 800 1024 8120 1160
rect 880 880 8120 1024
rect 880 752 8218 880
rect 880 744 8120 752
rect 800 579 8120 744
<< metal4 >>
rect 1714 1040 2034 8752
rect 2576 1040 2896 8752
rect 3439 1040 3759 8752
rect 4301 1040 4621 8752
rect 5164 1040 5484 8752
rect 6026 1040 6346 8752
rect 6889 1040 7209 8752
rect 7751 1040 8071 8752
<< obsm4 >>
rect 4107 8832 5645 9213
rect 4107 3027 4221 8832
rect 4701 3027 5084 8832
rect 5564 3027 5645 8832
<< labels >>
rlabel metal4 s 2576 1040 2896 8752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4301 1040 4621 8752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6026 1040 6346 8752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7751 1040 8071 8752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1714 1040 2034 8752 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3439 1040 3759 8752 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5164 1040 5484 8752 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6889 1040 7209 8752 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 7930 9200 7986 10000 6 mgmt_gpio_in[0]
port 3 nsew signal input
rlabel metal2 s 2410 9200 2466 10000 6 mgmt_gpio_in[10]
port 4 nsew signal input
rlabel metal2 s 1858 9200 1914 10000 6 mgmt_gpio_in[11]
port 5 nsew signal input
rlabel metal2 s 1306 9200 1362 10000 6 mgmt_gpio_in[12]
port 6 nsew signal input
rlabel metal2 s 754 9200 810 10000 6 mgmt_gpio_in[13]
port 7 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 mgmt_gpio_in[14]
port 8 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 mgmt_gpio_in[15]
port 9 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 mgmt_gpio_in[16]
port 10 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 mgmt_gpio_in[17]
port 11 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 mgmt_gpio_in[18]
port 12 nsew signal input
rlabel metal2 s 7378 9200 7434 10000 6 mgmt_gpio_in[1]
port 13 nsew signal input
rlabel metal2 s 6826 9200 6882 10000 6 mgmt_gpio_in[2]
port 14 nsew signal input
rlabel metal2 s 6274 9200 6330 10000 6 mgmt_gpio_in[3]
port 15 nsew signal input
rlabel metal2 s 5722 9200 5778 10000 6 mgmt_gpio_in[4]
port 16 nsew signal input
rlabel metal2 s 5170 9200 5226 10000 6 mgmt_gpio_in[5]
port 17 nsew signal input
rlabel metal2 s 4618 9200 4674 10000 6 mgmt_gpio_in[6]
port 18 nsew signal input
rlabel metal2 s 4066 9200 4122 10000 6 mgmt_gpio_in[7]
port 19 nsew signal input
rlabel metal2 s 3514 9200 3570 10000 6 mgmt_gpio_in[8]
port 20 nsew signal input
rlabel metal2 s 2962 9200 3018 10000 6 mgmt_gpio_in[9]
port 21 nsew signal input
rlabel metal3 s 8200 1776 9000 1896 6 mgmt_gpio_in_buf[0]
port 22 nsew signal output
rlabel metal3 s 8200 5856 9000 5976 6 mgmt_gpio_in_buf[10]
port 23 nsew signal output
rlabel metal3 s 8200 6264 9000 6384 6 mgmt_gpio_in_buf[11]
port 24 nsew signal output
rlabel metal3 s 8200 6672 9000 6792 6 mgmt_gpio_in_buf[12]
port 25 nsew signal output
rlabel metal3 s 8200 7080 9000 7200 6 mgmt_gpio_in_buf[13]
port 26 nsew signal output
rlabel metal3 s 8200 7488 9000 7608 6 mgmt_gpio_in_buf[14]
port 27 nsew signal output
rlabel metal3 s 8200 7896 9000 8016 6 mgmt_gpio_in_buf[15]
port 28 nsew signal output
rlabel metal3 s 8200 8304 9000 8424 6 mgmt_gpio_in_buf[16]
port 29 nsew signal output
rlabel metal3 s 8200 8712 9000 8832 6 mgmt_gpio_in_buf[17]
port 30 nsew signal output
rlabel metal3 s 8200 9120 9000 9240 6 mgmt_gpio_in_buf[18]
port 31 nsew signal output
rlabel metal3 s 8200 2184 9000 2304 6 mgmt_gpio_in_buf[1]
port 32 nsew signal output
rlabel metal3 s 8200 2592 9000 2712 6 mgmt_gpio_in_buf[2]
port 33 nsew signal output
rlabel metal3 s 8200 3000 9000 3120 6 mgmt_gpio_in_buf[3]
port 34 nsew signal output
rlabel metal3 s 8200 3408 9000 3528 6 mgmt_gpio_in_buf[4]
port 35 nsew signal output
rlabel metal3 s 8200 3816 9000 3936 6 mgmt_gpio_in_buf[5]
port 36 nsew signal output
rlabel metal3 s 8200 4224 9000 4344 6 mgmt_gpio_in_buf[6]
port 37 nsew signal output
rlabel metal3 s 8200 4632 9000 4752 6 mgmt_gpio_in_buf[7]
port 38 nsew signal output
rlabel metal3 s 8200 5040 9000 5160 6 mgmt_gpio_in_buf[8]
port 39 nsew signal output
rlabel metal3 s 8200 5448 9000 5568 6 mgmt_gpio_in_buf[9]
port 40 nsew signal output
rlabel metal3 s 8200 552 9000 672 6 mgmt_gpio_oeb[0]
port 41 nsew signal input
rlabel metal3 s 8200 960 9000 1080 6 mgmt_gpio_oeb[1]
port 42 nsew signal input
rlabel metal3 s 8200 1368 9000 1488 6 mgmt_gpio_oeb[2]
port 43 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 mgmt_gpio_oeb_buf[0]
port 44 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 mgmt_gpio_oeb_buf[1]
port 45 nsew signal output
rlabel metal3 s 0 824 800 944 6 mgmt_gpio_oeb_buf[2]
port 46 nsew signal output
rlabel metal2 s 294 0 350 800 6 mgmt_gpio_out[0]
port 47 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 mgmt_gpio_out[10]
port 48 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 mgmt_gpio_out[11]
port 49 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 mgmt_gpio_out[12]
port 50 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 mgmt_gpio_out[13]
port 51 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 mgmt_gpio_out[14]
port 52 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 mgmt_gpio_out[15]
port 53 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 mgmt_gpio_out[16]
port 54 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 mgmt_gpio_out[17]
port 55 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 mgmt_gpio_out[18]
port 56 nsew signal input
rlabel metal2 s 754 0 810 800 6 mgmt_gpio_out[1]
port 57 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 mgmt_gpio_out[2]
port 58 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 mgmt_gpio_out[3]
port 59 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 mgmt_gpio_out[4]
port 60 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 mgmt_gpio_out[5]
port 61 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 mgmt_gpio_out[6]
port 62 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 mgmt_gpio_out[7]
port 63 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 mgmt_gpio_out[8]
port 64 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 mgmt_gpio_out[9]
port 65 nsew signal input
rlabel metal2 s 8206 9200 8262 10000 6 mgmt_gpio_out_buf[0]
port 66 nsew signal output
rlabel metal2 s 2686 9200 2742 10000 6 mgmt_gpio_out_buf[10]
port 67 nsew signal output
rlabel metal2 s 2134 9200 2190 10000 6 mgmt_gpio_out_buf[11]
port 68 nsew signal output
rlabel metal2 s 1582 9200 1638 10000 6 mgmt_gpio_out_buf[12]
port 69 nsew signal output
rlabel metal2 s 1030 9200 1086 10000 6 mgmt_gpio_out_buf[13]
port 70 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 mgmt_gpio_out_buf[14]
port 71 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 mgmt_gpio_out_buf[15]
port 72 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 mgmt_gpio_out_buf[16]
port 73 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 mgmt_gpio_out_buf[17]
port 74 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 mgmt_gpio_out_buf[18]
port 75 nsew signal output
rlabel metal2 s 7654 9200 7710 10000 6 mgmt_gpio_out_buf[1]
port 76 nsew signal output
rlabel metal2 s 7102 9200 7158 10000 6 mgmt_gpio_out_buf[2]
port 77 nsew signal output
rlabel metal2 s 6550 9200 6606 10000 6 mgmt_gpio_out_buf[3]
port 78 nsew signal output
rlabel metal2 s 5998 9200 6054 10000 6 mgmt_gpio_out_buf[4]
port 79 nsew signal output
rlabel metal2 s 5446 9200 5502 10000 6 mgmt_gpio_out_buf[5]
port 80 nsew signal output
rlabel metal2 s 4894 9200 4950 10000 6 mgmt_gpio_out_buf[6]
port 81 nsew signal output
rlabel metal2 s 4342 9200 4398 10000 6 mgmt_gpio_out_buf[7]
port 82 nsew signal output
rlabel metal2 s 3790 9200 3846 10000 6 mgmt_gpio_out_buf[8]
port 83 nsew signal output
rlabel metal2 s 3238 9200 3294 10000 6 mgmt_gpio_out_buf[9]
port 84 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 9000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 243482
string GDS_FILE /home/hosni/caravel_sky130/caravel_redesign-2/caravel/openlane/mprj_io_buffer/runs/23_02_27_07_42/results/signoff/mprj_io_buffer.magic.gds
string GDS_START 27902
<< end >>

