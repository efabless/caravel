VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_id_programming
  CLASS BLOCK ;
  FOREIGN user_id_programming ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.545 BY 35.385 ;
  PIN mask_rev[0]
    PORT
      LAYER met2 ;
        RECT 20.330 31.385 20.610 35.385 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    PORT
      LAYER met2 ;
        RECT 26.770 31.385 27.050 35.385 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END mask_rev[14]
  PIN mask_rev[16]
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    PORT
      LAYER met2 ;
        RECT 8.370 31.385 8.650 35.385 ;
    END
  END mask_rev[17]
  PIN mask_rev[19]
    PORT
      LAYER met2 ;
        RECT 14.810 31.385 15.090 35.385 ;
    END
  END mask_rev[19]
  PIN mask_rev[23]
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    PORT
      LAYER met2 ;
        RECT 29.530 31.385 29.810 35.385 ;
    END
  END mask_rev[24]
  PIN mask_rev[26]
    PORT
      LAYER met2 ;
        RECT 24.010 31.385 24.290 35.385 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    PORT
      LAYER met2 ;
        RECT 5.610 31.385 5.890 35.385 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    PORT
      LAYER met2 ;
        RECT 32.290 31.385 32.570 35.385 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END mask_rev[29]
  PIN mask_rev[31]
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END mask_rev[3]
  PIN mask_rev[7]
    PORT
      LAYER met2 ;
        RECT 17.570 31.385 17.850 35.385 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    PORT
      LAYER met2 ;
        RECT 11.130 31.385 11.410 35.385 ;
    END
  END mask_rev[9]
  PIN mask_rev[15]
    PORT
      LAYER met3 ;
        RECT 31.545 8.200 35.545 8.800 ;
    END
  END mask_rev[15]
  PIN mask_rev[18]
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END mask_rev[18]
  PIN mask_rev[1]
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    PORT
      LAYER met3 ;
        RECT 31.545 12.280 35.545 12.880 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    PORT
      LAYER met3 ;
        RECT 31.545 4.120 35.545 4.720 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END mask_rev[22]
  PIN mask_rev[25]
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END mask_rev[25]
  PIN mask_rev[2]
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    PORT
      LAYER met3 ;
        RECT 31.545 25.880 35.545 26.480 ;
    END
  END mask_rev[30]
  PIN mask_rev[4]
    PORT
      LAYER met3 ;
        RECT 31.545 17.720 35.545 18.320 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    PORT
      LAYER met3 ;
        RECT 31.545 21.800 35.545 22.400 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END mask_rev[6]
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 20.720 29.900 22.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 12.560 29.900 14.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.970 5.200 22.570 30.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.845 5.200 14.445 30.160 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 16.640 29.900 18.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 24.800 29.900 26.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 8.480 29.900 10.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.780 5.200 10.380 30.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.910 5.200 18.510 30.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.035 5.200 26.635 30.160 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 29.900 30.005 ;
      LAYER met1 ;
        RECT 2.830 5.200 32.590 30.160 ;
      LAYER met2 ;
        RECT 2.860 31.105 5.330 31.385 ;
        RECT 6.170 31.105 8.090 31.385 ;
        RECT 8.930 31.105 10.850 31.385 ;
        RECT 11.690 31.105 14.530 31.385 ;
        RECT 15.370 31.105 17.290 31.385 ;
        RECT 18.130 31.105 20.050 31.385 ;
        RECT 20.890 31.105 23.730 31.385 ;
        RECT 24.570 31.105 26.490 31.385 ;
        RECT 27.330 31.105 29.250 31.385 ;
        RECT 30.090 31.105 32.010 31.385 ;
        RECT 2.860 4.280 32.560 31.105 ;
        RECT 3.410 4.000 5.330 4.280 ;
        RECT 6.170 4.000 8.090 4.280 ;
        RECT 8.930 4.000 10.850 4.280 ;
        RECT 11.690 4.000 14.530 4.280 ;
        RECT 15.370 4.000 17.290 4.280 ;
        RECT 18.130 4.000 20.050 4.280 ;
        RECT 20.890 4.000 23.730 4.280 ;
        RECT 24.570 4.000 26.490 4.280 ;
        RECT 27.330 4.000 29.250 4.280 ;
        RECT 30.090 4.000 32.560 4.280 ;
      LAYER met3 ;
        RECT 4.400 29.560 31.545 30.410 ;
        RECT 4.000 26.880 31.545 29.560 ;
        RECT 4.400 25.480 31.145 26.880 ;
        RECT 4.000 22.800 31.545 25.480 ;
        RECT 4.400 21.400 31.145 22.800 ;
        RECT 4.000 18.720 31.545 21.400 ;
        RECT 4.000 17.360 31.145 18.720 ;
        RECT 4.400 17.320 31.145 17.360 ;
        RECT 4.400 15.960 31.545 17.320 ;
        RECT 4.000 13.280 31.545 15.960 ;
        RECT 4.400 11.880 31.145 13.280 ;
        RECT 4.000 9.200 31.545 11.880 ;
        RECT 4.400 7.800 31.145 9.200 ;
        RECT 4.000 5.120 31.545 7.800 ;
        RECT 4.000 4.255 31.145 5.120 ;
  END
END user_id_programming
END LIBRARY
