VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO empty_macro
  CLASS BLOCK ;
  FOREIGN empty_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 25.000 ;
END empty_macro
END LIBRARY

