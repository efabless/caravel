magic
tech sky130A
magscale 1 2
timestamp 1638470713
<< pwell >>
rect 397 -17 431 17
rect 673 -17 707 17
rect 1411 -10 1443 12
rect 1685 -17 1719 17
rect 2881 -17 2915 17
rect 4077 -17 4111 17
rect 4812 -11 4836 11
rect 5090 -17 5124 17
rect 5272 -11 5296 11
rect 5457 -17 5491 17
rect 5551 -10 5583 12
rect 6008 -17 6042 17
rect 6101 -17 6135 17
rect 6470 -17 6504 17
rect 6837 -17 6871 17
rect 7667 -10 7699 12
rect 7849 -17 7883 17
rect 8493 -17 8527 17
rect 8861 -17 8895 17
rect 9505 -17 9539 17
rect 9872 -11 9896 11
rect 10057 -17 10091 17
rect 11253 -17 11287 17
rect 12449 -17 12483 17
rect 13092 -11 13116 11
rect 13368 -17 13402 17
rect 13460 -11 13484 11
rect 13645 -17 13679 17
rect 14840 -11 14864 11
rect 15025 -17 15059 17
rect 15117 -17 15151 17
rect 15852 -11 15876 11
rect 16037 -17 16071 17
rect 17233 -17 17267 17
rect 17879 -10 17911 12
rect 18245 -17 18279 17
rect 18429 -17 18463 17
rect 18797 -17 18831 17
<< obsli1 >>
rect 213 0 18860 10897
rect 368 -17 18860 0
<< obsm1 >>
rect 201 0 18860 10928
rect 368 -48 18860 0
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
<< obsm2 >>
rect 664 11144 1342 11257
rect 1510 11144 4194 11257
rect 4362 11144 7046 11257
rect 7214 11144 9898 11257
rect 10066 11144 12750 11257
rect 12918 11144 15602 11257
rect 15770 11144 18454 11257
rect 18622 11144 18842 11257
rect 664 0 18842 11144
rect 5028 -48 5336 0
rect 8128 -48 8436 0
rect 11228 -48 11536 0
rect 14328 -48 14636 0
rect 17428 -48 17736 0
<< metal3 >>
rect 19200 11160 20000 11280
rect 19200 9664 20000 9784
rect 19200 8168 20000 8288
rect 19200 6672 20000 6792
rect 19200 5176 20000 5296
rect 19200 3680 20000 3800
rect 19200 2184 20000 2304
rect 19200 688 20000 808
<< obsm3 >>
rect 2497 11080 19120 11253
rect 2497 9864 19200 11080
rect 2497 9584 19120 9864
rect 2497 8368 19200 9584
rect 2497 8088 19120 8368
rect 2497 6872 19200 8088
rect 2497 6592 19120 6872
rect 2497 5376 19200 6592
rect 2497 5096 19120 5376
rect 2497 3880 19200 5096
rect 2497 3600 19120 3880
rect 2497 2384 19200 3600
rect 2497 2104 19120 2384
rect 2497 888 19200 2104
rect 2497 608 19120 888
rect 2497 0 19200 608
rect 5022 -33 5342 0
rect 8122 -33 8442 0
rect 11222 -33 11542 0
rect 14322 -33 14642 0
rect 17422 -33 17742 0
<< metal4 >>
rect 3472 -48 3792 10928
rect 5022 -48 5342 10928
rect 6572 -48 6892 10928
rect 8122 -48 8442 10928
rect 9672 -48 9992 10928
rect 11222 -48 11542 10928
rect 12772 -48 13092 10928
rect 14322 -48 14642 10928
rect 15872 -48 16192 10928
rect 17422 -48 17742 10928
<< metal5 >>
rect 368 9882 18860 10202
rect 368 8192 18860 8512
rect 368 6502 18860 6822
rect 368 4812 18860 5132
rect 368 3122 18860 3442
<< labels >>
rlabel metal5 s 368 4812 18860 5132 6 VGND
port 1 nsew ground input
rlabel metal5 s 368 8192 18860 8512 6 VGND
port 1 nsew ground input
rlabel metal4 s 5022 -48 5342 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 8122 -48 8442 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 11222 -48 11542 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 14322 -48 14642 10928 6 VGND
port 1 nsew ground input
rlabel metal4 s 17422 -48 17742 10928 6 VGND
port 1 nsew ground input
rlabel metal5 s 368 3122 18860 3442 6 VPWR
port 2 nsew power input
rlabel metal5 s 368 6502 18860 6822 6 VPWR
port 2 nsew power input
rlabel metal5 s 368 9882 18860 10202 6 VPWR
port 2 nsew power input
rlabel metal4 s 3472 -48 3792 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 6572 -48 6892 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 9672 -48 9992 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 12772 -48 13092 10928 6 VPWR
port 2 nsew power input
rlabel metal4 s 15872 -48 16192 10928 6 VPWR
port 2 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 3 nsew signal output
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 4 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 5 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 6 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 7 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 8 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 9 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 10 nsew signal output
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 11 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 12 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 13 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 14 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 15 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 16 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 17 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 20000 12000
string LEFview TRUE
string GDS_FILE ../gds/caravel_clocking.gds
string GDS_END 1177254
string GDS_START 407686
<< end >>

