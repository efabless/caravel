* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbn_2 abstract view
.subckt sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_16 abstract view
.subckt sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_0 abstract view
.subckt sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_0 abstract view
.subckt sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__macro_sparecell abstract view
.subckt sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
.ends

* Black-box entry subcircuit for gpio_logic_high abstract view
.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
XFILLER_3_89 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_062_ _106_/Q user_gpio_out vssd vssd vccd vccd _062_/Y sky130_fd_sc_hd__nand2b_2
X_131_ _131_/CLK hold4/X _086_/A vssd vssd vccd vccd hold3/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_114_ _101__9/Y hold4/X _084_/X _085_/Y vssd vssd vccd vccd _114_/Q _114_/Q_N sky130_fd_sc_hd__dfbbn_2
Xoutput20 _134_/X vssd vssd vccd vccd resetn_out sky130_fd_sc_hd__buf_16
X_104__12 _100__8/A vssd vssd vccd vccd _104__12/Y sky130_fd_sc_hd__inv_2
Xoutput7 _116_/Q vssd vssd vccd vccd pad_gpio_ana_en sky130_fd_sc_hd__buf_16
X_130_ _130_/CLK hold9/X _086_/A vssd vssd vccd vccd hold4/A sky130_fd_sc_hd__dfrtp_4
X_094__2 _101__9/A vssd vssd vccd vccd _094__2/Y sky130_fd_sc_hd__inv_2
X_061_ user_gpio_oeb _060_/X _106_/Q vssd vssd vccd vccd _061_/X sky130_fd_sc_hd__mux2_4
X_113_ _100__8/Y hold9/X _082_/X _083_/Y vssd vssd vccd vccd _113_/Q _113_/Q_N sky130_fd_sc_hd__dfbbn_2
Xclkbuf_1_0__f_serial_load clkbuf_0_serial_load/X vssd vssd vccd vccd _100__8/A sky130_fd_sc_hd__clkbuf_16
X_059__14 _130_/CLK vssd vssd vccd vccd _132_/CLK sky130_fd_sc_hd__inv_2
Xoutput21 _132_/Q vssd vssd vccd vccd serial_data_out sky130_fd_sc_hd__buf_16
Xoutput8 _118_/Q vssd vssd vccd vccd pad_gpio_ana_pol sky130_fd_sc_hd__buf_16
Xoutput10 _113_/Q vssd vssd vccd vccd pad_gpio_dm[0] sky130_fd_sc_hd__buf_16
X_060_ _112_/Q _063_/C vssd vssd vccd vccd _060_/X sky130_fd_sc_hd__and2_0
X_112_ _099__7/Y hold6/X _080_/X _081_/Y vssd vssd vccd vccd _112_/Q _112_/Q_N sky130_fd_sc_hd__dfbbn_2
Xhold10 _127_/Q vssd vssd vccd vccd _128_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput22 _067_/X vssd vssd vccd vccd user_gpio_in sky130_fd_sc_hd__buf_16
Xoutput9 _117_/Q vssd vssd vccd vccd pad_gpio_ana_sel sky130_fd_sc_hd__buf_16
Xoutput11 _114_/Q vssd vssd vccd vccd pad_gpio_dm[1] sky130_fd_sc_hd__buf_16
X_111_ _098__6/Y hold8/X _078_/X _079_/Y vssd vssd vccd vccd _111_/Q _111_/Q_N sky130_fd_sc_hd__dfbbn_2
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold11 _126_/Q vssd vssd vccd vccd _127_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput12 _115_/Q vssd vssd vccd vccd pad_gpio_dm[2] sky130_fd_sc_hd__buf_16
X_110_ _097__5/Y hold7/X _076_/X _077_/Y vssd vssd vccd vccd _110_/Q _110_/Q_N sky130_fd_sc_hd__dfbbn_2
Xhold12 _125_/Q vssd vssd vccd vccd _126_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout29_A _082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__072__B gpio_defaults[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_097__5 _101__9/A vssd vssd vccd vccd _097__5/Y sky130_fd_sc_hd__inv_2
Xoutput13 _107_/Q vssd vssd vccd vccd pad_gpio_holdover sky130_fd_sc_hd__buf_16
XANTENNA__080__B gpio_defaults[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__075__B gpio_defaults[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold13 _124_/Q vssd vssd vccd vccd _125_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__083__B gpio_defaults[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput14 _111_/Q vssd vssd vccd vccd pad_gpio_ib_mode_sel sky130_fd_sc_hd__buf_16
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__078__B gpio_defaults[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__091__B gpio_defaults[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__086__B gpio_defaults[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput15 _110_/Q vssd vssd vccd vccd pad_gpio_inenb sky130_fd_sc_hd__buf_16
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__089__B gpio_defaults[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xconst_source vssd vssd vccd vccd one_buffer/A zero_buffer/A sky130_fd_sc_hd__conb_1
XANTENNA_fanout27_A _082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput16 _066_/Y vssd vssd vccd vccd pad_gpio_out sky130_fd_sc_hd__buf_16
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput17 _061_/X vssd vssd vccd vccd pad_gpio_outenb sky130_fd_sc_hd__buf_16
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xfanout30 fanout31/X vssd vssd vccd vccd _082_/A sky130_fd_sc_hd__buf_2
X_079_ _088_/A gpio_defaults[4] vssd vssd vccd vccd _079_/Y sky130_fd_sc_hd__nand2b_2
Xoutput18 _108_/Q vssd vssd vccd vccd pad_gpio_slow_sel sky130_fd_sc_hd__buf_16
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_100__8 _100__8/A vssd vssd vccd vccd _100__8/Y sky130_fd_sc_hd__inv_2
XANTENNA_input4_A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xfanout31 input4/X vssd vssd vccd vccd fanout31/X sky130_fd_sc_hd__buf_2
Xoutput19 _109_/Q vssd vssd vccd vccd pad_gpio_vtrip_sel sky130_fd_sc_hd__buf_16
X_078_ _088_/A gpio_defaults[4] vssd vssd vccd vccd _078_/X sky130_fd_sc_hd__or2_0
X_103__11 _100__8/A vssd vssd vccd vccd _103__11/Y sky130_fd_sc_hd__inv_2
XANTENNA__061__A0 user_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_34 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_129_ _131_/CLK hold2/X _074_/A vssd vssd vccd vccd hold9/A sky130_fd_sc_hd__dfrtp_4
X_077_ _076_/A gpio_defaults[3] vssd vssd vccd vccd _077_/Y sky130_fd_sc_hd__nand2b_2
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_093_ _092_/A gpio_defaults[7] vssd vssd vccd vccd _093_/Y sky130_fd_sc_hd__nand2b_2
X_076_ _076_/A gpio_defaults[3] vssd vssd vccd vccd _076_/X sky130_fd_sc_hd__or2_0
Xinput1 mgmt_gpio_oeb vssd vssd vccd vccd _063_/C sky130_fd_sc_hd__buf_2
X_128_ _131_/CLK _128_/D _074_/A vssd vssd vccd vccd hold2/A sky130_fd_sc_hd__dfrtp_4
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xfanout23 _092_/A vssd vssd vccd vccd _088_/A sky130_fd_sc_hd__buf_2
X_092_ _092_/A gpio_defaults[7] vssd vssd vccd vccd _092_/X sky130_fd_sc_hd__or2_0
XANTENNA_input2_A mgmt_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput2 mgmt_gpio_out vssd vssd vccd vccd input2/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_0_serial_load_A serial_load vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_075_ _074_/A gpio_defaults[9] vssd vssd vccd vccd _075_/Y sky130_fd_sc_hd__nand2b_2
X_127_ _130_/CLK _127_/D _092_/A vssd vssd vccd vccd _127_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xfanout24 fanout31/X vssd vssd vccd vccd _092_/A sky130_fd_sc_hd__buf_2
X_095__3 _100__8/A vssd vssd vccd vccd _095__3/Y sky130_fd_sc_hd__inv_2
XTAP_70 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_074_ _074_/A gpio_defaults[9] vssd vssd vccd vccd _074_/X sky130_fd_sc_hd__or2_0
X_091_ _088_/A gpio_defaults[6] vssd vssd vccd vccd _091_/Y sky130_fd_sc_hd__nand2b_2
Xinput3 pad_gpio_in vssd vssd vccd vccd _133_/A sky130_fd_sc_hd__buf_2
X_126_ _130_/CLK _126_/D _088_/A vssd vssd vccd vccd _126_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_109_ _096__4/Y hold2/X _074_/X _075_/Y vssd vssd vccd vccd _109_/Q _109_/Q_N sky130_fd_sc_hd__dfbbn_2
Xfanout25 _080_/A vssd vssd vccd vccd _076_/A sky130_fd_sc_hd__buf_2
XTAP_71 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 resetn vssd vssd vccd vccd input4/X sky130_fd_sc_hd__buf_2
X_090_ _092_/A gpio_defaults[6] vssd vssd vccd vccd _090_/X sky130_fd_sc_hd__or2_0
XFILLER_5_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_073_ _074_/A gpio_defaults[8] vssd vssd vccd vccd _073_/Y sky130_fd_sc_hd__nand2b_2
X_125_ _130_/CLK _125_/D _088_/A vssd vssd vccd vccd _125_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__062__B user_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__070__B gpio_defaults[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_108_ _095__3/Y _128_/D _072_/X _073_/Y vssd vssd vccd vccd _108_/Q _108_/Q_N sky130_fd_sc_hd__dfbbn_2
Xfanout26 fanout31/X vssd vssd vccd vccd _080_/A sky130_fd_sc_hd__buf_2
XTAP_72 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_072_ _074_/A gpio_defaults[8] vssd vssd vccd vccd _072_/X sky130_fd_sc_hd__or2_0
XTAP_61 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 serial_data_in vssd vssd vccd vccd _119_/D sky130_fd_sc_hd__buf_2
XTAP_50 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__073__B gpio_defaults[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_124_ _130_/CLK hold8/X _092_/A vssd vssd vccd vccd _124_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__068__B gpio_defaults[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_107_ _094__2/Y hold5/X _070_/X _071_/Y vssd vssd vccd vccd _107_/Q _107_/Q_N sky130_fd_sc_hd__dfbbn_2
Xfanout27 _082_/A vssd vssd vccd vccd _074_/A sky130_fd_sc_hd__buf_2
XANTENNA__076__B gpio_defaults[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__081__B gpio_defaults[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_73 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_071_ _076_/A gpio_defaults[2] vssd vssd vccd vccd _071_/Y sky130_fd_sc_hd__nand2b_2
XTAP_62 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ _058__1/Y hold1/X _068_/X _069_/Y vssd vssd vccd vccd _106_/Q _106_/Q_N sky130_fd_sc_hd__dfbbn_2
X_123_ _131_/CLK hold7/X _092_/A vssd vssd vccd vccd hold8/A sky130_fd_sc_hd__dfrtp_4
X_098__6 _100__8/A vssd vssd vccd vccd _098__6/Y sky130_fd_sc_hd__inv_2
XANTENNA__084__B gpio_defaults[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__079__B gpio_defaults[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xfanout28 _082_/A vssd vssd vccd vccd _086_/A sky130_fd_sc_hd__buf_2
XTAP_63 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ _076_/A gpio_defaults[2] vssd vssd vccd vccd _070_/X sky130_fd_sc_hd__or2_0
XANTENNA__092__B gpio_defaults[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_52 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__087__B gpio_defaults[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_122_ _130_/CLK hold5/X _076_/A vssd vssd vccd vccd hold7/A sky130_fd_sc_hd__dfrtp_4
Xspare_cell vssd vssd vccd vccd spare_cell/LO sky130_fd_sc_hd__macro_sparecell
Xserial_clock_out_buffer _131_/CLK vssd vssd vccd vccd serial_clock_out sky130_fd_sc_hd__clkbuf_16
Xfanout29 _082_/A vssd vssd vccd vccd _134_/A sky130_fd_sc_hd__buf_2
XTAP_64 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_121_ _130_/CLK hold6/X _076_/A vssd vssd vccd vccd hold5/A sky130_fd_sc_hd__dfrtp_4
XTAP_65 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_120_ _130_/CLK hold1/X _076_/A vssd vssd vccd vccd hold6/A sky130_fd_sc_hd__dfrtp_4
X_102__10 _101__9/A vssd vssd vccd vccd _102__10/Y sky130_fd_sc_hd__inv_2
X_058__1 _101__9/A vssd vssd vccd vccd _058__1/Y sky130_fd_sc_hd__inv_2
Xhold1 hold1/A vssd vssd vccd vccd hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_66 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd vssd vccd vccd hold2/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_serial_load serial_load vssd vssd vccd vccd clkbuf_0_serial_load/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _130_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_67 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xgpio_logic_high _067_/A vccd1 vssd1 gpio_logic_high
XTAP_45 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xone_buffer one_buffer/A vssd vssd vccd vccd one sky130_fd_sc_hd__buf_16
Xhold3 hold3/A vssd vssd vccd vccd hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_68 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_57 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_101__9 _101__9/A vssd vssd vccd vccd _101__9/Y sky130_fd_sc_hd__inv_2
XTAP_46 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout28_A _082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd vssd vccd vccd hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_69 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xhold5 hold5/A vssd vssd vccd vccd hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_59 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_48 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd vssd vccd vccd hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_089_ _088_/A gpio_defaults[5] vssd vssd vccd vccd _089_/Y sky130_fd_sc_hd__nand2b_2
Xzero_buffer zero_buffer/A vssd vssd vccd vccd zero sky130_fd_sc_hd__buf_16
XTAP_49 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0_serial_clock serial_clock vssd vssd vccd vccd clkbuf_0_serial_clock/X sky130_fd_sc_hd__clkbuf_16
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_105__13 _100__8/A vssd vssd vccd vccd _105__13/Y sky130_fd_sc_hd__inv_2
XANTENNA_input5_A serial_data_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_088_ _088_/A gpio_defaults[5] vssd vssd vccd vccd _088_/X sky130_fd_sc_hd__or2_0
XFILLER_3_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold7 hold7/A vssd vssd vccd vccd hold7/X sky130_fd_sc_hd__dlygate4sd3_1
X_096__4 _101__9/A vssd vssd vccd vccd _096__4/Y sky130_fd_sc_hd__inv_2
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold8 hold8/A vssd vssd vccd vccd hold8/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f_serial_load clkbuf_0_serial_load/X vssd vssd vccd vccd _101__9/A sky130_fd_sc_hd__clkbuf_16
X_087_ _134_/A gpio_defaults[12] vssd vssd vccd vccd _087_/Y sky130_fd_sc_hd__nand2b_2
XANTENNA__071__B gpio_defaults[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__082__A _082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _131_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__074__B gpio_defaults[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_086_ _086_/A gpio_defaults[12] vssd vssd vccd vccd _086_/X sky130_fd_sc_hd__or2_0
Xhold9 hold9/A vssd vssd vccd vccd hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__069__B gpio_defaults[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_069_ _086_/A gpio_defaults[0] vssd vssd vccd vccd _069_/Y sky130_fd_sc_hd__nand2b_2
XANTENNA__082__B gpio_defaults[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__077__B gpio_defaults[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input3_A pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_085_ _086_/A gpio_defaults[11] vssd vssd vccd vccd _085_/Y sky130_fd_sc_hd__nand2b_2
XANTENNA__090__B gpio_defaults[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__085__B gpio_defaults[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_068_ _086_/A gpio_defaults[0] vssd vssd vccd vccd _068_/X sky130_fd_sc_hd__or2_0
XFILLER_0_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__093__B gpio_defaults[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__088__B gpio_defaults[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_099__7 _101__9/A vssd vssd vccd vccd _099__7/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_084_ _086_/A gpio_defaults[11] vssd vssd vccd vccd _084_/X sky130_fd_sc_hd__or2_0
X_067_ _067_/A _133_/A vssd vssd vccd vccd _067_/X sky130_fd_sc_hd__and2_2
X_119_ _131_/CLK _119_/D _080_/A vssd vssd vccd vccd hold1/A sky130_fd_sc_hd__dfrtp_4
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_71 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_083_ _074_/A gpio_defaults[10] vssd vssd vccd vccd _083_/Y sky130_fd_sc_hd__nand2b_2
X_066_ _064_/X _065_/Y _062_/Y vssd vssd vccd vccd _066_/Y sky130_fd_sc_hd__o21ai_4
X_118_ _105__13/Y _127_/D _092_/X _093_/Y vssd vssd vccd vccd _118_/Q _118_/Q_N sky130_fd_sc_hd__dfbbn_2
XFILLER_0_31 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_065_ input2/X _064_/B _106_/Q vssd vssd vccd vccd _065_/Y sky130_fd_sc_hd__o21ai_2
X_082_ _082_/A gpio_defaults[10] vssd vssd vccd vccd _082_/X sky130_fd_sc_hd__or2_0
X_134_ _134_/A vssd vssd vccd vccd _134_/X sky130_fd_sc_hd__buf_2
Xserial_load_out_buffer _101__9/A vssd vssd vccd vccd serial_load_out sky130_fd_sc_hd__clkbuf_16
XANTENNA_input1_A mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_117_ _104__12/Y _126_/D _090_/X _091_/Y vssd vssd vccd vccd _117_/Q _117_/Q_N sky130_fd_sc_hd__dfbbn_2
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_081_ _080_/A gpio_defaults[1] vssd vssd vccd vccd _081_/Y sky130_fd_sc_hd__nand2b_2
X_064_ _113_/Q_N _064_/B vssd vssd vccd vccd _064_/X sky130_fd_sc_hd__and2b_2
X_133_ _133_/A vssd vssd vccd vccd _133_/X sky130_fd_sc_hd__buf_2
X_116_ _103__11/Y _125_/D _088_/X _089_/Y vssd vssd vccd vccd _116_/Q _116_/Q_N sky130_fd_sc_hd__dfbbn_2
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_serial_clock_A serial_clock vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_132_ _132_/CLK hold3/A _134_/A vssd vssd vccd vccd _132_/Q sky130_fd_sc_hd__dfrtp_2
X_080_ _080_/A gpio_defaults[1] vssd vssd vccd vccd _080_/X sky130_fd_sc_hd__or2_0
X_063_ _115_/Q _114_/Q _063_/C vssd vssd vccd vccd _064_/B sky130_fd_sc_hd__and3b_2
X_115_ _102__10/Y hold3/X _086_/X _087_/Y vssd vssd vccd vccd _115_/Q _115_/Q_N sky130_fd_sc_hd__dfbbn_2
Xoutput6 _133_/X vssd vssd vccd vccd mgmt_gpio_in sky130_fd_sc_hd__buf_16
.ends

