VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_control_block
  CLASS BLOCK ;
  FOREIGN gpio_control_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 65.000 ;
  PIN gpio_defaults[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 61.000 4.970 65.000 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 61.000 27.970 65.000 ;
    END
  END gpio_defaults[10]
  PIN gpio_defaults[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 61.000 30.270 65.000 ;
    END
  END gpio_defaults[11]
  PIN gpio_defaults[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 61.000 32.570 65.000 ;
    END
  END gpio_defaults[12]
  PIN gpio_defaults[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 61.000 7.270 65.000 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 61.000 9.570 65.000 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 61.000 11.870 65.000 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 61.000 14.170 65.000 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 61.000 16.470 65.000 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 61.000 18.770 65.000 ;
    END
  END gpio_defaults[6]
  PIN gpio_defaults[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 61.000 21.070 65.000 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 61.000 23.370 65.000 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 61.000 25.670 65.000 ;
    END
  END gpio_defaults[9]
  PIN mgmt_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 4.120 170.000 4.720 ;
    END
  END mgmt_gpio_in
  PIN mgmt_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 8.200 170.000 8.800 ;
    END
  END mgmt_gpio_oeb
  PIN mgmt_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 10.240 170.000 10.840 ;
    END
  END mgmt_gpio_out
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 6.160 170.000 6.760 ;
    END
  END one
  PIN pad_gpio_ana_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 12.280 170.000 12.880 ;
    END
  END pad_gpio_ana_en
  PIN pad_gpio_ana_pol
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 14.320 170.000 14.920 ;
    END
  END pad_gpio_ana_pol
  PIN pad_gpio_ana_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 16.360 170.000 16.960 ;
    END
  END pad_gpio_ana_sel
  PIN pad_gpio_dm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 18.400 170.000 19.000 ;
    END
  END pad_gpio_dm[0]
  PIN pad_gpio_dm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 20.440 170.000 21.040 ;
    END
  END pad_gpio_dm[1]
  PIN pad_gpio_dm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 22.480 170.000 23.080 ;
    END
  END pad_gpio_dm[2]
  PIN pad_gpio_holdover
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 24.520 170.000 25.120 ;
    END
  END pad_gpio_holdover
  PIN pad_gpio_ib_mode_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 26.560 170.000 27.160 ;
    END
  END pad_gpio_ib_mode_sel
  PIN pad_gpio_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 28.600 170.000 29.200 ;
    END
  END pad_gpio_in
  PIN pad_gpio_inenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 30.640 170.000 31.240 ;
    END
  END pad_gpio_inenb
  PIN pad_gpio_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 32.680 170.000 33.280 ;
    END
  END pad_gpio_out
  PIN pad_gpio_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 34.720 170.000 35.320 ;
    END
  END pad_gpio_outenb
  PIN pad_gpio_slow_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 36.760 170.000 37.360 ;
    END
  END pad_gpio_slow_sel
  PIN pad_gpio_vtrip_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 38.800 170.000 39.400 ;
    END
  END pad_gpio_vtrip_sel
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 40.840 170.000 41.440 ;
    END
  END resetn
  PIN resetn_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 42.880 170.000 43.480 ;
    END
  END resetn_out
  PIN serial_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 44.920 170.000 45.520 ;
    END
  END serial_clock
  PIN serial_clock_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 46.960 170.000 47.560 ;
    END
  END serial_clock_out
  PIN serial_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 49.000 170.000 49.600 ;
    END
  END serial_data_in
  PIN serial_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 51.040 170.000 51.640 ;
    END
  END serial_data_out
  PIN serial_load
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 53.080 170.000 53.680 ;
    END
  END serial_load
  PIN serial_load_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 55.120 170.000 55.720 ;
    END
  END serial_load_out
  PIN user_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 57.160 170.000 57.760 ;
    END
  END user_gpio_in
  PIN user_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 59.200 170.000 59.800 ;
    END
  END user_gpio_oeb
  PIN user_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 61.240 170.000 61.840 ;
    END
  END user_gpio_out
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 12.800 2.480 14.400 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.800 2.480 39.400 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 5.900 51.760 7.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 22.800 51.760 24.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 39.700 51.760 41.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 56.600 51.760 58.200 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.800 2.480 19.400 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.800 2.480 44.400 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 11.140 51.760 12.740 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 28.040 51.760 29.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 44.940 51.760 46.540 ;
    END
  END vccd1
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.300 2.480 26.900 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 14.350 51.760 15.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 31.250 51.760 32.850 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 48.150 51.760 49.750 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 30.300 2.480 31.900 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 19.590 51.760 21.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 36.490 51.760 38.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 53.390 51.760 54.990 ;
    END
  END vssd1
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 2.080 170.000 2.680 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 0.000 64.930 4.265 65.070 ;
      LAYER li1 ;
        RECT 4.265 64.930 169.810 65.000 ;
      LAYER li1 ;
        RECT 0.000 64.845 49.815 64.930 ;
      LAYER li1 ;
        RECT 49.815 64.845 169.810 64.930 ;
      LAYER li1 ;
        RECT 0.000 59.925 169.810 64.845 ;
        RECT 0.000 59.755 4.745 59.925 ;
      LAYER li1 ;
        RECT 4.745 59.755 169.810 59.925 ;
      LAYER li1 ;
        RECT 0.000 59.585 169.810 59.755 ;
        RECT 0.000 57.645 6.100 59.585 ;
      LAYER li1 ;
        RECT 6.100 57.645 169.810 59.585 ;
      LAYER li1 ;
        RECT 0.000 57.405 8.925 57.645 ;
      LAYER li1 ;
        RECT 8.925 57.405 169.810 57.645 ;
      LAYER li1 ;
        RECT 0.000 30.025 4.265 57.405 ;
      LAYER li1 ;
        RECT 4.265 30.025 169.810 57.405 ;
      LAYER li1 ;
        RECT 0.000 30.005 16.795 30.025 ;
      LAYER li1 ;
        RECT 16.795 30.005 169.810 30.025 ;
      LAYER li1 ;
        RECT 0.000 29.835 4.745 30.005 ;
      LAYER li1 ;
        RECT 4.745 29.835 169.810 30.005 ;
      LAYER li1 ;
        RECT 0.000 29.665 16.795 29.835 ;
      LAYER li1 ;
        RECT 16.795 29.665 169.810 29.835 ;
      LAYER li1 ;
        RECT 0.000 27.455 6.065 29.665 ;
      LAYER li1 ;
        RECT 6.065 27.455 169.810 29.665 ;
      LAYER li1 ;
        RECT 0.000 27.285 16.795 27.455 ;
      LAYER li1 ;
        RECT 16.795 27.285 169.810 27.455 ;
      LAYER li1 ;
        RECT 0.000 27.115 4.745 27.285 ;
      LAYER li1 ;
        RECT 4.745 27.115 169.810 27.285 ;
      LAYER li1 ;
        RECT 0.000 26.945 16.795 27.115 ;
      LAYER li1 ;
        RECT 16.795 26.945 169.810 27.115 ;
      LAYER li1 ;
        RECT 0.000 26.185 16.905 26.945 ;
      LAYER li1 ;
        RECT 16.905 26.185 169.810 26.945 ;
      LAYER li1 ;
        RECT 0.000 26.015 17.450 26.185 ;
      LAYER li1 ;
        RECT 17.450 26.015 169.810 26.185 ;
      LAYER li1 ;
        RECT 0.000 25.835 16.795 26.015 ;
      LAYER li1 ;
        RECT 16.795 25.835 169.810 26.015 ;
      LAYER li1 ;
        RECT 0.000 25.465 16.645 25.835 ;
      LAYER li1 ;
        RECT 16.645 25.465 169.810 25.835 ;
      LAYER li1 ;
        RECT 0.000 25.285 16.795 25.465 ;
      LAYER li1 ;
        RECT 16.795 25.285 169.810 25.465 ;
      LAYER li1 ;
        RECT 0.000 25.115 17.450 25.285 ;
      LAYER li1 ;
        RECT 17.450 25.115 169.810 25.285 ;
      LAYER li1 ;
        RECT 0.000 24.735 16.905 25.115 ;
      LAYER li1 ;
        RECT 16.905 24.735 169.810 25.115 ;
      LAYER li1 ;
        RECT 0.000 24.565 16.795 24.735 ;
      LAYER li1 ;
        RECT 16.795 24.565 169.810 24.735 ;
      LAYER li1 ;
        RECT 0.000 24.395 15.325 24.565 ;
      LAYER li1 ;
        RECT 15.325 24.395 169.810 24.565 ;
      LAYER li1 ;
        RECT 0.000 24.225 16.795 24.395 ;
      LAYER li1 ;
        RECT 16.795 24.225 169.810 24.395 ;
      LAYER li1 ;
        RECT 0.000 22.015 16.645 24.225 ;
      LAYER li1 ;
        RECT 16.645 22.015 169.810 24.225 ;
      LAYER li1 ;
        RECT 0.000 21.845 16.795 22.015 ;
      LAYER li1 ;
        RECT 16.795 21.845 169.810 22.015 ;
      LAYER li1 ;
        RECT 0.000 21.675 15.325 21.845 ;
      LAYER li1 ;
        RECT 15.325 21.675 169.810 21.845 ;
      LAYER li1 ;
        RECT 0.000 20.865 16.950 21.675 ;
      LAYER li1 ;
        RECT 16.950 20.865 169.810 21.675 ;
      LAYER li1 ;
        RECT 0.000 20.365 16.795 20.865 ;
      LAYER li1 ;
        RECT 16.795 20.365 169.810 20.865 ;
      LAYER li1 ;
        RECT 0.000 19.805 16.645 20.365 ;
      LAYER li1 ;
        RECT 16.645 19.805 169.810 20.365 ;
      LAYER li1 ;
        RECT 0.000 19.635 16.795 19.805 ;
      LAYER li1 ;
        RECT 16.795 19.635 169.810 19.805 ;
      LAYER li1 ;
        RECT 0.000 19.125 16.950 19.635 ;
      LAYER li1 ;
        RECT 16.950 19.125 169.810 19.635 ;
      LAYER li1 ;
        RECT 0.000 18.955 15.325 19.125 ;
      LAYER li1 ;
        RECT 15.325 18.955 169.810 19.125 ;
      LAYER li1 ;
        RECT 0.000 18.785 16.795 18.955 ;
      LAYER li1 ;
        RECT 16.795 18.785 169.810 18.955 ;
      LAYER li1 ;
        RECT 0.000 16.575 16.645 18.785 ;
      LAYER li1 ;
        RECT 16.645 16.575 169.810 18.785 ;
      LAYER li1 ;
        RECT 0.000 16.405 16.795 16.575 ;
      LAYER li1 ;
        RECT 16.795 16.405 169.810 16.575 ;
      LAYER li1 ;
        RECT 0.000 16.235 15.325 16.405 ;
      LAYER li1 ;
        RECT 15.325 16.235 169.810 16.405 ;
      LAYER li1 ;
        RECT 0.000 15.425 16.950 16.235 ;
      LAYER li1 ;
        RECT 16.950 15.425 169.810 16.235 ;
      LAYER li1 ;
        RECT 0.000 14.925 16.795 15.425 ;
      LAYER li1 ;
        RECT 16.795 14.925 169.810 15.425 ;
      LAYER li1 ;
        RECT 0.000 14.365 16.645 14.925 ;
      LAYER li1 ;
        RECT 16.645 14.365 169.810 14.925 ;
      LAYER li1 ;
        RECT 0.000 14.195 16.795 14.365 ;
      LAYER li1 ;
        RECT 16.795 14.195 169.810 14.365 ;
      LAYER li1 ;
        RECT 0.000 13.685 16.950 14.195 ;
      LAYER li1 ;
        RECT 16.950 13.685 169.810 14.195 ;
      LAYER li1 ;
        RECT 0.000 13.515 15.325 13.685 ;
      LAYER li1 ;
        RECT 15.325 13.515 169.810 13.685 ;
      LAYER li1 ;
        RECT 0.000 13.005 16.950 13.515 ;
      LAYER li1 ;
        RECT 16.950 13.005 169.810 13.515 ;
      LAYER li1 ;
        RECT 0.000 12.835 16.795 13.005 ;
      LAYER li1 ;
        RECT 16.795 12.835 169.810 13.005 ;
      LAYER li1 ;
        RECT 0.000 12.275 16.645 12.835 ;
      LAYER li1 ;
        RECT 16.645 12.275 169.810 12.835 ;
      LAYER li1 ;
        RECT 0.000 11.775 16.795 12.275 ;
      LAYER li1 ;
        RECT 16.795 11.775 169.810 12.275 ;
      LAYER li1 ;
        RECT 0.000 10.965 16.950 11.775 ;
      LAYER li1 ;
        RECT 16.950 10.965 169.810 11.775 ;
      LAYER li1 ;
        RECT 0.000 10.795 15.325 10.965 ;
      LAYER li1 ;
        RECT 15.325 10.795 169.810 10.965 ;
      LAYER li1 ;
        RECT 0.000 10.020 16.795 10.795 ;
      LAYER li1 ;
        RECT 16.795 10.020 169.810 10.795 ;
      LAYER li1 ;
        RECT 0.000 9.825 16.970 10.020 ;
      LAYER li1 ;
        RECT 16.970 9.825 169.810 10.020 ;
      LAYER li1 ;
        RECT 0.000 9.655 17.920 9.825 ;
      LAYER li1 ;
        RECT 17.920 9.655 169.810 9.825 ;
      LAYER li1 ;
        RECT 0.000 9.000 16.840 9.655 ;
      LAYER li1 ;
        RECT 16.840 9.000 169.810 9.655 ;
      LAYER li1 ;
        RECT 0.000 8.670 16.905 9.000 ;
      LAYER li1 ;
        RECT 16.905 8.670 169.810 9.000 ;
      LAYER li1 ;
        RECT 0.000 8.245 16.795 8.670 ;
      LAYER li1 ;
        RECT 16.795 8.245 169.810 8.670 ;
      LAYER li1 ;
        RECT 0.000 8.075 15.325 8.245 ;
      LAYER li1 ;
        RECT 15.325 8.075 169.810 8.245 ;
      LAYER li1 ;
        RECT 0.000 7.905 16.795 8.075 ;
      LAYER li1 ;
        RECT 16.795 7.905 169.810 8.075 ;
      LAYER li1 ;
        RECT 0.000 5.695 16.645 7.905 ;
      LAYER li1 ;
        RECT 16.645 5.695 169.810 7.905 ;
      LAYER li1 ;
        RECT 0.000 5.525 16.795 5.695 ;
      LAYER li1 ;
        RECT 16.795 5.525 169.810 5.695 ;
      LAYER li1 ;
        RECT 0.000 5.355 4.745 5.525 ;
      LAYER li1 ;
        RECT 4.745 5.355 169.810 5.525 ;
      LAYER li1 ;
        RECT 0.000 5.185 16.795 5.355 ;
      LAYER li1 ;
        RECT 16.795 5.185 169.810 5.355 ;
      LAYER li1 ;
        RECT 0.000 2.975 6.525 5.185 ;
      LAYER li1 ;
        RECT 6.525 2.975 169.810 5.185 ;
      LAYER li1 ;
        RECT 0.000 2.805 16.795 2.975 ;
      LAYER li1 ;
        RECT 16.795 2.805 169.810 2.975 ;
      LAYER li1 ;
        RECT 0.000 2.635 4.745 2.805 ;
      LAYER li1 ;
        RECT 4.745 2.635 169.810 2.805 ;
      LAYER li1 ;
        RECT 0.000 0.000 16.795 2.635 ;
      LAYER li1 ;
        RECT 16.795 0.000 169.810 2.635 ;
      LAYER met1 ;
        RECT 4.300 0.000 170.000 65.000 ;
      LAYER met2 ;
        RECT 5.250 60.720 6.710 65.000 ;
        RECT 7.550 60.720 9.010 65.000 ;
        RECT 9.850 60.720 11.310 65.000 ;
        RECT 12.150 60.720 13.610 65.000 ;
        RECT 14.450 60.720 15.910 65.000 ;
        RECT 16.750 60.720 18.210 65.000 ;
        RECT 19.050 60.720 20.510 65.000 ;
        RECT 21.350 60.720 22.810 65.000 ;
        RECT 23.650 60.720 25.110 65.000 ;
        RECT 25.950 60.720 27.410 65.000 ;
        RECT 28.250 60.720 29.710 65.000 ;
        RECT 30.550 60.720 32.010 65.000 ;
        RECT 32.850 60.720 170.000 65.000 ;
        RECT 4.700 0.000 170.000 60.720 ;
      LAYER met3 ;
        RECT 6.280 60.840 69.600 61.705 ;
        RECT 6.280 60.200 70.000 60.840 ;
        RECT 6.280 58.800 69.600 60.200 ;
        RECT 6.280 58.160 70.000 58.800 ;
        RECT 6.280 56.760 69.600 58.160 ;
        RECT 6.280 56.120 70.000 56.760 ;
        RECT 6.280 54.720 69.600 56.120 ;
        RECT 6.280 54.080 70.000 54.720 ;
        RECT 6.280 52.680 69.600 54.080 ;
        RECT 6.280 52.040 70.000 52.680 ;
        RECT 6.280 50.640 69.600 52.040 ;
        RECT 6.280 50.000 70.000 50.640 ;
        RECT 6.280 48.600 69.600 50.000 ;
        RECT 6.280 47.960 70.000 48.600 ;
        RECT 6.280 46.560 69.600 47.960 ;
        RECT 6.280 45.920 70.000 46.560 ;
        RECT 6.280 44.520 69.600 45.920 ;
        RECT 6.280 43.880 70.000 44.520 ;
        RECT 6.280 42.480 69.600 43.880 ;
        RECT 6.280 41.840 70.000 42.480 ;
        RECT 6.280 40.440 69.600 41.840 ;
        RECT 6.280 39.800 70.000 40.440 ;
        RECT 6.280 38.400 69.600 39.800 ;
        RECT 6.280 37.760 70.000 38.400 ;
        RECT 6.280 36.360 69.600 37.760 ;
        RECT 6.280 35.720 70.000 36.360 ;
        RECT 6.280 34.320 69.600 35.720 ;
        RECT 6.280 33.680 70.000 34.320 ;
        RECT 6.280 32.280 69.600 33.680 ;
        RECT 6.280 31.640 70.000 32.280 ;
        RECT 6.280 30.240 69.600 31.640 ;
        RECT 6.280 29.600 70.000 30.240 ;
        RECT 6.280 28.200 69.600 29.600 ;
        RECT 6.280 27.560 70.000 28.200 ;
        RECT 6.280 26.160 69.600 27.560 ;
        RECT 6.280 25.520 70.000 26.160 ;
        RECT 6.280 24.120 69.600 25.520 ;
        RECT 6.280 23.480 70.000 24.120 ;
        RECT 6.280 22.080 69.600 23.480 ;
        RECT 6.280 21.440 70.000 22.080 ;
        RECT 6.280 20.040 69.600 21.440 ;
        RECT 6.280 19.400 70.000 20.040 ;
        RECT 6.280 18.000 69.600 19.400 ;
        RECT 6.280 17.360 70.000 18.000 ;
        RECT 6.280 15.960 69.600 17.360 ;
        RECT 6.280 15.320 70.000 15.960 ;
        RECT 6.280 13.920 69.600 15.320 ;
        RECT 6.280 13.280 70.000 13.920 ;
        RECT 6.280 11.880 69.600 13.280 ;
        RECT 6.280 11.240 70.000 11.880 ;
        RECT 6.280 9.840 69.600 11.240 ;
        RECT 6.280 9.200 70.000 9.840 ;
        RECT 6.280 7.800 69.600 9.200 ;
        RECT 6.280 7.160 70.000 7.800 ;
        RECT 6.280 5.760 69.600 7.160 ;
        RECT 6.280 5.120 70.000 5.760 ;
        RECT 6.280 3.720 69.600 5.120 ;
        RECT 6.280 3.080 70.000 3.720 ;
        RECT 6.280 1.680 69.600 3.080 ;
        RECT 6.280 0.175 70.000 1.680 ;
      LAYER met4 ;
        RECT 6.280 60.480 170.000 65.000 ;
        RECT 6.280 2.080 12.400 60.480 ;
        RECT 14.800 2.080 17.400 60.480 ;
        RECT 19.800 2.080 24.900 60.480 ;
        RECT 27.300 2.080 29.900 60.480 ;
        RECT 32.300 2.080 37.400 60.480 ;
        RECT 39.800 2.080 42.400 60.480 ;
        RECT 44.800 2.080 170.000 60.480 ;
        RECT 6.280 0.000 170.000 2.080 ;
      LAYER met5 ;
        RECT 67.000 0.000 170.000 65.000 ;
  END
END gpio_control_block
END LIBRARY

