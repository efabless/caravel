magic
tech sky130A
timestamp 0
<< properties >>
string FIXED_BBOX 0 0 0 0
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29976804
string GDS_FILE /home/hosni/caravan/caravan-mpw9-PnR/caravel/openlane/housekeeping_alt/runs/23_05_23_06_27/results/signoff/housekeeping_alt.magic.gds
string GDS_START 1712610
<< end >>

