magic
tech sky130A
magscale 1 2
timestamp 1636370563
<< locali >>
rect 8309 13175 8343 13413
rect 1961 8959 1995 9061
rect 14013 7531 14047 12325
rect 14105 7871 14139 9877
rect 3065 6715 3099 6885
rect 14013 5899 14047 7361
rect 8769 5559 8803 5797
rect 14013 527 14047 2805
<< viali >>
rect 3525 13481 3559 13515
rect 3893 13481 3927 13515
rect 6193 13481 6227 13515
rect 8493 13481 8527 13515
rect 6929 13413 6963 13447
rect 8309 13413 8343 13447
rect 9689 13413 9723 13447
rect 3157 13277 3191 13311
rect 5273 13277 5307 13311
rect 6377 13277 6411 13311
rect 6750 13277 6784 13311
rect 7113 13277 7147 13311
rect 7389 13277 7423 13311
rect 7757 13277 7791 13311
rect 6561 13209 6595 13243
rect 6653 13209 6687 13243
rect 8677 13345 8711 13379
rect 9137 13345 9171 13379
rect 10241 13345 10275 13379
rect 9229 13277 9263 13311
rect 10701 13277 10735 13311
rect 12081 13277 12115 13311
rect 12725 13277 12759 13311
rect 10793 13209 10827 13243
rect 10885 13209 10919 13243
rect 12541 13209 12575 13243
rect 12633 13209 12667 13243
rect 13185 13209 13219 13243
rect 13277 13209 13311 13243
rect 3341 13141 3375 13175
rect 5365 13141 5399 13175
rect 7205 13141 7239 13175
rect 7665 13141 7699 13175
rect 8217 13141 8251 13175
rect 8309 13141 8343 13175
rect 9321 13141 9355 13175
rect 9873 13141 9907 13175
rect 10057 13141 10091 13175
rect 11069 13141 11103 13175
rect 4077 12937 4111 12971
rect 6009 12937 6043 12971
rect 8125 12937 8159 12971
rect 8309 12937 8343 12971
rect 9413 12937 9447 12971
rect 13369 12937 13403 12971
rect 6653 12869 6687 12903
rect 8953 12869 8987 12903
rect 11345 12869 11379 12903
rect 2329 12801 2363 12835
rect 8493 12801 8527 12835
rect 9045 12801 9079 12835
rect 9781 12801 9815 12835
rect 11253 12801 11287 12835
rect 11713 12801 11747 12835
rect 12909 12801 12943 12835
rect 13553 12801 13587 12835
rect 2605 12733 2639 12767
rect 4261 12733 4295 12767
rect 4537 12733 4571 12767
rect 6377 12733 6411 12767
rect 8861 12733 8895 12767
rect 9505 12665 9539 12699
rect 13001 12665 13035 12699
rect 4629 12393 4663 12427
rect 10149 12393 10183 12427
rect 11621 12393 11655 12427
rect 13369 12393 13403 12427
rect 3893 12325 3927 12359
rect 6561 12325 6595 12359
rect 14013 12325 14047 12359
rect 1685 12257 1719 12291
rect 4261 12257 4295 12291
rect 5365 12257 5399 12291
rect 5825 12257 5859 12291
rect 5917 12257 5951 12291
rect 6397 12257 6431 12291
rect 7297 12257 7331 12291
rect 7573 12257 7607 12291
rect 8033 12257 8067 12291
rect 1409 12189 1443 12223
rect 3433 12189 3467 12223
rect 3801 12189 3835 12223
rect 4077 12189 4111 12223
rect 4808 12189 4842 12223
rect 5181 12189 5215 12223
rect 5457 12189 5491 12223
rect 6009 12189 6043 12223
rect 6285 12189 6319 12223
rect 6837 12189 6871 12223
rect 7021 12189 7055 12223
rect 7113 12189 7147 12223
rect 7389 12189 7423 12223
rect 7665 12189 7699 12223
rect 8400 12189 8434 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 8769 12189 8803 12223
rect 8953 12189 8987 12223
rect 9229 12189 9263 12223
rect 9505 12189 9539 12223
rect 9597 12189 9631 12223
rect 10333 12189 10367 12223
rect 11069 12189 11103 12223
rect 11253 12189 11287 12223
rect 11529 12189 11563 12223
rect 11989 12189 12023 12223
rect 12265 12189 12299 12223
rect 13001 12189 13035 12223
rect 13277 12189 13311 12223
rect 4905 12121 4939 12155
rect 4997 12121 5031 12155
rect 8125 12121 8159 12155
rect 9321 12121 9355 12155
rect 12173 12121 12207 12155
rect 13185 12121 13219 12155
rect 3157 12053 3191 12087
rect 3617 12053 3651 12087
rect 9965 12053 9999 12087
rect 11345 12053 11379 12087
rect 2605 11849 2639 11883
rect 6745 11849 6779 11883
rect 10149 11849 10183 11883
rect 11621 11849 11655 11883
rect 5825 11781 5859 11815
rect 8493 11781 8527 11815
rect 8953 11781 8987 11815
rect 9321 11781 9355 11815
rect 11161 11781 11195 11815
rect 13093 11781 13127 11815
rect 2421 11713 2455 11747
rect 2789 11713 2823 11747
rect 5365 11713 5399 11747
rect 5457 11713 5491 11747
rect 6009 11713 6043 11747
rect 6101 11713 6135 11747
rect 6377 11713 6411 11747
rect 6653 11713 6687 11747
rect 7113 11713 7147 11747
rect 7849 11713 7883 11747
rect 8585 11713 8619 11747
rect 9137 11713 9171 11747
rect 9413 11713 9447 11747
rect 11069 11713 11103 11747
rect 11713 11713 11747 11747
rect 12265 11713 12299 11747
rect 1501 11645 1535 11679
rect 3157 11645 3191 11679
rect 3433 11645 3467 11679
rect 5733 11645 5767 11679
rect 6469 11645 6503 11679
rect 7941 11645 7975 11679
rect 8217 11645 8251 11679
rect 9873 11645 9907 11679
rect 10057 11645 10091 11679
rect 10609 11645 10643 11679
rect 12357 11645 12391 11679
rect 12909 11645 12943 11679
rect 12081 11577 12115 11611
rect 12817 11577 12851 11611
rect 2881 11509 2915 11543
rect 4905 11509 4939 11543
rect 5181 11509 5215 11543
rect 5641 11509 5675 11543
rect 7021 11509 7055 11543
rect 8677 11509 8711 11543
rect 9505 11509 9539 11543
rect 10517 11509 10551 11543
rect 11253 11509 11287 11543
rect 13185 11509 13219 11543
rect 3525 11305 3559 11339
rect 6469 11305 6503 11339
rect 7481 11305 7515 11339
rect 2789 11237 2823 11271
rect 3801 11237 3835 11271
rect 5457 11237 5491 11271
rect 5825 11237 5859 11271
rect 6285 11237 6319 11271
rect 7021 11237 7055 11271
rect 11529 11237 11563 11271
rect 13185 11237 13219 11271
rect 6653 11169 6687 11203
rect 7665 11169 7699 11203
rect 7941 11169 7975 11203
rect 9321 11169 9355 11203
rect 2973 11101 3007 11135
rect 3617 11101 3651 11135
rect 4076 11101 4110 11135
rect 4168 11095 4202 11129
rect 4261 11101 4295 11135
rect 4445 11095 4479 11129
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 5641 11101 5675 11135
rect 5733 11101 5767 11135
rect 5917 11101 5951 11135
rect 6101 11101 6135 11135
rect 6469 11101 6503 11135
rect 6745 11101 6779 11135
rect 6929 11101 6963 11135
rect 7205 11101 7239 11135
rect 7297 11101 7331 11135
rect 8033 11101 8067 11135
rect 8953 11101 8987 11135
rect 9118 11101 9152 11135
rect 9229 11101 9263 11135
rect 9505 11101 9539 11135
rect 9781 11101 9815 11135
rect 10241 11101 10275 11135
rect 11529 11101 11563 11135
rect 11897 11101 11931 11135
rect 13185 11101 13219 11135
rect 3341 11033 3375 11067
rect 4923 11033 4957 11067
rect 5089 11033 5123 11067
rect 9965 11033 9999 11067
rect 10149 11033 10183 11067
rect 3065 10965 3099 10999
rect 3157 10965 3191 10999
rect 4813 10965 4847 10999
rect 8677 10965 8711 10999
rect 9597 10965 9631 10999
rect 3157 10761 3191 10795
rect 8401 10761 8435 10795
rect 9597 10761 9631 10795
rect 9965 10761 9999 10795
rect 10057 10761 10091 10795
rect 10425 10761 10459 10795
rect 12357 10761 12391 10795
rect 5641 10693 5675 10727
rect 6469 10693 6503 10727
rect 7205 10693 7239 10727
rect 11253 10693 11287 10727
rect 12081 10693 12115 10727
rect 12449 10693 12483 10727
rect 13185 10693 13219 10727
rect 13461 10693 13495 10727
rect 1409 10625 1443 10659
rect 3709 10625 3743 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4996 10625 5030 10659
rect 5273 10625 5307 10659
rect 5457 10625 5491 10659
rect 5733 10625 5767 10659
rect 6377 10625 6411 10659
rect 6745 10625 6779 10659
rect 7481 10625 7515 10659
rect 8125 10625 8159 10659
rect 8585 10625 8619 10659
rect 8733 10628 8767 10662
rect 8953 10625 8987 10659
rect 9110 10625 9144 10659
rect 10793 10625 10827 10659
rect 11529 10625 11563 10659
rect 11805 10625 11839 10659
rect 12541 10625 12575 10659
rect 1685 10557 1719 10591
rect 3617 10557 3651 10591
rect 3801 10557 3835 10591
rect 3893 10557 3927 10591
rect 4537 10557 4571 10591
rect 4629 10557 4663 10591
rect 6837 10557 6871 10591
rect 7113 10557 7147 10591
rect 7593 10557 7627 10591
rect 7941 10557 7975 10591
rect 8493 10557 8527 10591
rect 8861 10557 8895 10591
rect 9873 10557 9907 10591
rect 11345 10557 11379 10591
rect 11897 10557 11931 10591
rect 7757 10489 7791 10523
rect 9321 10489 9355 10523
rect 3433 10421 3467 10455
rect 4261 10421 4295 10455
rect 5089 10421 5123 10455
rect 5825 10421 5859 10455
rect 10517 10421 10551 10455
rect 11713 10421 11747 10455
rect 1961 10217 1995 10251
rect 2329 10217 2363 10251
rect 2513 10217 2547 10251
rect 4537 10217 4571 10251
rect 6929 10217 6963 10251
rect 8033 10217 8067 10251
rect 8309 10217 8343 10251
rect 8677 10217 8711 10251
rect 10517 10217 10551 10251
rect 6377 10149 6411 10183
rect 10425 10149 10459 10183
rect 11805 10149 11839 10183
rect 13093 10149 13127 10183
rect 4261 10081 4295 10115
rect 7205 10081 7239 10115
rect 7665 10081 7699 10115
rect 11713 10081 11747 10115
rect 2053 10013 2087 10047
rect 2145 10013 2179 10047
rect 3249 10013 3283 10047
rect 3341 10013 3375 10047
rect 3525 10013 3559 10047
rect 3617 10013 3651 10047
rect 4169 10013 4203 10047
rect 4721 10013 4755 10047
rect 4905 10013 4939 10047
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 6198 10013 6232 10047
rect 6837 10013 6871 10047
rect 7297 10013 7331 10047
rect 7757 10013 7791 10047
rect 8493 10013 8527 10047
rect 8769 10013 8803 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 9965 10013 9999 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 10701 10013 10735 10047
rect 11437 10013 11471 10047
rect 12265 10013 12299 10047
rect 12633 10013 12667 10047
rect 13461 10013 13495 10047
rect 5641 9945 5675 9979
rect 6009 9945 6043 9979
rect 6101 9945 6135 9979
rect 7941 9945 7975 9979
rect 9045 9945 9079 9979
rect 11621 9945 11655 9979
rect 13185 9945 13219 9979
rect 3065 9877 3099 9911
rect 6653 9877 6687 9911
rect 13277 9877 13311 9911
rect 8125 9673 8159 9707
rect 8861 9673 8895 9707
rect 3801 9605 3835 9639
rect 6653 9605 6687 9639
rect 8677 9605 8711 9639
rect 10701 9605 10735 9639
rect 10885 9605 10919 9639
rect 11069 9605 11103 9639
rect 12909 9605 12943 9639
rect 3612 9537 3646 9571
rect 3709 9537 3743 9571
rect 3985 9537 4019 9571
rect 4452 9537 4486 9571
rect 4721 9537 4755 9571
rect 4905 9537 4939 9571
rect 4997 9537 5031 9571
rect 5141 9537 5175 9571
rect 6009 9537 6043 9571
rect 8309 9537 8343 9571
rect 8493 9537 8527 9571
rect 8769 9537 8803 9571
rect 9137 9537 9171 9571
rect 10149 9537 10183 9571
rect 11529 9537 11563 9571
rect 12173 9537 12207 9571
rect 12449 9537 12483 9571
rect 13277 9537 13311 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3157 9469 3191 9503
rect 4077 9469 4111 9503
rect 4353 9469 4387 9503
rect 6377 9469 6411 9503
rect 12725 9469 12759 9503
rect 3433 9401 3467 9435
rect 6193 9401 6227 9435
rect 12541 9401 12575 9435
rect 13461 9401 13495 9435
rect 5273 9333 5307 9367
rect 5825 9333 5859 9367
rect 13093 9333 13127 9367
rect 2237 9129 2271 9163
rect 3525 9129 3559 9163
rect 6653 9129 6687 9163
rect 6929 9129 6963 9163
rect 8769 9129 8803 9163
rect 9689 9129 9723 9163
rect 1961 9061 1995 9095
rect 2421 9061 2455 9095
rect 4077 9061 4111 9095
rect 10333 9061 10367 9095
rect 12817 9061 12851 9095
rect 5181 8993 5215 9027
rect 9045 8993 9079 9027
rect 9873 8993 9907 9027
rect 11437 8993 11471 9027
rect 1961 8925 1995 8959
rect 2053 8925 2087 8959
rect 3433 8925 3467 8959
rect 3801 8925 3835 8959
rect 4905 8925 4939 8959
rect 6837 8925 6871 8959
rect 7481 8925 7515 8959
rect 10885 8925 10919 8959
rect 11529 8925 11563 8959
rect 12725 8925 12759 8959
rect 13461 8925 13495 8959
rect 7941 8857 7975 8891
rect 8033 8857 8067 8891
rect 10425 8857 10459 8891
rect 10609 8857 10643 8891
rect 11345 8857 11379 8891
rect 13185 8857 13219 8891
rect 3985 8789 4019 8823
rect 8493 8789 8527 8823
rect 9229 8789 9263 8823
rect 9321 8789 9355 8823
rect 10517 8789 10551 8823
rect 13277 8789 13311 8823
rect 4629 8585 4663 8619
rect 5733 8585 5767 8619
rect 6101 8585 6135 8619
rect 8861 8585 8895 8619
rect 11529 8585 11563 8619
rect 12817 8585 12851 8619
rect 2329 8517 2363 8551
rect 3157 8517 3191 8551
rect 6377 8517 6411 8551
rect 8585 8517 8619 8551
rect 8769 8517 8803 8551
rect 9045 8517 9079 8551
rect 9689 8517 9723 8551
rect 10517 8517 10551 8551
rect 10793 8517 10827 8551
rect 11345 8517 11379 8551
rect 11989 8517 12023 8551
rect 12541 8517 12575 8551
rect 1777 8449 1811 8483
rect 1869 8449 1903 8483
rect 2145 8449 2179 8483
rect 2421 8449 2455 8483
rect 2565 8449 2599 8483
rect 5641 8449 5675 8483
rect 5917 8449 5951 8483
rect 7021 8449 7055 8483
rect 8125 8449 8159 8483
rect 9229 8449 9263 8483
rect 9873 8449 9907 8483
rect 11069 8449 11103 8483
rect 11897 8449 11931 8483
rect 13185 8449 13219 8483
rect 2881 8381 2915 8415
rect 9781 8381 9815 8415
rect 12081 8381 12115 8415
rect 13277 8381 13311 8415
rect 13369 8381 13403 8415
rect 2053 8313 2087 8347
rect 10885 8313 10919 8347
rect 12725 8313 12759 8347
rect 2697 8245 2731 8279
rect 1501 8041 1535 8075
rect 6653 8041 6687 8075
rect 7113 8041 7147 8075
rect 8769 8041 8803 8075
rect 9689 8041 9723 8075
rect 11621 8041 11655 8075
rect 12449 8041 12483 8075
rect 6929 7973 6963 8007
rect 8401 7973 8435 8007
rect 9229 7973 9263 8007
rect 10425 7973 10459 8007
rect 12265 7973 12299 8007
rect 3249 7905 3283 7939
rect 6101 7905 6135 7939
rect 7573 7905 7607 7939
rect 7757 7905 7791 7939
rect 11805 7905 11839 7939
rect 12357 7905 12391 7939
rect 13369 7905 13403 7939
rect 3433 7837 3467 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 7481 7837 7515 7871
rect 7941 7837 7975 7871
rect 8217 7837 8251 7871
rect 8309 7837 8343 7871
rect 8493 7837 8527 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 9873 7837 9907 7871
rect 10241 7837 10275 7871
rect 10977 7837 11011 7871
rect 11069 7837 11103 7871
rect 11437 7837 11471 7871
rect 12725 7837 12759 7871
rect 13277 7837 13311 7871
rect 2973 7769 3007 7803
rect 5365 7769 5399 7803
rect 13185 7769 13219 7803
rect 3617 7701 3651 7735
rect 3893 7701 3927 7735
rect 7021 7701 7055 7735
rect 10057 7701 10091 7735
rect 10149 7701 10183 7735
rect 10793 7701 10827 7735
rect 12817 7701 12851 7735
rect 14105 9877 14139 9911
rect 14105 7837 14139 7871
rect 3157 7497 3191 7531
rect 9413 7497 9447 7531
rect 10977 7497 11011 7531
rect 11345 7497 11379 7531
rect 11713 7497 11747 7531
rect 12817 7497 12851 7531
rect 14013 7497 14047 7531
rect 3525 7429 3559 7463
rect 6653 7429 6687 7463
rect 7849 7429 7883 7463
rect 11897 7429 11931 7463
rect 3341 7361 3375 7395
rect 3617 7361 3651 7395
rect 3714 7361 3748 7395
rect 4445 7361 4479 7395
rect 4628 7361 4662 7395
rect 4813 7361 4847 7395
rect 4997 7361 5031 7395
rect 5549 7361 5583 7395
rect 5917 7361 5951 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 7205 7361 7239 7395
rect 8125 7361 8159 7395
rect 8217 7361 8251 7395
rect 8309 7361 8343 7395
rect 8769 7361 8803 7395
rect 9137 7361 9171 7395
rect 9689 7361 9723 7395
rect 9873 7361 9907 7395
rect 10149 7361 10183 7395
rect 12357 7361 12391 7395
rect 12449 7361 12483 7395
rect 13185 7361 13219 7395
rect 13277 7361 13311 7395
rect 14013 7361 14047 7395
rect 1409 7293 1443 7327
rect 1685 7293 1719 7327
rect 4721 7293 4755 7327
rect 5457 7293 5491 7327
rect 9045 7293 9079 7327
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 12541 7293 12575 7327
rect 13369 7293 13403 7327
rect 3893 7225 3927 7259
rect 10057 7225 10091 7259
rect 4077 7157 4111 7191
rect 5089 7157 5123 7191
rect 5825 7157 5859 7191
rect 6101 7157 6135 7191
rect 6561 7157 6595 7191
rect 8861 7157 8895 7191
rect 8953 7157 8987 7191
rect 11989 7157 12023 7191
rect 2237 6953 2271 6987
rect 3433 6953 3467 6987
rect 4353 6953 4387 6987
rect 5720 6953 5754 6987
rect 10977 6953 11011 6987
rect 2329 6885 2363 6919
rect 3065 6885 3099 6919
rect 3801 6885 3835 6919
rect 4997 6885 5031 6919
rect 7849 6885 7883 6919
rect 9689 6885 9723 6919
rect 2053 6749 2087 6783
rect 2513 6749 2547 6783
rect 4629 6817 4663 6851
rect 8217 6817 8251 6851
rect 8585 6817 8619 6851
rect 10333 6817 10367 6851
rect 11713 6817 11747 6851
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4813 6749 4847 6783
rect 4905 6749 4939 6783
rect 5089 6749 5123 6783
rect 5457 6749 5491 6783
rect 7389 6749 7423 6783
rect 8401 6749 8435 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 9873 6749 9907 6783
rect 10149 6749 10183 6783
rect 11989 6749 12023 6783
rect 12909 6749 12943 6783
rect 2697 6681 2731 6715
rect 3065 6681 3099 6715
rect 7941 6681 7975 6715
rect 13553 6681 13587 6715
rect 2789 6613 2823 6647
rect 3249 6613 3283 6647
rect 3985 6613 4019 6647
rect 7205 6613 7239 6647
rect 10517 6613 10551 6647
rect 10609 6613 10643 6647
rect 11069 6613 11103 6647
rect 11437 6613 11471 6647
rect 11529 6613 11563 6647
rect 5733 6409 5767 6443
rect 6745 6409 6779 6443
rect 8401 6409 8435 6443
rect 11345 6409 11379 6443
rect 5365 6341 5399 6375
rect 5457 6341 5491 6375
rect 7849 6341 7883 6375
rect 9965 6341 9999 6375
rect 10149 6341 10183 6375
rect 10793 6341 10827 6375
rect 11161 6341 11195 6375
rect 12541 6341 12575 6375
rect 13093 6341 13127 6375
rect 13369 6341 13403 6375
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 3893 6273 3927 6307
rect 4077 6273 4111 6307
rect 4261 6273 4295 6307
rect 4537 6273 4571 6307
rect 4629 6273 4663 6307
rect 5089 6273 5123 6307
rect 5237 6273 5271 6307
rect 5595 6273 5629 6307
rect 6009 6273 6043 6307
rect 6837 6273 6871 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 7757 6273 7791 6307
rect 8217 6273 8251 6307
rect 8861 6273 8895 6307
rect 9229 6273 9263 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 10609 6273 10643 6307
rect 11621 6273 11655 6307
rect 12265 6273 12299 6307
rect 1409 6205 1443 6239
rect 1685 6205 1719 6239
rect 3709 6205 3743 6239
rect 7021 6205 7055 6239
rect 9045 6205 9079 6239
rect 12633 6205 12667 6239
rect 13185 6205 13219 6239
rect 9505 6137 9539 6171
rect 3157 6069 3191 6103
rect 4353 6069 4387 6103
rect 4813 6069 4847 6103
rect 6101 6069 6135 6103
rect 6377 6069 6411 6103
rect 7573 6069 7607 6103
rect 8033 6069 8067 6103
rect 8953 6069 8987 6103
rect 9137 6069 9171 6103
rect 10885 6069 10919 6103
rect 13461 6069 13495 6103
rect 2329 5865 2363 5899
rect 3249 5865 3283 5899
rect 4629 5865 4663 5899
rect 4813 5865 4847 5899
rect 5181 5865 5215 5899
rect 6653 5865 6687 5899
rect 7297 5865 7331 5899
rect 9505 5865 9539 5899
rect 9689 5865 9723 5899
rect 9873 5865 9907 5899
rect 10425 5865 10459 5899
rect 12817 5865 12851 5899
rect 13277 5865 13311 5899
rect 13553 5865 13587 5899
rect 14013 5865 14047 5899
rect 3525 5797 3559 5831
rect 6193 5797 6227 5831
rect 6929 5797 6963 5831
rect 7481 5797 7515 5831
rect 8125 5797 8159 5831
rect 8677 5797 8711 5831
rect 8769 5797 8803 5831
rect 9045 5797 9079 5831
rect 11529 5797 11563 5831
rect 12173 5797 12207 5831
rect 2973 5729 3007 5763
rect 3893 5729 3927 5763
rect 4353 5729 4387 5763
rect 4537 5729 4571 5763
rect 5641 5729 5675 5763
rect 6377 5729 6411 5763
rect 8217 5729 8251 5763
rect 2145 5661 2179 5695
rect 2881 5661 2915 5695
rect 3433 5661 3467 5695
rect 3985 5661 4019 5695
rect 4445 5661 4479 5695
rect 5549 5661 5583 5695
rect 6193 5661 6227 5695
rect 6561 5661 6595 5695
rect 7205 5661 7239 5695
rect 7297 5661 7331 5695
rect 7389 5661 7423 5695
rect 8033 5661 8067 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 5825 5593 5859 5627
rect 10977 5729 11011 5763
rect 9229 5661 9263 5695
rect 9321 5661 9355 5695
rect 9873 5661 9907 5695
rect 10057 5661 10091 5695
rect 10333 5661 10367 5695
rect 11253 5661 11287 5695
rect 11437 5661 11471 5695
rect 11713 5661 11747 5695
rect 12633 5661 12667 5695
rect 9505 5593 9539 5627
rect 12265 5593 12299 5627
rect 12725 5593 12759 5627
rect 13185 5593 13219 5627
rect 2421 5525 2455 5559
rect 7849 5525 7883 5559
rect 8769 5525 8803 5559
rect 10241 5525 10275 5559
rect 10793 5525 10827 5559
rect 10885 5525 10919 5559
rect 12449 5525 12483 5559
rect 13001 5525 13035 5559
rect 1501 5321 1535 5355
rect 3893 5321 3927 5355
rect 5549 5321 5583 5355
rect 7849 5321 7883 5355
rect 8677 5321 8711 5355
rect 11345 5321 11379 5355
rect 6469 5253 6503 5287
rect 7021 5253 7055 5287
rect 9689 5253 9723 5287
rect 10977 5253 11011 5287
rect 3801 5185 3835 5219
rect 4169 5185 4203 5219
rect 4353 5185 4387 5219
rect 4905 5185 4939 5219
rect 4997 5185 5031 5219
rect 5365 5185 5399 5219
rect 5457 5185 5491 5219
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 6653 5185 6687 5219
rect 6837 5185 6871 5219
rect 7389 5185 7423 5219
rect 8932 5185 8966 5219
rect 9413 5185 9447 5219
rect 9873 5185 9907 5219
rect 10148 5185 10182 5219
rect 10333 5185 10367 5219
rect 10885 5185 10919 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 13461 5185 13495 5219
rect 2973 5117 3007 5151
rect 3249 5117 3283 5151
rect 5089 5117 5123 5151
rect 5181 5117 5215 5151
rect 7941 5117 7975 5151
rect 8125 5117 8159 5151
rect 9229 5117 9263 5151
rect 10057 5117 10091 5151
rect 10701 5117 10735 5151
rect 4537 5049 4571 5083
rect 5917 5049 5951 5083
rect 7481 5049 7515 5083
rect 8493 5049 8527 5083
rect 9137 5049 9171 5083
rect 9965 5049 9999 5083
rect 13277 5049 13311 5083
rect 4721 4981 4755 5015
rect 7297 4981 7331 5015
rect 9045 4981 9079 5015
rect 10517 4981 10551 5015
rect 11805 4981 11839 5015
rect 2053 4777 2087 4811
rect 2973 4777 3007 4811
rect 4629 4777 4663 4811
rect 6469 4777 6503 4811
rect 7941 4777 7975 4811
rect 8033 4777 8067 4811
rect 9229 4777 9263 4811
rect 6009 4709 6043 4743
rect 7849 4709 7883 4743
rect 8401 4709 8435 4743
rect 9505 4709 9539 4743
rect 10425 4709 10459 4743
rect 13093 4709 13127 4743
rect 2697 4641 2731 4675
rect 3065 4641 3099 4675
rect 3525 4641 3559 4675
rect 4241 4641 4275 4675
rect 4537 4641 4571 4675
rect 5089 4641 5123 4675
rect 6653 4641 6687 4675
rect 9597 4641 9631 4675
rect 10885 4641 10919 4675
rect 11345 4641 11379 4675
rect 12633 4641 12667 4675
rect 13185 4641 13219 4675
rect 1869 4573 1903 4607
rect 2329 4573 2363 4607
rect 2605 4573 2639 4607
rect 3433 4573 3467 4607
rect 4997 4573 5031 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6285 4573 6319 4607
rect 6745 4573 6779 4607
rect 6837 4573 6871 4607
rect 6929 4573 6963 4607
rect 7113 4573 7147 4607
rect 7389 4573 7423 4607
rect 7757 4573 7791 4607
rect 8146 4573 8180 4607
rect 8585 4573 8619 4607
rect 9413 4573 9447 4607
rect 9689 4573 9723 4607
rect 9873 4573 9907 4607
rect 10241 4573 10275 4607
rect 10333 4573 10367 4607
rect 10517 4573 10551 4607
rect 10701 4573 10735 4607
rect 11529 4573 11563 4607
rect 12173 4573 12207 4607
rect 12449 4573 12483 4607
rect 13461 4573 13495 4607
rect 3801 4505 3835 4539
rect 3985 4505 4019 4539
rect 7205 4505 7239 4539
rect 7573 4505 7607 4539
rect 8677 4505 8711 4539
rect 11437 4505 11471 4539
rect 1777 4437 1811 4471
rect 2237 4437 2271 4471
rect 4353 4437 4387 4471
rect 4445 4437 4479 4471
rect 10057 4437 10091 4471
rect 13277 4437 13311 4471
rect 5181 4233 5215 4267
rect 5641 4233 5675 4267
rect 6101 4233 6135 4267
rect 8493 4233 8527 4267
rect 3341 4165 3375 4199
rect 9689 4165 9723 4199
rect 9873 4165 9907 4199
rect 10333 4165 10367 4199
rect 10517 4165 10551 4199
rect 13277 4165 13311 4199
rect 2237 4097 2271 4131
rect 3065 4097 3099 4131
rect 3985 4097 4019 4131
rect 4169 4097 4203 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 4813 4097 4847 4131
rect 4905 4097 4939 4131
rect 5549 4097 5583 4131
rect 6009 4097 6043 4131
rect 6745 4097 6779 4131
rect 7389 4097 7423 4131
rect 7849 4097 7883 4131
rect 8953 4097 8987 4131
rect 9505 4097 9539 4131
rect 9597 4097 9631 4131
rect 11253 4097 11287 4131
rect 11529 4097 11563 4131
rect 11897 4097 11931 4131
rect 12817 4097 12851 4131
rect 2953 4029 2987 4063
rect 3433 4029 3467 4063
rect 5733 4029 5767 4063
rect 6377 4029 6411 4063
rect 6653 4029 6687 4063
rect 7297 4029 7331 4063
rect 8309 4029 8343 4063
rect 8401 4029 8435 4063
rect 9137 4029 9171 4063
rect 12173 4029 12207 4063
rect 12725 4029 12759 4063
rect 12909 4029 12943 4063
rect 2605 3961 2639 3995
rect 4077 3961 4111 3995
rect 4629 3961 4663 3995
rect 8861 3961 8895 3995
rect 10701 3961 10735 3995
rect 12633 3961 12667 3995
rect 2421 3893 2455 3927
rect 2789 3893 2823 3927
rect 4997 3893 5031 3927
rect 7021 3893 7055 3927
rect 7665 3893 7699 3927
rect 7941 3893 7975 3927
rect 9873 3893 9907 3927
rect 10057 3893 10091 3927
rect 12081 3893 12115 3927
rect 13185 3893 13219 3927
rect 3249 3689 3283 3723
rect 4169 3689 4203 3723
rect 4997 3689 5031 3723
rect 9689 3689 9723 3723
rect 10153 3621 10187 3655
rect 10517 3621 10551 3655
rect 13277 3621 13311 3655
rect 1777 3553 1811 3587
rect 5181 3553 5215 3587
rect 5457 3553 5491 3587
rect 6561 3553 6595 3587
rect 8033 3553 8067 3587
rect 9045 3553 9079 3587
rect 10241 3553 10275 3587
rect 1501 3485 1535 3519
rect 4261 3485 4295 3519
rect 4353 3485 4387 3519
rect 4446 3485 4480 3519
rect 4721 3485 4755 3519
rect 4857 3485 4891 3519
rect 5549 3485 5583 3519
rect 6285 3485 6319 3519
rect 8513 3485 8547 3519
rect 8769 3485 8803 3519
rect 10057 3485 10091 3519
rect 10346 3485 10380 3519
rect 10977 3485 11011 3519
rect 11713 3485 11747 3519
rect 11989 3485 12023 3519
rect 13185 3485 13219 3519
rect 4629 3417 4663 3451
rect 8217 3417 8251 3451
rect 8401 3417 8435 3451
rect 10701 3417 10735 3451
rect 10885 3417 10919 3451
rect 11897 3417 11931 3451
rect 8585 3349 8619 3383
rect 9229 3349 9263 3383
rect 9321 3349 9355 3383
rect 9873 3349 9907 3383
rect 1593 3145 1627 3179
rect 3801 3145 3835 3179
rect 8033 3145 8067 3179
rect 8769 3145 8803 3179
rect 9321 3145 9355 3179
rect 11161 3145 11195 3179
rect 12173 3145 12207 3179
rect 4261 3077 4295 3111
rect 8677 3077 8711 3111
rect 9965 3077 9999 3111
rect 10149 3077 10183 3111
rect 12081 3077 12115 3111
rect 1777 3009 1811 3043
rect 2053 3009 2087 3043
rect 3985 3009 4019 3043
rect 6377 3009 6411 3043
rect 7021 3009 7055 3043
rect 7389 3009 7423 3043
rect 7573 3009 7607 3043
rect 8125 3009 8159 3043
rect 9045 3009 9079 3043
rect 9505 3009 9539 3043
rect 9781 3009 9815 3043
rect 10333 3009 10367 3043
rect 10793 3009 10827 3043
rect 11529 3009 11563 3043
rect 11989 3009 12023 3043
rect 12541 3009 12575 3043
rect 2329 2941 2363 2975
rect 6929 2941 6963 2975
rect 7113 2941 7147 2975
rect 8309 2941 8343 2975
rect 9601 2941 9635 2975
rect 10609 2941 10643 2975
rect 10701 2941 10735 2975
rect 11253 2941 11287 2975
rect 12633 2941 12667 2975
rect 12725 2941 12759 2975
rect 13185 2941 13219 2975
rect 5733 2873 5767 2907
rect 6837 2873 6871 2907
rect 9689 2873 9723 2907
rect 7665 2805 7699 2839
rect 13001 2805 13035 2839
rect 13461 2805 13495 2839
rect 14013 2805 14047 2839
rect 3065 2601 3099 2635
rect 4077 2601 4111 2635
rect 4905 2601 4939 2635
rect 5089 2601 5123 2635
rect 8401 2601 8435 2635
rect 8493 2601 8527 2635
rect 10701 2601 10735 2635
rect 7205 2533 7239 2567
rect 10977 2533 11011 2567
rect 11253 2533 11287 2567
rect 11437 2533 11471 2567
rect 4537 2465 4571 2499
rect 7757 2465 7791 2499
rect 9505 2465 9539 2499
rect 11897 2465 11931 2499
rect 12081 2465 12115 2499
rect 2881 2397 2915 2431
rect 3249 2397 3283 2431
rect 3617 2397 3651 2431
rect 3801 2397 3835 2431
rect 4445 2397 4479 2431
rect 4721 2397 4755 2431
rect 5641 2397 5675 2431
rect 5733 2397 5767 2431
rect 7205 2397 7239 2431
rect 7481 2397 7515 2431
rect 7665 2397 7699 2431
rect 7849 2397 7883 2431
rect 8217 2397 8251 2431
rect 9321 2397 9355 2431
rect 9781 2397 9815 2431
rect 10517 2397 10551 2431
rect 11621 2397 11655 2431
rect 12173 2397 12207 2431
rect 12633 2397 12667 2431
rect 13461 2397 13495 2431
rect 10241 2329 10275 2363
rect 10333 2329 10367 2363
rect 13093 2329 13127 2363
rect 13185 2329 13219 2363
rect 3985 2261 4019 2295
rect 5457 2261 5491 2295
rect 8217 2261 8251 2295
rect 8953 2261 8987 2295
rect 9413 2261 9447 2295
rect 10885 2261 10919 2295
rect 12541 2261 12575 2295
rect 13369 2261 13403 2295
rect 3157 2057 3191 2091
rect 5089 2057 5123 2091
rect 10977 2057 11011 2091
rect 11345 2057 11379 2091
rect 13185 2057 13219 2091
rect 3617 1989 3651 2023
rect 6009 1989 6043 2023
rect 7573 1989 7607 2023
rect 7757 1989 7791 2023
rect 10517 1989 10551 2023
rect 13461 1989 13495 2023
rect 1409 1921 1443 1955
rect 5273 1921 5307 1955
rect 6193 1921 6227 1955
rect 6469 1921 6503 1955
rect 7941 1921 7975 1955
rect 9413 1921 9447 1955
rect 9597 1921 9631 1955
rect 10241 1921 10275 1955
rect 11529 1921 11563 1955
rect 13001 1921 13035 1955
rect 13369 1921 13403 1955
rect 1685 1853 1719 1887
rect 3341 1853 3375 1887
rect 10701 1853 10735 1887
rect 10885 1853 10919 1887
rect 9229 1785 9263 1819
rect 12817 1785 12851 1819
rect 6469 1717 6503 1751
rect 2237 1513 2271 1547
rect 3157 1513 3191 1547
rect 7849 1513 7883 1547
rect 9873 1513 9907 1547
rect 10701 1513 10735 1547
rect 6837 1445 6871 1479
rect 9413 1445 9447 1479
rect 5365 1377 5399 1411
rect 5641 1377 5675 1411
rect 8217 1377 8251 1411
rect 8953 1377 8987 1411
rect 10517 1377 10551 1411
rect 11161 1377 11195 1411
rect 11529 1377 11563 1411
rect 2053 1309 2087 1343
rect 2421 1309 2455 1343
rect 2881 1309 2915 1343
rect 3341 1309 3375 1343
rect 6377 1309 6411 1343
rect 7205 1309 7239 1343
rect 7297 1309 7331 1343
rect 7481 1309 7515 1343
rect 7665 1309 7699 1343
rect 7941 1309 7975 1343
rect 8677 1309 8711 1343
rect 9781 1309 9815 1343
rect 10885 1309 10919 1343
rect 11989 1309 12023 1343
rect 12449 1309 12483 1343
rect 13093 1309 13127 1343
rect 13369 1309 13403 1343
rect 6929 1241 6963 1275
rect 8125 1241 8159 1275
rect 9505 1241 9539 1275
rect 9597 1241 9631 1275
rect 10333 1241 10367 1275
rect 11069 1241 11103 1275
rect 12081 1241 12115 1275
rect 12173 1241 12207 1275
rect 12357 1241 12391 1275
rect 3065 1173 3099 1207
rect 3893 1173 3927 1207
rect 7021 1173 7055 1207
rect 8585 1173 8619 1207
rect 10241 1173 10275 1207
rect 14013 493 14047 527
<< metal1 >>
rect 1104 13626 13892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 13892 13626
rect 1104 13552 13892 13574
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 3559 13484 3893 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3881 13481 3893 13484
rect 3927 13512 3939 13515
rect 5534 13512 5540 13524
rect 3927 13484 5540 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3418 13308 3424 13320
rect 3191 13280 3424 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3418 13268 3424 13280
rect 3476 13308 3482 13320
rect 3528 13308 3556 13475
rect 5534 13472 5540 13484
rect 5592 13512 5598 13524
rect 6181 13515 6239 13521
rect 6181 13512 6193 13515
rect 5592 13484 6193 13512
rect 5592 13472 5598 13484
rect 6181 13481 6193 13484
rect 6227 13512 6239 13515
rect 6227 13484 7052 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 6914 13444 6920 13456
rect 6875 13416 6920 13444
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 7024 13444 7052 13484
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 8481 13515 8539 13521
rect 8481 13512 8493 13515
rect 8260 13484 8493 13512
rect 8260 13472 8266 13484
rect 8481 13481 8493 13484
rect 8527 13481 8539 13515
rect 8481 13475 8539 13481
rect 8297 13447 8355 13453
rect 8297 13444 8309 13447
rect 7024 13416 8309 13444
rect 8297 13413 8309 13416
rect 8343 13413 8355 13447
rect 8297 13407 8355 13413
rect 9677 13447 9735 13453
rect 9677 13413 9689 13447
rect 9723 13444 9735 13447
rect 9766 13444 9772 13456
rect 9723 13416 9772 13444
rect 9723 13413 9735 13416
rect 9677 13407 9735 13413
rect 9766 13404 9772 13416
rect 9824 13444 9830 13456
rect 9824 13416 10272 13444
rect 9824 13404 9830 13416
rect 5902 13336 5908 13388
rect 5960 13376 5966 13388
rect 5960 13348 6781 13376
rect 5960 13336 5966 13348
rect 3476 13280 3556 13308
rect 5261 13311 5319 13317
rect 3476 13268 3482 13280
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5994 13308 6000 13320
rect 5307 13280 6000 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5994 13268 6000 13280
rect 6052 13268 6058 13320
rect 6753 13317 6781 13348
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 10244 13385 10272 13416
rect 8665 13379 8723 13385
rect 8665 13376 8677 13379
rect 6880 13348 8677 13376
rect 6880 13336 6886 13348
rect 8665 13345 8677 13348
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13376 9183 13379
rect 10229 13379 10287 13385
rect 9171 13348 9904 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 6738 13311 6796 13317
rect 6738 13277 6750 13311
rect 6784 13277 6796 13311
rect 7101 13311 7159 13317
rect 7101 13308 7113 13311
rect 6738 13271 6796 13277
rect 6932 13280 7113 13308
rect 5166 13200 5172 13252
rect 5224 13240 5230 13252
rect 6380 13240 6408 13271
rect 6546 13240 6552 13252
rect 5224 13212 6408 13240
rect 6507 13212 6552 13240
rect 5224 13200 5230 13212
rect 6546 13200 6552 13212
rect 6604 13200 6610 13252
rect 6641 13243 6699 13249
rect 6641 13209 6653 13243
rect 6687 13240 6699 13243
rect 6822 13240 6828 13252
rect 6687 13212 6828 13240
rect 6687 13209 6699 13212
rect 6641 13203 6699 13209
rect 6822 13200 6828 13212
rect 6880 13200 6886 13252
rect 3326 13172 3332 13184
rect 3287 13144 3332 13172
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 5350 13172 5356 13184
rect 5311 13144 5356 13172
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 6564 13172 6592 13200
rect 6932 13172 6960 13280
rect 7101 13277 7113 13280
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 7377 13311 7435 13317
rect 7377 13277 7389 13311
rect 7423 13308 7435 13311
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7423 13280 7757 13308
rect 7423 13277 7435 13280
rect 7377 13271 7435 13277
rect 7745 13277 7757 13280
rect 7791 13308 7803 13311
rect 7926 13308 7932 13320
rect 7791 13280 7932 13308
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8680 13308 8708 13339
rect 9217 13311 9275 13317
rect 9217 13308 9229 13311
rect 8680 13280 9229 13308
rect 9217 13277 9229 13280
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 6564 13144 6960 13172
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 7193 13175 7251 13181
rect 7193 13172 7205 13175
rect 7064 13144 7205 13172
rect 7064 13132 7070 13144
rect 7193 13141 7205 13144
rect 7239 13141 7251 13175
rect 7193 13135 7251 13141
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 7653 13175 7711 13181
rect 7653 13172 7665 13175
rect 7616 13144 7665 13172
rect 7616 13132 7622 13144
rect 7653 13141 7665 13144
rect 7699 13141 7711 13175
rect 7653 13135 7711 13141
rect 8205 13175 8263 13181
rect 8205 13141 8217 13175
rect 8251 13172 8263 13175
rect 8297 13175 8355 13181
rect 8297 13172 8309 13175
rect 8251 13144 8309 13172
rect 8251 13141 8263 13144
rect 8205 13135 8263 13141
rect 8297 13141 8309 13144
rect 8343 13172 8355 13175
rect 8570 13172 8576 13184
rect 8343 13144 8576 13172
rect 8343 13141 8355 13144
rect 8297 13135 8355 13141
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 9309 13175 9367 13181
rect 9309 13141 9321 13175
rect 9355 13172 9367 13175
rect 9490 13172 9496 13184
rect 9355 13144 9496 13172
rect 9355 13141 9367 13144
rect 9309 13135 9367 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 9876 13181 9904 13348
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13308 10747 13311
rect 11330 13308 11336 13320
rect 10735 13280 11336 13308
rect 10735 13277 10747 13280
rect 10689 13271 10747 13277
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 12066 13308 12072 13320
rect 12027 13280 12072 13308
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12710 13308 12716 13320
rect 12671 13280 12716 13308
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 10781 13243 10839 13249
rect 10781 13209 10793 13243
rect 10827 13240 10839 13243
rect 10873 13243 10931 13249
rect 10873 13240 10885 13243
rect 10827 13212 10885 13240
rect 10827 13209 10839 13212
rect 10781 13203 10839 13209
rect 10873 13209 10885 13212
rect 10919 13209 10931 13243
rect 12526 13240 12532 13252
rect 12487 13212 12532 13240
rect 10873 13203 10931 13209
rect 12526 13200 12532 13212
rect 12584 13200 12590 13252
rect 12618 13200 12624 13252
rect 12676 13240 12682 13252
rect 13170 13240 13176 13252
rect 12676 13212 12721 13240
rect 13131 13212 13176 13240
rect 12676 13200 12682 13212
rect 13170 13200 13176 13212
rect 13228 13200 13234 13252
rect 13265 13243 13323 13249
rect 13265 13209 13277 13243
rect 13311 13240 13323 13243
rect 13354 13240 13360 13252
rect 13311 13212 13360 13240
rect 13311 13209 13323 13212
rect 13265 13203 13323 13209
rect 13354 13200 13360 13212
rect 13412 13200 13418 13252
rect 9861 13175 9919 13181
rect 9861 13141 9873 13175
rect 9907 13172 9919 13175
rect 10042 13172 10048 13184
rect 9907 13144 10048 13172
rect 9907 13141 9919 13144
rect 9861 13135 9919 13141
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 11054 13172 11060 13184
rect 11015 13144 11060 13172
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 1104 13082 13892 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 13892 13082
rect 1104 13008 13892 13030
rect 2498 12968 2504 12980
rect 2332 12940 2504 12968
rect 2332 12841 2360 12940
rect 2498 12928 2504 12940
rect 2556 12968 2562 12980
rect 4065 12971 4123 12977
rect 2556 12940 4016 12968
rect 2556 12928 2562 12940
rect 3326 12860 3332 12912
rect 3384 12860 3390 12912
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3988 12696 4016 12940
rect 4065 12937 4077 12971
rect 4111 12968 4123 12971
rect 4706 12968 4712 12980
rect 4111 12940 4712 12968
rect 4111 12937 4123 12940
rect 4065 12931 4123 12937
rect 4706 12928 4712 12940
rect 4764 12968 4770 12980
rect 5994 12968 6000 12980
rect 4764 12940 5856 12968
rect 5955 12940 6000 12968
rect 4764 12928 4770 12940
rect 5534 12860 5540 12912
rect 5592 12860 5598 12912
rect 5828 12900 5856 12940
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 7926 12968 7932 12980
rect 6880 12940 7932 12968
rect 6880 12928 6886 12940
rect 7926 12928 7932 12940
rect 7984 12968 7990 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 7984 12940 8125 12968
rect 7984 12928 7990 12940
rect 8113 12937 8125 12940
rect 8159 12937 8171 12971
rect 8113 12931 8171 12937
rect 8297 12971 8355 12977
rect 8297 12937 8309 12971
rect 8343 12937 8355 12971
rect 8297 12931 8355 12937
rect 9401 12971 9459 12977
rect 9401 12937 9413 12971
rect 9447 12968 9459 12971
rect 12066 12968 12072 12980
rect 9447 12940 12072 12968
rect 9447 12937 9459 12940
rect 9401 12931 9459 12937
rect 6546 12900 6552 12912
rect 5828 12872 6552 12900
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 6641 12903 6699 12909
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 6914 12900 6920 12912
rect 6687 12872 6920 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 8312 12900 8340 12931
rect 8941 12903 8999 12909
rect 8941 12900 8953 12903
rect 7866 12872 8340 12900
rect 8404 12872 8953 12900
rect 8110 12792 8116 12844
rect 8168 12832 8174 12844
rect 8404 12832 8432 12872
rect 8941 12869 8953 12872
rect 8987 12869 8999 12903
rect 11330 12900 11336 12912
rect 11291 12872 11336 12900
rect 8941 12863 8999 12869
rect 11330 12860 11336 12872
rect 11388 12860 11394 12912
rect 8168 12804 8432 12832
rect 8481 12835 8539 12841
rect 8168 12792 8174 12804
rect 8481 12801 8493 12835
rect 8527 12832 8539 12835
rect 8570 12832 8576 12844
rect 8527 12804 8576 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9122 12832 9128 12844
rect 9079 12804 9128 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 9766 12832 9772 12844
rect 9727 12804 9772 12832
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 11238 12832 11244 12844
rect 11199 12804 11244 12832
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11716 12841 11744 12940
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 13354 12968 13360 12980
rect 13315 12940 13360 12968
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 12894 12832 12900 12844
rect 12855 12804 12900 12832
rect 11701 12795 11759 12801
rect 12894 12792 12900 12804
rect 12952 12832 12958 12844
rect 13541 12835 13599 12841
rect 13541 12832 13553 12835
rect 12952 12804 13553 12832
rect 12952 12792 12958 12804
rect 13541 12801 13553 12804
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 4614 12764 4620 12776
rect 4571 12736 4620 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 4264 12696 4292 12727
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 6365 12767 6423 12773
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6365 12727 6423 12733
rect 8849 12767 8907 12773
rect 8849 12733 8861 12767
rect 8895 12764 8907 12767
rect 10042 12764 10048 12776
rect 8895 12736 10048 12764
rect 8895 12733 8907 12736
rect 8849 12727 8907 12733
rect 3988 12668 4292 12696
rect 4264 12628 4292 12668
rect 6380 12628 6408 12727
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 8386 12656 8392 12708
rect 8444 12696 8450 12708
rect 9214 12696 9220 12708
rect 8444 12668 9220 12696
rect 8444 12656 8450 12668
rect 9214 12656 9220 12668
rect 9272 12696 9278 12708
rect 9493 12699 9551 12705
rect 9493 12696 9505 12699
rect 9272 12668 9505 12696
rect 9272 12656 9278 12668
rect 9493 12665 9505 12668
rect 9539 12665 9551 12699
rect 9493 12659 9551 12665
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12986 12696 12992 12708
rect 12584 12668 12992 12696
rect 12584 12656 12590 12668
rect 12986 12656 12992 12668
rect 13044 12656 13050 12708
rect 4264 12600 6408 12628
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 10870 12628 10876 12640
rect 10100 12600 10876 12628
rect 10100 12588 10106 12600
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 1104 12538 13892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 13892 12538
rect 1104 12464 13892 12486
rect 4614 12424 4620 12436
rect 4575 12396 4620 12424
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 5902 12384 5908 12436
rect 5960 12384 5966 12436
rect 10134 12424 10140 12436
rect 10095 12396 10140 12424
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 11609 12427 11667 12433
rect 11609 12424 11621 12427
rect 10928 12396 11621 12424
rect 10928 12384 10934 12396
rect 11609 12393 11621 12396
rect 11655 12393 11667 12427
rect 11609 12387 11667 12393
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 13357 12427 13415 12433
rect 13357 12424 13369 12427
rect 12676 12396 13369 12424
rect 12676 12384 12682 12396
rect 13357 12393 13369 12396
rect 13403 12393 13415 12427
rect 13357 12387 13415 12393
rect 3510 12316 3516 12368
rect 3568 12356 3574 12368
rect 3881 12359 3939 12365
rect 3881 12356 3893 12359
rect 3568 12328 3893 12356
rect 3568 12316 3574 12328
rect 3881 12325 3893 12328
rect 3927 12325 3939 12359
rect 5920 12356 5948 12384
rect 3881 12319 3939 12325
rect 5000 12328 5948 12356
rect 6549 12359 6607 12365
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 1719 12260 4261 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 1412 12096 1440 12183
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3418 12220 3424 12232
rect 3016 12192 3424 12220
rect 3016 12180 3022 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 4614 12220 4620 12232
rect 4111 12192 4620 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 2682 12112 2688 12164
rect 2740 12112 2746 12164
rect 3804 12152 3832 12183
rect 4614 12180 4620 12192
rect 4672 12220 4678 12232
rect 4796 12223 4854 12229
rect 4796 12220 4808 12223
rect 4672 12192 4808 12220
rect 4672 12180 4678 12192
rect 4796 12189 4808 12192
rect 4842 12220 4854 12223
rect 5000 12220 5028 12328
rect 6549 12325 6561 12359
rect 6595 12356 6607 12359
rect 9306 12356 9312 12368
rect 6595 12328 9312 12356
rect 6595 12325 6607 12328
rect 6549 12319 6607 12325
rect 9306 12316 9312 12328
rect 9364 12356 9370 12368
rect 12710 12356 12716 12368
rect 9364 12328 9628 12356
rect 9364 12316 9370 12328
rect 5350 12288 5356 12300
rect 5311 12260 5356 12288
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5813 12291 5871 12297
rect 5813 12257 5825 12291
rect 5859 12288 5871 12291
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5859 12260 5917 12288
rect 5859 12257 5871 12260
rect 5813 12251 5871 12257
rect 5905 12257 5917 12260
rect 5951 12288 5963 12291
rect 6385 12291 6443 12297
rect 6385 12288 6397 12291
rect 5951 12260 6397 12288
rect 5951 12257 5963 12260
rect 5905 12251 5963 12257
rect 6385 12257 6397 12260
rect 6431 12257 6443 12291
rect 6385 12251 6443 12257
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12288 7343 12291
rect 7558 12288 7564 12300
rect 7331 12260 7564 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8772 12260 9352 12288
rect 5166 12220 5172 12232
rect 4842 12192 5028 12220
rect 5127 12192 5172 12220
rect 4842 12189 4854 12192
rect 4796 12183 4854 12189
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5445 12223 5503 12229
rect 5445 12189 5457 12223
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 3160 12124 3832 12152
rect 4893 12155 4951 12161
rect 3160 12096 3188 12124
rect 4893 12121 4905 12155
rect 4939 12121 4951 12155
rect 4893 12115 4951 12121
rect 4985 12155 5043 12161
rect 4985 12121 4997 12155
rect 5031 12152 5043 12155
rect 5074 12152 5080 12164
rect 5031 12124 5080 12152
rect 5031 12121 5043 12124
rect 4985 12115 5043 12121
rect 1394 12084 1400 12096
rect 1307 12056 1400 12084
rect 1394 12044 1400 12056
rect 1452 12084 1458 12096
rect 2498 12084 2504 12096
rect 1452 12056 2504 12084
rect 1452 12044 1458 12056
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 3142 12084 3148 12096
rect 3055 12056 3148 12084
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 3878 12084 3884 12096
rect 3651 12056 3884 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4908 12084 4936 12115
rect 5074 12112 5080 12124
rect 5132 12152 5138 12164
rect 5460 12152 5488 12183
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5592 12192 6009 12220
rect 5592 12180 5598 12192
rect 5997 12189 6009 12192
rect 6043 12220 6055 12223
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 6043 12192 6285 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6273 12189 6285 12192
rect 6319 12220 6331 12223
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6319 12192 6837 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 7006 12220 7012 12232
rect 6967 12192 7012 12220
rect 6825 12183 6883 12189
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7101 12223 7159 12229
rect 7101 12189 7113 12223
rect 7147 12220 7159 12223
rect 7190 12220 7196 12232
rect 7147 12192 7196 12220
rect 7147 12189 7159 12192
rect 7101 12183 7159 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12220 7435 12223
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7423 12192 7665 12220
rect 7423 12189 7435 12192
rect 7377 12183 7435 12189
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 7653 12183 7711 12189
rect 5132 12124 5488 12152
rect 5132 12112 5138 12124
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 7392 12152 7420 12183
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 6788 12124 7420 12152
rect 8113 12155 8171 12161
rect 6788 12112 6794 12124
rect 8113 12121 8125 12155
rect 8159 12121 8171 12155
rect 8496 12152 8524 12183
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 8772 12229 8800 12260
rect 8757 12223 8815 12229
rect 8628 12192 8673 12220
rect 8628 12180 8634 12192
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12189 8999 12223
rect 9214 12220 9220 12232
rect 9127 12192 9220 12220
rect 8941 12183 8999 12189
rect 8662 12152 8668 12164
rect 8496 12124 8668 12152
rect 8113 12115 8171 12121
rect 5994 12084 6000 12096
rect 4908 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 8128 12084 8156 12115
rect 8662 12112 8668 12124
rect 8720 12152 8726 12164
rect 8956 12152 8984 12183
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 8720 12124 8984 12152
rect 8720 12112 8726 12124
rect 8754 12084 8760 12096
rect 8128 12056 8760 12084
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 9232 12084 9260 12180
rect 9324 12161 9352 12260
rect 9600 12229 9628 12328
rect 12406 12328 12716 12356
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 11388 12260 12020 12288
rect 11388 12248 11394 12260
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12189 9643 12223
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 9585 12183 9643 12189
rect 9309 12155 9367 12161
rect 9309 12121 9321 12155
rect 9355 12152 9367 12155
rect 9398 12152 9404 12164
rect 9355 12124 9404 12152
rect 9355 12121 9367 12124
rect 9309 12115 9367 12121
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 9508 12152 9536 12183
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11054 12220 11060 12232
rect 11015 12192 11060 12220
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 11238 12180 11244 12192
rect 11296 12220 11302 12232
rect 11992 12229 12020 12260
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11296 12192 11529 12220
rect 11296 12180 11302 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12253 12223 12311 12229
rect 12253 12189 12265 12223
rect 12299 12220 12311 12223
rect 12406 12220 12434 12328
rect 12710 12316 12716 12328
rect 12768 12356 12774 12368
rect 14001 12359 14059 12365
rect 14001 12356 14013 12359
rect 12768 12328 14013 12356
rect 12768 12316 12774 12328
rect 14001 12325 14013 12328
rect 14047 12325 14059 12359
rect 14001 12319 14059 12325
rect 13170 12248 13176 12300
rect 13228 12248 13234 12300
rect 12299 12192 12434 12220
rect 12989 12223 13047 12229
rect 12299 12189 12311 12192
rect 12253 12183 12311 12189
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13188 12220 13216 12248
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 13035 12192 13277 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 9674 12152 9680 12164
rect 9508 12124 9680 12152
rect 9674 12112 9680 12124
rect 9732 12152 9738 12164
rect 10134 12152 10140 12164
rect 9732 12124 10140 12152
rect 9732 12112 9738 12124
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 12161 12155 12219 12161
rect 12161 12121 12173 12155
rect 12207 12152 12219 12155
rect 12894 12152 12900 12164
rect 12207 12124 12900 12152
rect 12207 12121 12219 12124
rect 12161 12115 12219 12121
rect 12894 12112 12900 12124
rect 12952 12152 12958 12164
rect 13173 12155 13231 12161
rect 13173 12152 13185 12155
rect 12952 12124 13185 12152
rect 12952 12112 12958 12124
rect 13173 12121 13185 12124
rect 13219 12121 13231 12155
rect 13173 12115 13231 12121
rect 9950 12084 9956 12096
rect 9232 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 11204 12056 11345 12084
rect 11204 12044 11210 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 11333 12047 11391 12053
rect 1104 11994 13892 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 13892 11994
rect 1104 11920 13892 11942
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 2682 11880 2688 11892
rect 2639 11852 2688 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 3804 11852 4752 11880
rect 3804 11812 3832 11852
rect 2424 11784 3832 11812
rect 2424 11753 2452 11784
rect 3878 11772 3884 11824
rect 3936 11772 3942 11824
rect 4724 11812 4752 11852
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 6730 11880 6736 11892
rect 5132 11852 6132 11880
rect 6691 11852 6736 11880
rect 5132 11840 5138 11852
rect 5813 11815 5871 11821
rect 5813 11812 5825 11815
rect 4724 11784 5304 11812
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 2866 11744 2872 11756
rect 2823 11716 2872 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 1486 11676 1492 11688
rect 1447 11648 1492 11676
rect 1486 11636 1492 11648
rect 1544 11636 1550 11688
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 3145 11679 3203 11685
rect 3145 11676 3157 11679
rect 2556 11648 3157 11676
rect 2556 11636 2562 11648
rect 3145 11645 3157 11648
rect 3191 11645 3203 11679
rect 3145 11639 3203 11645
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3786 11676 3792 11688
rect 3467 11648 3792 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 5276 11676 5304 11784
rect 5368 11784 5825 11812
rect 5368 11753 5396 11784
rect 5813 11781 5825 11784
rect 5859 11781 5871 11815
rect 5813 11775 5871 11781
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 5534 11744 5540 11756
rect 5491 11716 5540 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 5994 11744 6000 11756
rect 5955 11716 6000 11744
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 6104 11753 6132 11852
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 8628 11852 8984 11880
rect 8628 11840 8634 11852
rect 8956 11821 8984 11852
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 9824 11852 10149 11880
rect 9824 11840 9830 11852
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11609 11883 11667 11889
rect 11609 11880 11621 11883
rect 11296 11852 11621 11880
rect 11296 11840 11302 11852
rect 11609 11849 11621 11852
rect 11655 11849 11667 11883
rect 11609 11843 11667 11849
rect 8481 11815 8539 11821
rect 8481 11781 8493 11815
rect 8527 11812 8539 11815
rect 8941 11815 8999 11821
rect 8527 11784 8892 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11744 6147 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 6135 11716 6377 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 6604 11716 6653 11744
rect 6604 11704 6610 11716
rect 6641 11713 6653 11716
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 5721 11679 5779 11685
rect 5276 11648 5672 11676
rect 5644 11608 5672 11648
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 6457 11679 6515 11685
rect 6457 11676 6469 11679
rect 5767 11648 6469 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 6457 11645 6469 11648
rect 6503 11676 6515 11679
rect 6730 11676 6736 11688
rect 6503 11648 6736 11676
rect 6503 11645 6515 11648
rect 6457 11639 6515 11645
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 7116 11676 7144 11707
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 7248 11716 7849 11744
rect 7248 11704 7254 11716
rect 7837 11713 7849 11716
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8754 11744 8760 11756
rect 8619 11716 8760 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 8864 11744 8892 11784
rect 8941 11781 8953 11815
rect 8987 11812 8999 11815
rect 8987 11784 9260 11812
rect 8987 11781 8999 11784
rect 8941 11775 8999 11781
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 8864 11716 9137 11744
rect 9125 11713 9137 11716
rect 9171 11713 9183 11747
rect 9232 11744 9260 11784
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 10042 11812 10048 11824
rect 9364 11784 9409 11812
rect 9876 11784 10048 11812
rect 9364 11772 9370 11784
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 9232 11716 9413 11744
rect 9125 11707 9183 11713
rect 9401 11713 9413 11716
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 7374 11676 7380 11688
rect 7116 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 8018 11676 8024 11688
rect 7975 11648 8024 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 8662 11676 8668 11688
rect 8251 11648 8668 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 8772 11676 8800 11704
rect 9140 11676 9168 11707
rect 9674 11676 9680 11688
rect 8772 11648 8892 11676
rect 9140 11648 9680 11676
rect 8864 11608 8892 11648
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 9876 11685 9904 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 11146 11812 11152 11824
rect 11107 11784 11152 11812
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 12986 11812 12992 11824
rect 12268 11784 12992 11812
rect 10870 11744 10876 11756
rect 10244 11716 10876 11744
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11645 9919 11679
rect 10042 11676 10048 11688
rect 10003 11648 10048 11676
rect 9861 11639 9919 11645
rect 10042 11636 10048 11648
rect 10100 11676 10106 11688
rect 10244 11676 10272 11716
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11054 11744 11060 11756
rect 11015 11716 11060 11744
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 12268 11753 12296 11784
rect 12986 11772 12992 11784
rect 13044 11812 13050 11824
rect 13081 11815 13139 11821
rect 13081 11812 13093 11815
rect 13044 11784 13093 11812
rect 13044 11772 13050 11784
rect 13081 11781 13093 11784
rect 13127 11781 13139 11815
rect 13081 11775 13139 11781
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11296 11716 11713 11744
rect 11296 11704 11302 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 10100 11648 10272 11676
rect 10100 11636 10106 11648
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 10376 11648 10609 11676
rect 10376 11636 10382 11648
rect 10597 11645 10609 11648
rect 10643 11676 10655 11679
rect 11330 11676 11336 11688
rect 10643 11648 11336 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12345 11679 12403 11685
rect 12345 11676 12357 11679
rect 11940 11648 12357 11676
rect 11940 11636 11946 11648
rect 12345 11645 12357 11648
rect 12391 11645 12403 11679
rect 12894 11676 12900 11688
rect 12855 11648 12900 11676
rect 12345 11639 12403 11645
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 9122 11608 9128 11620
rect 5644 11580 8800 11608
rect 8864 11580 9128 11608
rect 2866 11540 2872 11552
rect 2827 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 4893 11543 4951 11549
rect 4893 11509 4905 11543
rect 4939 11540 4951 11543
rect 5074 11540 5080 11552
rect 4939 11512 5080 11540
rect 4939 11509 4951 11512
rect 4893 11503 4951 11509
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5258 11540 5264 11552
rect 5215 11512 5264 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5350 11500 5356 11552
rect 5408 11540 5414 11552
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 5408 11512 5641 11540
rect 5408 11500 5414 11512
rect 5629 11509 5641 11512
rect 5675 11509 5687 11543
rect 5629 11503 5687 11509
rect 6822 11500 6828 11552
rect 6880 11540 6886 11552
rect 7009 11543 7067 11549
rect 7009 11540 7021 11543
rect 6880 11512 7021 11540
rect 6880 11500 6886 11512
rect 7009 11509 7021 11512
rect 7055 11509 7067 11543
rect 8662 11540 8668 11552
rect 8623 11512 8668 11540
rect 7009 11503 7067 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 8772 11540 8800 11580
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 12069 11611 12127 11617
rect 12069 11608 12081 11611
rect 9232 11580 12081 11608
rect 9232 11540 9260 11580
rect 12069 11577 12081 11580
rect 12115 11577 12127 11611
rect 12069 11571 12127 11577
rect 12805 11611 12863 11617
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 12986 11608 12992 11620
rect 12851 11580 12992 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 8772 11512 9260 11540
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 9364 11512 9505 11540
rect 9364 11500 9370 11512
rect 9493 11509 9505 11512
rect 9539 11509 9551 11543
rect 9493 11503 9551 11509
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10284 11512 10517 11540
rect 10284 11500 10290 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 10928 11512 11253 11540
rect 10928 11500 10934 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 13170 11540 13176 11552
rect 13131 11512 13176 11540
rect 11241 11503 11299 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 1104 11450 13892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 13892 11450
rect 1104 11376 13892 11398
rect 3510 11336 3516 11348
rect 3471 11308 3516 11336
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 4614 11336 4620 11348
rect 3615 11308 4620 11336
rect 2590 11228 2596 11280
rect 2648 11268 2654 11280
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 2648 11240 2789 11268
rect 2648 11228 2654 11240
rect 2777 11237 2789 11240
rect 2823 11237 2835 11271
rect 2777 11231 2835 11237
rect 3615 11200 3643 11308
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 5828 11308 6408 11336
rect 3786 11268 3792 11280
rect 3747 11240 3792 11268
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 5828 11277 5856 11308
rect 5445 11271 5503 11277
rect 5445 11268 5457 11271
rect 3936 11240 5457 11268
rect 3936 11228 3942 11240
rect 5445 11237 5457 11240
rect 5491 11237 5503 11271
rect 5445 11231 5503 11237
rect 5813 11271 5871 11277
rect 5813 11237 5825 11271
rect 5859 11237 5871 11271
rect 5813 11231 5871 11237
rect 6273 11271 6331 11277
rect 6273 11237 6285 11271
rect 6319 11237 6331 11271
rect 6380 11268 6408 11308
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 6512 11308 6557 11336
rect 6512 11296 6518 11308
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 7248 11308 7481 11336
rect 7248 11296 7254 11308
rect 7469 11305 7481 11308
rect 7515 11305 7527 11339
rect 7469 11299 7527 11305
rect 6380 11240 6684 11268
rect 6273 11231 6331 11237
rect 2976 11172 3643 11200
rect 2976 11141 3004 11172
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 6288 11200 6316 11231
rect 6656 11212 6684 11240
rect 6914 11228 6920 11280
rect 6972 11268 6978 11280
rect 7009 11271 7067 11277
rect 7009 11268 7021 11271
rect 6972 11240 7021 11268
rect 6972 11228 6978 11240
rect 7009 11237 7021 11240
rect 7055 11268 7067 11271
rect 7055 11240 7972 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 6638 11200 6644 11212
rect 4856 11172 6316 11200
rect 6599 11172 6644 11200
rect 4856 11160 4862 11172
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 7944 11209 7972 11240
rect 11238 11228 11244 11280
rect 11296 11268 11302 11280
rect 11517 11271 11575 11277
rect 11517 11268 11529 11271
rect 11296 11240 11529 11268
rect 11296 11228 11302 11240
rect 11517 11237 11529 11240
rect 11563 11237 11575 11271
rect 11517 11231 11575 11237
rect 12986 11228 12992 11280
rect 13044 11268 13050 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 13044 11240 13185 11268
rect 13044 11228 13050 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 7208 11172 7665 11200
rect 7208 11144 7236 11172
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 7653 11163 7711 11169
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 9306 11200 9312 11212
rect 8720 11172 9076 11200
rect 9267 11172 9312 11200
rect 8720 11160 8726 11172
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 3234 11132 3240 11144
rect 2961 11095 3019 11101
rect 3068 11104 3240 11132
rect 3068 11005 3096 11104
rect 3234 11092 3240 11104
rect 3292 11132 3298 11144
rect 3510 11132 3516 11144
rect 3292 11104 3516 11132
rect 3292 11092 3298 11104
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 3660 11104 3705 11132
rect 3660 11092 3666 11104
rect 3970 11092 3976 11144
rect 4028 11134 4034 11144
rect 4064 11135 4122 11141
rect 4064 11134 4076 11135
rect 4028 11106 4076 11134
rect 4028 11092 4034 11106
rect 4064 11101 4076 11106
rect 4110 11101 4122 11135
rect 4156 11129 4214 11135
rect 4156 11122 4168 11129
rect 4202 11122 4214 11129
rect 4064 11095 4122 11101
rect 3329 11067 3387 11073
rect 3329 11033 3341 11067
rect 3375 11064 3387 11067
rect 3878 11064 3884 11076
rect 3375 11036 3884 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4154 11070 4160 11122
rect 4212 11070 4218 11122
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4525 11135 4583 11141
rect 4304 11104 4349 11132
rect 4433 11129 4491 11135
rect 4525 11129 4537 11135
rect 4304 11092 4310 11104
rect 4433 11095 4445 11129
rect 4479 11101 4537 11129
rect 4571 11101 4583 11135
rect 4706 11132 4712 11144
rect 4667 11104 4712 11132
rect 4479 11095 4491 11101
rect 4525 11095 4583 11101
rect 4433 11089 4491 11095
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 4890 11024 4896 11076
rect 4948 11073 4954 11076
rect 4948 11067 4969 11073
rect 4957 11033 4969 11067
rect 5074 11064 5080 11076
rect 5035 11036 5080 11064
rect 4948 11027 4969 11033
rect 4948 11024 4954 11027
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 5644 11064 5672 11095
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 5776 11104 5821 11132
rect 5776 11092 5782 11104
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 6086 11132 6092 11144
rect 5960 11104 6005 11132
rect 6047 11104 6092 11132
rect 5960 11092 5966 11104
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11101 6515 11135
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6457 11095 6515 11101
rect 6472 11064 6500 11095
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6880 11104 6929 11132
rect 6880 11092 6886 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 7190 11132 7196 11144
rect 7103 11104 7196 11132
rect 6917 11095 6975 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 6840 11064 6868 11092
rect 5644 11036 6868 11064
rect 7098 11024 7104 11076
rect 7156 11064 7162 11076
rect 7300 11064 7328 11095
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7432 11104 8033 11132
rect 7432 11092 7438 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8938 11132 8944 11144
rect 8899 11104 8944 11132
rect 8021 11095 8079 11101
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 9048 11132 9076 11172
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 9106 11135 9164 11141
rect 9106 11132 9118 11135
rect 9048 11104 9118 11132
rect 9106 11101 9118 11104
rect 9152 11101 9164 11135
rect 9106 11095 9164 11101
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9272 11104 9317 11132
rect 9272 11092 9278 11104
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9493 11135 9551 11141
rect 9493 11132 9505 11135
rect 9456 11104 9505 11132
rect 9456 11092 9462 11104
rect 9493 11101 9505 11104
rect 9539 11101 9551 11135
rect 9766 11132 9772 11144
rect 9727 11104 9772 11132
rect 9493 11095 9551 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10226 11132 10232 11144
rect 10187 11104 10232 11132
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 13170 11132 13176 11144
rect 13131 11104 13176 11132
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 7156 11036 7328 11064
rect 7156 11024 7162 11036
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 9953 11067 10011 11073
rect 9953 11064 9965 11067
rect 9364 11036 9965 11064
rect 9364 11024 9370 11036
rect 9953 11033 9965 11036
rect 9999 11033 10011 11067
rect 10134 11064 10140 11076
rect 10095 11036 10140 11064
rect 9953 11027 10011 11033
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 3053 10999 3111 11005
rect 3053 10965 3065 10999
rect 3099 10965 3111 10999
rect 3053 10959 3111 10965
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 3970 10996 3976 11008
rect 3200 10968 3976 10996
rect 3200 10956 3206 10968
rect 3970 10956 3976 10968
rect 4028 10996 4034 11008
rect 4154 10996 4160 11008
rect 4028 10968 4160 10996
rect 4028 10956 4034 10968
rect 4154 10956 4160 10968
rect 4212 10956 4218 11008
rect 4801 10999 4859 11005
rect 4801 10965 4813 10999
rect 4847 10996 4859 10999
rect 5534 10996 5540 11008
rect 4847 10968 5540 10996
rect 4847 10965 4859 10968
rect 4801 10959 4859 10965
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 6454 10996 6460 11008
rect 5776 10968 6460 10996
rect 5776 10956 5782 10968
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8665 10999 8723 11005
rect 8665 10996 8677 10999
rect 8168 10968 8677 10996
rect 8168 10956 8174 10968
rect 8665 10965 8677 10968
rect 8711 10996 8723 10999
rect 9398 10996 9404 11008
rect 8711 10968 9404 10996
rect 8711 10965 8723 10968
rect 8665 10959 8723 10965
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 9582 10996 9588 11008
rect 9543 10968 9588 10996
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 1104 10906 13892 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 13892 10906
rect 1104 10832 13892 10854
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 4890 10792 4896 10804
rect 3191 10764 4896 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 8389 10795 8447 10801
rect 8389 10761 8401 10795
rect 8435 10792 8447 10795
rect 9214 10792 9220 10804
rect 8435 10764 9220 10792
rect 8435 10761 8447 10764
rect 8389 10755 8447 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 9456 10764 9597 10792
rect 9456 10752 9462 10764
rect 9585 10761 9597 10764
rect 9631 10792 9643 10795
rect 9674 10792 9680 10804
rect 9631 10764 9680 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 9953 10795 10011 10801
rect 9953 10792 9965 10795
rect 9916 10764 9965 10792
rect 9916 10752 9922 10764
rect 9953 10761 9965 10764
rect 9999 10761 10011 10795
rect 9953 10755 10011 10761
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10134 10792 10140 10804
rect 10091 10764 10140 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 2314 10684 2320 10736
rect 2372 10684 2378 10736
rect 3602 10684 3608 10736
rect 3660 10724 3666 10736
rect 4798 10724 4804 10736
rect 3660 10696 4804 10724
rect 3660 10684 3666 10696
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 3712 10665 3740 10696
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 5626 10724 5632 10736
rect 4999 10696 5632 10724
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3697 10619 3755 10625
rect 3804 10628 4077 10656
rect 3804 10600 3832 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4999 10665 5027 10696
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 6086 10684 6092 10736
rect 6144 10724 6150 10736
rect 6457 10727 6515 10733
rect 6457 10724 6469 10727
rect 6144 10696 6469 10724
rect 6144 10684 6150 10696
rect 6457 10693 6469 10696
rect 6503 10693 6515 10727
rect 6457 10687 6515 10693
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 7190 10724 7196 10736
rect 6604 10696 6776 10724
rect 7151 10696 7196 10724
rect 6604 10684 6610 10696
rect 4984 10659 5042 10665
rect 4212 10628 4257 10656
rect 4212 10616 4218 10628
rect 4984 10625 4996 10659
rect 5030 10625 5042 10659
rect 4984 10619 5042 10625
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5445 10659 5503 10665
rect 5316 10628 5361 10656
rect 5316 10616 5322 10628
rect 5445 10625 5457 10659
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10557 3663 10591
rect 3786 10588 3792 10600
rect 3747 10560 3792 10588
rect 3605 10551 3663 10557
rect 3620 10520 3648 10551
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 4525 10591 4583 10597
rect 3936 10560 3981 10588
rect 3936 10548 3942 10560
rect 4525 10557 4537 10591
rect 4571 10557 4583 10591
rect 4525 10551 4583 10557
rect 4540 10520 4568 10551
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5460 10588 5488 10619
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5592 10628 5733 10656
rect 5592 10616 5598 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10656 6423 10659
rect 6638 10656 6644 10668
rect 6411 10628 6644 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 6638 10616 6644 10628
rect 6696 10616 6702 10668
rect 6748 10665 6776 10696
rect 7190 10684 7196 10696
rect 7248 10724 7254 10736
rect 9416 10724 9444 10752
rect 7248 10696 7512 10724
rect 7248 10684 7254 10696
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7282 10656 7288 10668
rect 6779 10628 7288 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7484 10665 7512 10696
rect 7944 10696 8984 10724
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 6822 10588 6828 10600
rect 4672 10560 5488 10588
rect 6783 10560 6828 10588
rect 4672 10548 4678 10560
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7098 10588 7104 10600
rect 7059 10560 7104 10588
rect 7098 10548 7104 10560
rect 7156 10588 7162 10600
rect 7944 10597 7972 10696
rect 8956 10668 8984 10696
rect 9121 10696 9444 10724
rect 9968 10724 9996 10755
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10413 10795 10471 10801
rect 10413 10761 10425 10795
rect 10459 10792 10471 10795
rect 11882 10792 11888 10804
rect 10459 10764 11888 10792
rect 10459 10761 10471 10764
rect 10413 10755 10471 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12345 10795 12403 10801
rect 12345 10761 12357 10795
rect 12391 10792 12403 10795
rect 12894 10792 12900 10804
rect 12391 10764 12900 10792
rect 12391 10761 12403 10764
rect 12345 10755 12403 10761
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 11238 10724 11244 10736
rect 9968 10696 10916 10724
rect 11199 10696 11244 10724
rect 8110 10656 8116 10668
rect 8071 10628 8116 10656
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 8570 10656 8576 10668
rect 8531 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8662 10616 8668 10668
rect 8720 10662 8779 10668
rect 8720 10628 8733 10662
rect 8767 10628 8779 10662
rect 8938 10656 8944 10668
rect 8851 10628 8944 10656
rect 8720 10622 8779 10628
rect 8720 10616 8726 10622
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9121 10665 9149 10696
rect 9098 10659 9156 10665
rect 9098 10625 9110 10659
rect 9144 10625 9156 10659
rect 9098 10619 9156 10625
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10284 10628 10793 10656
rect 10284 10616 10290 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 10888 10656 10916 10696
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 12069 10727 12127 10733
rect 12069 10724 12081 10727
rect 11348 10696 12081 10724
rect 11348 10656 11376 10696
rect 12069 10693 12081 10696
rect 12115 10693 12127 10727
rect 12069 10687 12127 10693
rect 12437 10727 12495 10733
rect 12437 10693 12449 10727
rect 12483 10724 12495 10727
rect 13078 10724 13084 10736
rect 12483 10696 13084 10724
rect 12483 10693 12495 10696
rect 12437 10687 12495 10693
rect 13078 10684 13084 10696
rect 13136 10724 13142 10736
rect 13173 10727 13231 10733
rect 13173 10724 13185 10727
rect 13136 10696 13185 10724
rect 13136 10684 13142 10696
rect 13173 10693 13185 10696
rect 13219 10693 13231 10727
rect 13173 10687 13231 10693
rect 13262 10684 13268 10736
rect 13320 10724 13326 10736
rect 13449 10727 13507 10733
rect 13449 10724 13461 10727
rect 13320 10696 13461 10724
rect 13320 10684 13326 10696
rect 13449 10693 13461 10696
rect 13495 10693 13507 10727
rect 13449 10687 13507 10693
rect 11514 10656 11520 10668
rect 10888 10628 11376 10656
rect 11475 10628 11520 10656
rect 10781 10619 10839 10625
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11790 10656 11796 10668
rect 11751 10628 11796 10656
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12618 10656 12624 10668
rect 12575 10628 12624 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 7581 10591 7639 10597
rect 7581 10588 7593 10591
rect 7156 10560 7593 10588
rect 7156 10548 7162 10560
rect 7581 10557 7593 10560
rect 7627 10557 7639 10591
rect 7581 10551 7639 10557
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10557 8539 10591
rect 8846 10588 8852 10600
rect 8807 10560 8852 10588
rect 8481 10551 8539 10557
rect 5258 10520 5264 10532
rect 3620 10492 4292 10520
rect 4540 10492 5264 10520
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4264 10461 4292 10492
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 7745 10523 7803 10529
rect 7745 10489 7757 10523
rect 7791 10520 7803 10523
rect 7944 10520 7972 10551
rect 7791 10492 7972 10520
rect 8496 10520 8524 10551
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 9950 10588 9956 10600
rect 9907 10560 9956 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10588 11391 10591
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11379 10560 11897 10588
rect 11379 10557 11391 10560
rect 11333 10551 11391 10557
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 9309 10523 9367 10529
rect 9309 10520 9321 10523
rect 8496 10492 9321 10520
rect 7791 10489 7803 10492
rect 7745 10483 7803 10489
rect 9309 10489 9321 10492
rect 9355 10520 9367 10523
rect 9398 10520 9404 10532
rect 9355 10492 9404 10520
rect 9355 10489 9367 10492
rect 9309 10483 9367 10489
rect 9398 10480 9404 10492
rect 9456 10480 9462 10532
rect 9646 10492 10456 10520
rect 4249 10455 4307 10461
rect 4249 10421 4261 10455
rect 4295 10452 4307 10455
rect 4706 10452 4712 10464
rect 4295 10424 4712 10452
rect 4295 10421 4307 10424
rect 4249 10415 4307 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5074 10452 5080 10464
rect 5035 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5718 10452 5724 10464
rect 5408 10424 5724 10452
rect 5408 10412 5414 10424
rect 5718 10412 5724 10424
rect 5776 10452 5782 10464
rect 5813 10455 5871 10461
rect 5813 10452 5825 10455
rect 5776 10424 5825 10452
rect 5776 10412 5782 10424
rect 5813 10421 5825 10424
rect 5859 10421 5871 10455
rect 5813 10415 5871 10421
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 9646 10452 9674 10492
rect 10428 10464 10456 10492
rect 8720 10424 9674 10452
rect 8720 10412 8726 10424
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10468 10424 10517 10452
rect 10468 10412 10474 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 11698 10452 11704 10464
rect 11659 10424 11704 10452
rect 10505 10415 10563 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 1104 10362 13892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 13892 10362
rect 1104 10288 13892 10310
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 1949 10251 2007 10257
rect 1949 10248 1961 10251
rect 1728 10220 1961 10248
rect 1728 10208 1734 10220
rect 1949 10217 1961 10220
rect 1995 10217 2007 10251
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 1949 10211 2007 10217
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2501 10251 2559 10257
rect 2501 10217 2513 10251
rect 2547 10248 2559 10251
rect 2866 10248 2872 10260
rect 2547 10220 2872 10248
rect 2547 10217 2559 10220
rect 2501 10211 2559 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 4614 10248 4620 10260
rect 4571 10220 4620 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 5350 10248 5356 10260
rect 5000 10220 5356 10248
rect 4338 10180 4344 10192
rect 3528 10152 4344 10180
rect 3418 10112 3424 10124
rect 2056 10084 3424 10112
rect 2056 10053 2084 10084
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10044 2191 10047
rect 2866 10044 2872 10056
rect 2179 10016 2872 10044
rect 2179 10013 2191 10016
rect 2133 10007 2191 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3234 10044 3240 10056
rect 3195 10016 3240 10044
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3528 10053 3556 10152
rect 4338 10140 4344 10152
rect 4396 10180 4402 10192
rect 5000 10180 5028 10220
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 6914 10248 6920 10260
rect 5500 10220 6776 10248
rect 6875 10220 6920 10248
rect 5500 10208 5506 10220
rect 6362 10180 6368 10192
rect 4396 10152 5028 10180
rect 6323 10152 6368 10180
rect 4396 10140 4402 10152
rect 6362 10140 6368 10152
rect 6420 10140 6426 10192
rect 6748 10180 6776 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 8021 10251 8079 10257
rect 8021 10248 8033 10251
rect 7156 10220 8033 10248
rect 7156 10208 7162 10220
rect 8021 10217 8033 10220
rect 8067 10217 8079 10251
rect 8021 10211 8079 10217
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 8168 10220 8309 10248
rect 8168 10208 8174 10220
rect 8297 10217 8309 10220
rect 8343 10217 8355 10251
rect 8297 10211 8355 10217
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8628 10220 8677 10248
rect 8628 10208 8634 10220
rect 8665 10217 8677 10220
rect 8711 10217 8723 10251
rect 10042 10248 10048 10260
rect 8665 10211 8723 10217
rect 8864 10220 10048 10248
rect 8864 10180 8892 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10505 10251 10563 10257
rect 10505 10248 10517 10251
rect 10244 10220 10517 10248
rect 6748 10152 8892 10180
rect 8938 10140 8944 10192
rect 8996 10140 9002 10192
rect 9950 10140 9956 10192
rect 10008 10180 10014 10192
rect 10244 10180 10272 10220
rect 10505 10217 10517 10220
rect 10551 10248 10563 10251
rect 10870 10248 10876 10260
rect 10551 10220 10876 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 10410 10180 10416 10192
rect 10008 10152 10272 10180
rect 10371 10152 10416 10180
rect 10008 10140 10014 10152
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 11790 10180 11796 10192
rect 11440 10152 11796 10180
rect 4249 10115 4307 10121
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 4614 10112 4620 10124
rect 4295 10084 4620 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 4614 10072 4620 10084
rect 4672 10112 4678 10124
rect 4672 10084 4936 10112
rect 4672 10072 4678 10084
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10013 3571 10047
rect 3513 10007 3571 10013
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10044 3663 10047
rect 3694 10044 3700 10056
rect 3651 10016 3700 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 2222 9936 2228 9988
rect 2280 9976 2286 9988
rect 2958 9976 2964 9988
rect 2280 9948 2964 9976
rect 2280 9936 2286 9948
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 3142 9936 3148 9988
rect 3200 9976 3206 9988
rect 3344 9976 3372 10007
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4157 10007 4215 10013
rect 3786 9976 3792 9988
rect 3200 9948 3792 9976
rect 3200 9936 3206 9948
rect 3786 9936 3792 9948
rect 3844 9976 3850 9988
rect 4172 9976 4200 10007
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4908 10053 4936 10084
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 5684 10084 5758 10112
rect 5684 10072 5690 10084
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 4893 10007 4951 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5442 10044 5448 10056
rect 5403 10016 5448 10044
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5730 10053 5758 10084
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 7190 10112 7196 10124
rect 6052 10084 6224 10112
rect 7151 10084 7196 10112
rect 6052 10072 6058 10084
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 6196 10053 6224 10084
rect 7190 10072 7196 10084
rect 7248 10112 7254 10124
rect 7653 10115 7711 10121
rect 7248 10084 7420 10112
rect 7248 10072 7254 10084
rect 6186 10047 6244 10053
rect 5868 10016 5913 10044
rect 5868 10004 5874 10016
rect 6186 10013 6198 10047
rect 6232 10013 6244 10047
rect 6186 10007 6244 10013
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 6914 10044 6920 10056
rect 6871 10016 6920 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 3844 9948 4200 9976
rect 3844 9936 3850 9948
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 5997 9979 6055 9985
rect 5684 9948 5729 9976
rect 5684 9936 5690 9948
rect 5997 9945 6009 9979
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6089 9979 6147 9985
rect 6089 9945 6101 9979
rect 6135 9976 6147 9979
rect 6840 9976 6868 10007
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7282 10044 7288 10056
rect 7243 10016 7288 10044
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7392 10044 7420 10084
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 8570 10112 8576 10124
rect 7699 10084 8576 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 8956 10112 8984 10140
rect 8772 10084 8984 10112
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7392 10016 7757 10044
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8772 10053 8800 10084
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 8168 10016 8493 10044
rect 8168 10004 8174 10016
rect 8481 10013 8493 10016
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10013 8815 10047
rect 8938 10044 8944 10056
rect 8899 10016 8944 10044
rect 8757 10007 8815 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9398 10044 9404 10056
rect 9359 10016 9404 10044
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9508 10016 9689 10044
rect 6135 9948 6868 9976
rect 7300 9976 7328 10004
rect 7929 9979 7987 9985
rect 7929 9976 7941 9979
rect 7300 9948 7941 9976
rect 6135 9945 6147 9948
rect 6089 9939 6147 9945
rect 7929 9945 7941 9948
rect 7975 9945 7987 9979
rect 7929 9939 7987 9945
rect 3050 9908 3056 9920
rect 3011 9880 3056 9908
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 6012 9908 6040 9939
rect 8662 9936 8668 9988
rect 8720 9976 8726 9988
rect 9033 9979 9091 9985
rect 9033 9976 9045 9979
rect 8720 9948 9045 9976
rect 8720 9936 8726 9948
rect 9033 9945 9045 9948
rect 9079 9945 9091 9979
rect 9033 9939 9091 9945
rect 6270 9908 6276 9920
rect 6012 9880 6276 9908
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 6641 9911 6699 9917
rect 6641 9877 6653 9911
rect 6687 9908 6699 9911
rect 6822 9908 6828 9920
rect 6687 9880 6828 9908
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 9508 9908 9536 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10044 10011 10047
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9999 10016 10149 10044
rect 9999 10013 10011 10016
rect 9953 10007 10011 10013
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10044 10287 10047
rect 10428 10044 10456 10140
rect 10275 10016 10456 10044
rect 10689 10047 10747 10053
rect 10275 10013 10287 10016
rect 10229 10007 10287 10013
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 11146 10044 11152 10056
rect 10735 10016 11152 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 11440 10053 11468 10152
rect 11790 10140 11796 10152
rect 11848 10140 11854 10192
rect 13078 10180 13084 10192
rect 13039 10152 13084 10180
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 11698 10112 11704 10124
rect 11659 10084 11704 10112
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12618 10044 12624 10056
rect 12579 10016 12624 10044
rect 12253 10007 12311 10013
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 11514 9976 11520 9988
rect 11112 9948 11520 9976
rect 11112 9936 11118 9948
rect 11514 9936 11520 9948
rect 11572 9976 11578 9988
rect 11609 9979 11667 9985
rect 11609 9976 11621 9979
rect 11572 9948 11621 9976
rect 11572 9936 11578 9948
rect 11609 9945 11621 9948
rect 11655 9945 11667 9979
rect 11609 9939 11667 9945
rect 8628 9880 9536 9908
rect 8628 9868 8634 9880
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 12268 9908 12296 10007
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 13320 10016 13461 10044
rect 13320 10004 13326 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13173 9979 13231 9985
rect 13173 9945 13185 9979
rect 13219 9945 13231 9979
rect 13173 9939 13231 9945
rect 11204 9880 12296 9908
rect 13188 9908 13216 9939
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 13188 9880 13277 9908
rect 11204 9868 11210 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 13265 9871 13323 9877
rect 14093 9911 14151 9917
rect 14093 9877 14105 9911
rect 14139 9908 14151 9911
rect 14182 9908 14188 9920
rect 14139 9880 14188 9908
rect 14139 9877 14151 9880
rect 14093 9871 14151 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 1104 9818 13892 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 13892 9818
rect 1104 9744 13892 9766
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 6546 9704 6552 9716
rect 3016 9676 6552 9704
rect 3016 9664 3022 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 8113 9707 8171 9713
rect 8113 9704 8125 9707
rect 6972 9676 8125 9704
rect 6972 9664 6978 9676
rect 8113 9673 8125 9676
rect 8159 9673 8171 9707
rect 8846 9704 8852 9716
rect 8807 9676 8852 9704
rect 8113 9667 8171 9673
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 2222 9596 2228 9648
rect 2280 9596 2286 9648
rect 3786 9636 3792 9648
rect 3747 9608 3792 9636
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 5534 9636 5540 9648
rect 3988 9608 4752 9636
rect 3602 9577 3608 9580
rect 3600 9568 3608 9577
rect 3563 9540 3608 9568
rect 3600 9531 3608 9540
rect 3602 9528 3608 9531
rect 3660 9528 3666 9580
rect 3988 9577 4016 9608
rect 4724 9580 4752 9608
rect 4908 9608 5540 9636
rect 4908 9580 4936 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 5868 9608 6040 9636
rect 5868 9596 5874 9608
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3697 9531 3755 9537
rect 3804 9540 3985 9568
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 3145 9503 3203 9509
rect 1719 9472 2774 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2746 9432 2774 9472
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3326 9500 3332 9512
rect 3191 9472 3332 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 3326 9460 3332 9472
rect 3384 9500 3390 9512
rect 3712 9500 3740 9531
rect 3804 9512 3832 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4440 9571 4498 9577
rect 4440 9537 4452 9571
rect 4486 9537 4498 9571
rect 4706 9568 4712 9580
rect 4619 9540 4712 9568
rect 4440 9531 4498 9537
rect 3384 9472 3740 9500
rect 3384 9460 3390 9472
rect 3786 9460 3792 9512
rect 3844 9460 3850 9512
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 3936 9472 4077 9500
rect 3936 9460 3942 9472
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 4338 9500 4344 9512
rect 4299 9472 4344 9500
rect 4065 9463 4123 9469
rect 4338 9460 4344 9472
rect 4396 9460 4402 9512
rect 4448 9500 4476 9531
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 4890 9568 4896 9580
rect 4851 9540 4896 9568
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5129 9571 5187 9577
rect 5040 9540 5085 9568
rect 5040 9528 5046 9540
rect 5129 9537 5141 9571
rect 5175 9568 5187 9571
rect 5902 9568 5908 9580
rect 5175 9540 5908 9568
rect 5175 9537 5212 9540
rect 5129 9531 5212 9537
rect 4798 9500 4804 9512
rect 4448 9472 4804 9500
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 3421 9435 3479 9441
rect 3421 9432 3433 9435
rect 2746 9404 3433 9432
rect 3421 9401 3433 9404
rect 3467 9401 3479 9435
rect 3421 9395 3479 9401
rect 3602 9392 3608 9444
rect 3660 9432 3666 9444
rect 5184 9432 5212 9531
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 6012 9577 6040 9608
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6420 9608 6653 9636
rect 6420 9596 6426 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 6641 9599 6699 9605
rect 8665 9639 8723 9645
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 8938 9636 8944 9648
rect 8711 9608 8944 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 10318 9596 10324 9648
rect 10376 9636 10382 9648
rect 10689 9639 10747 9645
rect 10689 9636 10701 9639
rect 10376 9608 10701 9636
rect 10376 9596 10382 9608
rect 10689 9605 10701 9608
rect 10735 9636 10747 9639
rect 10873 9639 10931 9645
rect 10873 9636 10885 9639
rect 10735 9608 10885 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 10873 9605 10885 9608
rect 10919 9605 10931 9639
rect 11054 9636 11060 9648
rect 11015 9608 11060 9636
rect 10873 9599 10931 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 12897 9639 12955 9645
rect 12897 9605 12909 9639
rect 12943 9636 12955 9639
rect 12986 9636 12992 9648
rect 12943 9608 12992 9636
rect 12943 9605 12955 9608
rect 12897 9599 12955 9605
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 8294 9568 8300 9580
rect 5997 9531 6055 9537
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 5592 9472 6377 9500
rect 5592 9460 5598 9472
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 7760 9500 7788 9554
rect 8255 9540 8300 9568
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 6365 9463 6423 9469
rect 6472 9472 7788 9500
rect 8496 9500 8524 9531
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8628 9540 8769 9568
rect 8628 9528 8634 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9568 9183 9571
rect 9674 9568 9680 9580
rect 9171 9540 9680 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 10134 9568 10140 9580
rect 10095 9540 10140 9568
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11296 9540 11529 9568
rect 11296 9528 11302 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 12124 9540 12173 9568
rect 12124 9528 12130 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9568 12495 9571
rect 13265 9571 13323 9577
rect 12483 9540 12756 9568
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 12728 9512 12756 9540
rect 13265 9537 13277 9571
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 8846 9500 8852 9512
rect 8496 9472 8852 9500
rect 3660 9404 5212 9432
rect 3660 9392 3666 9404
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 6181 9435 6239 9441
rect 5500 9404 5948 9432
rect 5500 9392 5506 9404
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3620 9364 3648 9392
rect 2832 9336 3648 9364
rect 2832 9324 2838 9336
rect 5166 9324 5172 9376
rect 5224 9364 5230 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 5224 9336 5273 9364
rect 5224 9324 5230 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5261 9327 5319 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 5920 9364 5948 9404
rect 6181 9401 6193 9435
rect 6227 9432 6239 9435
rect 6472 9432 6500 9472
rect 6227 9404 6500 9432
rect 6227 9401 6239 9404
rect 6181 9395 6239 9401
rect 6822 9364 6828 9376
rect 5920 9336 6828 9364
rect 6822 9324 6828 9336
rect 6880 9364 6886 9376
rect 8496 9364 8524 9472
rect 8846 9460 8852 9472
rect 8904 9500 8910 9512
rect 10502 9500 10508 9512
rect 8904 9472 10508 9500
rect 8904 9460 8910 9472
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 12710 9500 12716 9512
rect 12623 9472 12716 9500
rect 12710 9460 12716 9472
rect 12768 9500 12774 9512
rect 13280 9500 13308 9531
rect 12768 9472 13308 9500
rect 12768 9460 12774 9472
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 11974 9432 11980 9444
rect 10928 9404 11980 9432
rect 10928 9392 10934 9404
rect 11974 9392 11980 9404
rect 12032 9432 12038 9444
rect 12529 9435 12587 9441
rect 12529 9432 12541 9435
rect 12032 9404 12541 9432
rect 12032 9392 12038 9404
rect 12529 9401 12541 9404
rect 12575 9432 12587 9435
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 12575 9404 13461 9432
rect 12575 9401 12587 9404
rect 12529 9395 12587 9401
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 13078 9364 13084 9376
rect 6880 9336 8524 9364
rect 13039 9336 13084 9364
rect 6880 9324 6886 9336
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 1104 9274 13892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 13892 9274
rect 1104 9200 13892 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 4614 9160 4620 9172
rect 3559 9132 4620 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 6641 9163 6699 9169
rect 6641 9160 6653 9163
rect 5040 9132 6653 9160
rect 5040 9120 5046 9132
rect 6641 9129 6653 9132
rect 6687 9129 6699 9163
rect 6641 9123 6699 9129
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7190 9160 7196 9172
rect 6963 9132 7196 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 2409 9095 2467 9101
rect 2409 9092 2421 9095
rect 1995 9064 2421 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 2409 9061 2421 9064
rect 2455 9092 2467 9095
rect 2866 9092 2872 9104
rect 2455 9064 2872 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 2866 9052 2872 9064
rect 2924 9092 2930 9104
rect 3418 9092 3424 9104
rect 2924 9064 3424 9092
rect 2924 9052 2930 9064
rect 3418 9052 3424 9064
rect 3476 9092 3482 9104
rect 4065 9095 4123 9101
rect 4065 9092 4077 9095
rect 3476 9064 4077 9092
rect 3476 9052 3482 9064
rect 1854 8916 1860 8968
rect 1912 8956 1918 8968
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1912 8928 1961 8956
rect 1912 8916 1918 8928
rect 1949 8925 1961 8928
rect 1995 8956 2007 8959
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1995 8928 2053 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 3804 8965 3832 9064
rect 4065 9061 4077 9064
rect 4111 9061 4123 9095
rect 4065 9055 4123 9061
rect 5166 9024 5172 9036
rect 5127 8996 5172 9024
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 3384 8928 3433 8956
rect 3384 8916 3390 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 6656 8956 6684 9123
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 8846 9160 8852 9172
rect 8803 9132 8852 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9030 9024 9036 9036
rect 8991 8996 9036 9024
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 9692 9024 9720 9120
rect 10318 9092 10324 9104
rect 10279 9064 10324 9092
rect 10318 9052 10324 9064
rect 10376 9052 10382 9104
rect 12526 9052 12532 9104
rect 12584 9092 12590 9104
rect 12805 9095 12863 9101
rect 12805 9092 12817 9095
rect 12584 9064 12817 9092
rect 12584 9052 12590 9064
rect 12805 9061 12817 9064
rect 12851 9061 12863 9095
rect 12805 9055 12863 9061
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 9692 8996 9873 9024
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 13078 9024 13084 9036
rect 11471 8996 13084 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6656 8928 6837 8956
rect 4893 8919 4951 8925
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 4908 8888 4936 8919
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7064 8928 7481 8956
rect 7064 8916 7070 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8956 10931 8959
rect 11238 8956 11244 8968
rect 10919 8928 11244 8956
rect 10919 8925 10931 8928
rect 10873 8919 10931 8925
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11514 8956 11520 8968
rect 11475 8928 11520 8956
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12710 8956 12716 8968
rect 12671 8928 12716 8956
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13320 8928 13461 8956
rect 13320 8916 13326 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 5442 8888 5448 8900
rect 4908 8860 5448 8888
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 6178 8848 6184 8900
rect 6236 8848 6242 8900
rect 7926 8888 7932 8900
rect 7887 8860 7932 8888
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 10413 8891 10471 8897
rect 8076 8860 8121 8888
rect 8076 8848 8082 8860
rect 10413 8857 10425 8891
rect 10459 8888 10471 8891
rect 10597 8891 10655 8897
rect 10597 8888 10609 8891
rect 10459 8860 10609 8888
rect 10459 8857 10471 8860
rect 10413 8851 10471 8857
rect 10597 8857 10609 8860
rect 10643 8857 10655 8891
rect 10597 8851 10655 8857
rect 11333 8891 11391 8897
rect 11333 8857 11345 8891
rect 11379 8888 11391 8891
rect 12066 8888 12072 8900
rect 11379 8860 12072 8888
rect 11379 8857 11391 8860
rect 11333 8851 11391 8857
rect 12066 8848 12072 8860
rect 12124 8888 12130 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12124 8860 13185 8888
rect 12124 8848 12130 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 3786 8820 3792 8832
rect 3384 8792 3792 8820
rect 3384 8780 3390 8792
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 3973 8823 4031 8829
rect 3973 8820 3985 8823
rect 3936 8792 3985 8820
rect 3936 8780 3942 8792
rect 3973 8789 3985 8792
rect 4019 8789 4031 8823
rect 3973 8783 4031 8789
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 4212 8792 8493 8820
rect 4212 8780 4218 8792
rect 8481 8789 8493 8792
rect 8527 8820 8539 8823
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 8527 8792 9229 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 9309 8823 9367 8829
rect 9309 8789 9321 8823
rect 9355 8820 9367 8823
rect 9398 8820 9404 8832
rect 9355 8792 9404 8820
rect 9355 8789 9367 8792
rect 9309 8783 9367 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 10502 8820 10508 8832
rect 10463 8792 10508 8820
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 13078 8780 13084 8832
rect 13136 8820 13142 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 13136 8792 13277 8820
rect 13136 8780 13142 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 1104 8730 13892 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 13892 8730
rect 1104 8656 13892 8678
rect 3326 8616 3332 8628
rect 2148 8588 3332 8616
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 1854 8480 1860 8492
rect 1811 8452 1860 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2148 8489 2176 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 4617 8619 4675 8625
rect 3476 8588 4568 8616
rect 3476 8576 3482 8588
rect 2317 8551 2375 8557
rect 2317 8517 2329 8551
rect 2363 8548 2375 8551
rect 2866 8548 2872 8560
rect 2363 8520 2872 8548
rect 2363 8517 2375 8520
rect 2317 8511 2375 8517
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 3050 8508 3056 8560
rect 3108 8548 3114 8560
rect 3145 8551 3203 8557
rect 3145 8548 3157 8551
rect 3108 8520 3157 8548
rect 3108 8508 3114 8520
rect 3145 8517 3157 8520
rect 3191 8517 3203 8551
rect 3145 8511 3203 8517
rect 3878 8508 3884 8560
rect 3936 8508 3942 8560
rect 4540 8548 4568 8588
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 4890 8616 4896 8628
rect 4663 8588 4896 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5902 8616 5908 8628
rect 5767 8588 5908 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6178 8616 6184 8628
rect 6135 8588 6184 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8849 8619 8907 8625
rect 7984 8588 8616 8616
rect 7984 8576 7990 8588
rect 5810 8548 5816 8560
rect 4540 8520 5816 8548
rect 5810 8508 5816 8520
rect 5868 8548 5874 8560
rect 8588 8557 8616 8588
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 10134 8616 10140 8628
rect 8895 8588 10140 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 10134 8576 10140 8588
rect 10192 8616 10198 8628
rect 11514 8616 11520 8628
rect 10192 8588 10824 8616
rect 11475 8588 11520 8616
rect 10192 8576 10198 8588
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5868 8520 6377 8548
rect 5868 8508 5874 8520
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2406 8480 2412 8492
rect 2367 8452 2412 8480
rect 2133 8443 2191 8449
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 2553 8483 2611 8489
rect 2553 8449 2565 8483
rect 2599 8480 2611 8483
rect 2774 8480 2780 8492
rect 2599 8452 2780 8480
rect 2599 8449 2611 8452
rect 2553 8443 2611 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 5920 8489 5948 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 8573 8551 8631 8557
rect 8573 8517 8585 8551
rect 8619 8548 8631 8551
rect 8757 8551 8815 8557
rect 8757 8548 8769 8551
rect 8619 8520 8769 8548
rect 8619 8517 8631 8520
rect 8573 8511 8631 8517
rect 8757 8517 8769 8520
rect 8803 8517 8815 8551
rect 9030 8548 9036 8560
rect 8991 8520 9036 8548
rect 8757 8511 8815 8517
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 9677 8551 9735 8557
rect 9677 8517 9689 8551
rect 9723 8548 9735 8551
rect 10502 8548 10508 8560
rect 9723 8520 10508 8548
rect 9723 8517 9735 8520
rect 9677 8511 9735 8517
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10796 8557 10824 8588
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 12676 8588 12817 8616
rect 12676 8576 12682 8588
rect 12805 8585 12817 8588
rect 12851 8585 12863 8619
rect 12805 8579 12863 8585
rect 10781 8551 10839 8557
rect 10781 8517 10793 8551
rect 10827 8517 10839 8551
rect 10781 8511 10839 8517
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8548 11391 8551
rect 11422 8548 11428 8560
rect 11379 8520 11428 8548
rect 11379 8517 11391 8520
rect 11333 8511 11391 8517
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 4764 8452 5641 8480
rect 4764 8440 4770 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 7006 8480 7012 8492
rect 6967 8452 7012 8480
rect 5905 8443 5963 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 8110 8480 8116 8492
rect 8071 8452 8116 8480
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9263 8452 9873 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9861 8449 9873 8452
rect 9907 8480 9919 8483
rect 10410 8480 10416 8492
rect 9907 8452 10416 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10796 8480 10824 8511
rect 11422 8508 11428 8520
rect 11480 8548 11486 8560
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 11480 8520 11989 8548
rect 11480 8508 11486 8520
rect 11977 8517 11989 8520
rect 12023 8517 12035 8551
rect 12526 8548 12532 8560
rect 12487 8520 12532 8548
rect 11977 8511 12035 8517
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10796 8452 11069 8480
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11057 8443 11115 8449
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 13096 8452 13185 8480
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 9769 8415 9827 8421
rect 2915 8384 3004 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 1946 8304 1952 8356
rect 2004 8344 2010 8356
rect 2041 8347 2099 8353
rect 2041 8344 2053 8347
rect 2004 8316 2053 8344
rect 2004 8304 2010 8316
rect 2041 8313 2053 8316
rect 2087 8313 2099 8347
rect 2041 8307 2099 8313
rect 2976 8288 3004 8384
rect 9769 8381 9781 8415
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 9784 8344 9812 8375
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 12032 8384 12081 8412
rect 12032 8372 12038 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 9784 8316 10885 8344
rect 10873 8313 10885 8316
rect 10919 8313 10931 8347
rect 10873 8307 10931 8313
rect 12713 8347 12771 8353
rect 12713 8313 12725 8347
rect 12759 8344 12771 8347
rect 12894 8344 12900 8356
rect 12759 8316 12900 8344
rect 12759 8313 12771 8316
rect 12713 8307 12771 8313
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 2682 8276 2688 8288
rect 2643 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 2958 8236 2964 8288
rect 3016 8236 3022 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 9030 8276 9036 8288
rect 7800 8248 9036 8276
rect 7800 8236 7806 8248
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 13096 8276 13124 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13262 8412 13268 8424
rect 13223 8384 13268 8412
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 10836 8248 13124 8276
rect 10836 8236 10842 8248
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 13372 8276 13400 8375
rect 13228 8248 13400 8276
rect 13228 8236 13234 8248
rect 1104 8186 13892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 13892 8186
rect 1104 8112 13892 8134
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 2406 8072 2412 8084
rect 1535 8044 2412 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6604 8044 6653 8072
rect 6604 8032 6610 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 2958 7936 2964 7948
rect 1452 7908 2964 7936
rect 1452 7896 1458 7908
rect 2958 7896 2964 7908
rect 3016 7936 3022 7948
rect 3237 7939 3295 7945
rect 3237 7936 3249 7939
rect 3016 7908 3249 7936
rect 3016 7896 3022 7908
rect 3237 7905 3249 7908
rect 3283 7905 3295 7939
rect 3237 7899 3295 7905
rect 4614 7896 4620 7948
rect 4672 7936 4678 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 4672 7908 6101 7936
rect 4672 7896 4678 7908
rect 6089 7905 6101 7908
rect 6135 7936 6147 7939
rect 6178 7936 6184 7948
rect 6135 7908 6184 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6656 7936 6684 8035
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 7064 8044 7113 8072
rect 7064 8032 7070 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 7101 8035 7159 8041
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9030 8072 9036 8084
rect 8803 8044 9036 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 9723 8044 10364 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 6917 8007 6975 8013
rect 6917 7973 6929 8007
rect 6963 8004 6975 8007
rect 8018 8004 8024 8016
rect 6963 7976 8024 8004
rect 6963 7973 6975 7976
rect 6917 7967 6975 7973
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 8389 8007 8447 8013
rect 8389 7973 8401 8007
rect 8435 8004 8447 8007
rect 9217 8007 9275 8013
rect 9217 8004 9229 8007
rect 8435 7976 9229 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 9217 7973 9229 7976
rect 9263 8004 9275 8007
rect 9263 7976 9674 8004
rect 9263 7973 9275 7976
rect 9217 7967 9275 7973
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 6656 7908 7573 7936
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7561 7899 7619 7905
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8570 7936 8576 7948
rect 8312 7908 8576 7936
rect 3418 7868 3424 7880
rect 3379 7840 3424 7868
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 1946 7760 1952 7812
rect 2004 7760 2010 7812
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 2961 7803 3019 7809
rect 2961 7800 2973 7803
rect 2740 7772 2973 7800
rect 2740 7760 2746 7772
rect 2961 7769 2973 7772
rect 3007 7769 3019 7803
rect 5353 7803 5411 7809
rect 2961 7763 3019 7769
rect 3620 7772 4186 7800
rect 3620 7741 3648 7772
rect 5353 7769 5365 7803
rect 5399 7769 5411 7803
rect 5353 7763 5411 7769
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7701 3663 7735
rect 3878 7732 3884 7744
rect 3839 7704 3884 7732
rect 3605 7695 3663 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 5368 7732 5396 7763
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 5644 7800 5672 7831
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 5905 7871 5963 7877
rect 5776 7840 5821 7868
rect 5776 7828 5782 7840
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 7469 7871 7527 7877
rect 5951 7840 7420 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 5500 7772 5672 7800
rect 7392 7800 7420 7840
rect 7469 7837 7481 7871
rect 7515 7868 7527 7871
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7515 7840 7941 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8312 7877 8340 7908
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 8772 7908 9444 7936
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 8076 7840 8217 7868
rect 8076 7828 8082 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7864 8539 7871
rect 8772 7868 8800 7908
rect 9416 7880 9444 7908
rect 8588 7864 8800 7868
rect 8527 7840 8800 7864
rect 8527 7837 8616 7840
rect 8481 7836 8616 7837
rect 8481 7831 8539 7836
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 9088 7840 9137 7868
rect 9088 7828 9094 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9306 7868 9312 7880
rect 9267 7840 9312 7868
rect 9125 7831 9183 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9646 7868 9674 7976
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 9456 7840 9501 7868
rect 9646 7840 9873 7868
rect 9456 7828 9462 7840
rect 9861 7837 9873 7840
rect 9907 7868 9919 7871
rect 9950 7868 9956 7880
rect 9907 7840 9956 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 10100 7840 10241 7868
rect 10100 7828 10106 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 9582 7800 9588 7812
rect 7392 7772 9588 7800
rect 5500 7760 5506 7772
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 10336 7800 10364 8044
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 10928 8044 11621 8072
rect 10928 8032 10934 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12437 8075 12495 8081
rect 12437 8072 12449 8075
rect 12032 8044 12449 8072
rect 12032 8032 12038 8044
rect 12437 8041 12449 8044
rect 12483 8072 12495 8075
rect 13170 8072 13176 8084
rect 12483 8044 13176 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 10413 8007 10471 8013
rect 10413 7973 10425 8007
rect 10459 8004 10471 8007
rect 11882 8004 11888 8016
rect 10459 7976 11888 8004
rect 10459 7973 10471 7976
rect 10413 7967 10471 7973
rect 11882 7964 11888 7976
rect 11940 7964 11946 8016
rect 12253 8007 12311 8013
rect 12253 7973 12265 8007
rect 12299 8004 12311 8007
rect 12618 8004 12624 8016
rect 12299 7976 12624 8004
rect 12299 7973 12311 7976
rect 12253 7967 12311 7973
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 10778 7896 10784 7948
rect 10836 7936 10842 7948
rect 10836 7908 11008 7936
rect 10836 7896 10842 7908
rect 10980 7877 11008 7908
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 11572 7908 11805 7936
rect 11572 7896 11578 7908
rect 11793 7905 11805 7908
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 13078 7936 13084 7948
rect 12391 7908 13084 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 13188 7936 13216 8032
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13188 7908 13369 7936
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11425 7871 11483 7877
rect 11112 7840 11157 7868
rect 11112 7828 11118 7840
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11974 7868 11980 7880
rect 11471 7840 11980 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 12759 7840 13277 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 13265 7837 13277 7840
rect 13311 7868 13323 7871
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13311 7840 14105 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 13173 7803 13231 7809
rect 13173 7800 13185 7803
rect 10336 7772 13185 7800
rect 13173 7769 13185 7772
rect 13219 7769 13231 7803
rect 13173 7763 13231 7769
rect 4028 7704 5396 7732
rect 4028 7692 4034 7704
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7064 7704 7109 7732
rect 7064 7692 7070 7704
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 7984 7704 10057 7732
rect 7984 7692 7990 7704
rect 10045 7701 10057 7704
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 10781 7735 10839 7741
rect 10192 7704 10237 7732
rect 10192 7692 10198 7704
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 10962 7732 10968 7744
rect 10827 7704 10968 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 12805 7735 12863 7741
rect 12805 7732 12817 7735
rect 12768 7704 12817 7732
rect 12768 7692 12774 7704
rect 12805 7701 12817 7704
rect 12851 7701 12863 7735
rect 12805 7695 12863 7701
rect 1104 7642 13892 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 13892 7642
rect 1104 7568 13892 7590
rect 2958 7488 2964 7540
rect 3016 7528 3022 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 3016 7500 3157 7528
rect 3016 7488 3022 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 8662 7528 8668 7540
rect 3145 7491 3203 7497
rect 4908 7500 8668 7528
rect 2222 7420 2228 7472
rect 2280 7420 2286 7472
rect 3513 7463 3571 7469
rect 3513 7429 3525 7463
rect 3559 7460 3571 7463
rect 3878 7460 3884 7472
rect 3559 7432 3884 7460
rect 3559 7429 3571 7432
rect 3513 7423 3571 7429
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 3108 7364 3341 7392
rect 3108 7352 3114 7364
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2314 7324 2320 7336
rect 1719 7296 2320 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 3620 7324 3648 7355
rect 3694 7352 3700 7404
rect 3752 7401 3758 7404
rect 3752 7392 3760 7401
rect 4433 7395 4491 7401
rect 3752 7364 3797 7392
rect 3752 7355 3760 7364
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 4433 7355 4491 7361
rect 3752 7352 3758 7355
rect 3786 7324 3792 7336
rect 2464 7296 3792 7324
rect 2464 7284 2470 7296
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 3881 7259 3939 7265
rect 3881 7225 3893 7259
rect 3927 7256 3939 7259
rect 3970 7256 3976 7268
rect 3927 7228 3976 7256
rect 3927 7225 3939 7228
rect 3881 7219 3939 7225
rect 3970 7216 3976 7228
rect 4028 7216 4034 7268
rect 4448 7256 4476 7355
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 4908 7392 4936 7500
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 9490 7528 9496 7540
rect 9447 7500 9496 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 10134 7528 10140 7540
rect 10060 7500 10140 7528
rect 5718 7460 5724 7472
rect 5000 7432 5724 7460
rect 5000 7401 5028 7432
rect 5718 7420 5724 7432
rect 5776 7420 5782 7472
rect 5810 7420 5816 7472
rect 5868 7460 5874 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 5868 7432 6653 7460
rect 5868 7420 5874 7432
rect 4847 7364 4936 7392
rect 4985 7395 5043 7401
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5224 7364 5549 7392
rect 5224 7352 5230 7364
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5902 7392 5908 7404
rect 5863 7364 5908 7392
rect 5537 7355 5595 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6380 7401 6408 7432
rect 6641 7429 6653 7432
rect 6687 7429 6699 7463
rect 6641 7423 6699 7429
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 7834 7460 7840 7472
rect 7064 7432 7840 7460
rect 7064 7420 7070 7432
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 9030 7460 9036 7472
rect 8076 7432 8340 7460
rect 8943 7432 9036 7460
rect 8076 7420 8082 7432
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7392 7251 7395
rect 7466 7392 7472 7404
rect 7239 7364 7472 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 4706 7324 4712 7336
rect 4667 7296 4712 7324
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 4614 7256 4620 7268
rect 4448 7228 4620 7256
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 5460 7256 5488 7287
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 6012 7324 6040 7355
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 8110 7392 8116 7404
rect 8071 7364 8116 7392
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8312 7401 8340 7432
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8343 7364 8769 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 8757 7361 8769 7364
rect 8803 7392 8815 7395
rect 8846 7392 8852 7404
rect 8803 7364 8852 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 5684 7296 6040 7324
rect 5684 7284 5690 7296
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 7926 7324 7932 7336
rect 7432 7296 7932 7324
rect 7432 7284 7438 7296
rect 7926 7284 7932 7296
rect 7984 7324 7990 7336
rect 8220 7324 8248 7355
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 8956 7324 8984 7432
rect 9030 7420 9036 7432
rect 9088 7460 9094 7472
rect 10060 7460 10088 7500
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10962 7528 10968 7540
rect 10923 7500 10968 7528
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11146 7488 11152 7540
rect 11204 7528 11210 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 11204 7500 11345 7528
rect 11204 7488 11210 7500
rect 11333 7497 11345 7500
rect 11379 7497 11391 7531
rect 11333 7491 11391 7497
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 11974 7528 11980 7540
rect 11747 7500 11980 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 11716 7460 11744 7491
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12805 7531 12863 7537
rect 12805 7497 12817 7531
rect 12851 7528 12863 7531
rect 14001 7531 14059 7537
rect 14001 7528 14013 7531
rect 12851 7500 14013 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 14001 7497 14013 7500
rect 14047 7497 14059 7531
rect 14001 7491 14059 7497
rect 9088 7432 10088 7460
rect 10796 7432 11744 7460
rect 11885 7463 11943 7469
rect 9088 7420 9094 7432
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9398 7392 9404 7404
rect 9171 7364 9404 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9398 7352 9404 7364
rect 9456 7392 9462 7404
rect 9677 7395 9735 7401
rect 9677 7392 9689 7395
rect 9456 7364 9689 7392
rect 9456 7352 9462 7364
rect 9677 7361 9689 7364
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9824 7364 9873 7392
rect 9824 7352 9830 7364
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9950 7352 9956 7404
rect 10008 7392 10014 7404
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 10008 7364 10149 7392
rect 10008 7352 10014 7364
rect 10137 7361 10149 7364
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 7984 7296 8248 7324
rect 8864 7296 8984 7324
rect 9033 7327 9091 7333
rect 7984 7284 7990 7296
rect 8018 7256 8024 7268
rect 5460 7228 8024 7256
rect 8018 7216 8024 7228
rect 8076 7216 8082 7268
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3418 7188 3424 7200
rect 2832 7160 3424 7188
rect 2832 7148 2838 7160
rect 3418 7148 3424 7160
rect 3476 7188 3482 7200
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 3476 7160 4077 7188
rect 3476 7148 3482 7160
rect 4065 7157 4077 7160
rect 4111 7157 4123 7191
rect 5074 7188 5080 7200
rect 5035 7160 5080 7188
rect 4065 7151 4123 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5810 7188 5816 7200
rect 5771 7160 5816 7188
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 6086 7188 6092 7200
rect 6047 7160 6092 7188
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6512 7160 6561 7188
rect 6512 7148 6518 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 6549 7151 6607 7157
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 8864 7197 8892 7296
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9214 7324 9220 7336
rect 9079 7296 9220 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 10796 7333 10824 7432
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 11931 7432 12480 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 12452 7401 12480 7432
rect 12345 7395 12403 7401
rect 12345 7392 12357 7395
rect 11204 7364 12357 7392
rect 11204 7352 11210 7364
rect 12345 7361 12357 7364
rect 12391 7361 12403 7395
rect 12345 7355 12403 7361
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7392 12495 7395
rect 12802 7392 12808 7404
rect 12483 7364 12808 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 13170 7392 13176 7404
rect 13131 7364 13176 7392
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 13998 7392 14004 7404
rect 13311 7364 14004 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 10962 7324 10968 7336
rect 10919 7296 10968 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 12032 7296 12541 7324
rect 12032 7284 12038 7296
rect 12529 7293 12541 7296
rect 12575 7324 12587 7327
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 12575 7296 13369 7324
rect 12575 7293 12587 7296
rect 12529 7287 12587 7293
rect 13280 7268 13308 7296
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 10045 7259 10103 7265
rect 10045 7225 10057 7259
rect 10091 7256 10103 7259
rect 10134 7256 10140 7268
rect 10091 7228 10140 7256
rect 10091 7225 10103 7228
rect 10045 7219 10103 7225
rect 10134 7216 10140 7228
rect 10192 7216 10198 7268
rect 13262 7216 13268 7268
rect 13320 7216 13326 7268
rect 8849 7191 8907 7197
rect 8849 7188 8861 7191
rect 8628 7160 8861 7188
rect 8628 7148 8634 7160
rect 8849 7157 8861 7160
rect 8895 7157 8907 7191
rect 8849 7151 8907 7157
rect 8941 7191 8999 7197
rect 8941 7157 8953 7191
rect 8987 7188 8999 7191
rect 9030 7188 9036 7200
rect 8987 7160 9036 7188
rect 8987 7157 8999 7160
rect 8941 7151 8999 7157
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 11974 7188 11980 7200
rect 11935 7160 11980 7188
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 1104 7098 13892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 13892 7098
rect 1104 7024 13892 7046
rect 2222 6984 2228 6996
rect 2183 6956 2228 6984
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 2924 6956 3433 6984
rect 2924 6944 2930 6956
rect 3421 6953 3433 6956
rect 3467 6953 3479 6987
rect 3421 6947 3479 6953
rect 4341 6987 4399 6993
rect 4341 6953 4353 6987
rect 4387 6984 4399 6987
rect 4614 6984 4620 6996
rect 4387 6956 4620 6984
rect 4387 6953 4399 6956
rect 4341 6947 4399 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 5708 6987 5766 6993
rect 5708 6953 5720 6987
rect 5754 6984 5766 6987
rect 5810 6984 5816 6996
rect 5754 6956 5816 6984
rect 5754 6953 5766 6956
rect 5708 6947 5766 6953
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 10042 6984 10048 6996
rect 9364 6956 10048 6984
rect 9364 6944 9370 6956
rect 2314 6916 2320 6928
rect 2275 6888 2320 6916
rect 2314 6876 2320 6888
rect 2372 6876 2378 6928
rect 3053 6919 3111 6925
rect 3053 6885 3065 6919
rect 3099 6916 3111 6919
rect 3326 6916 3332 6928
rect 3099 6888 3332 6916
rect 3099 6885 3111 6888
rect 3053 6879 3111 6885
rect 3326 6876 3332 6888
rect 3384 6916 3390 6928
rect 3602 6916 3608 6928
rect 3384 6888 3608 6916
rect 3384 6876 3390 6888
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 3786 6916 3792 6928
rect 3747 6888 3792 6916
rect 3786 6876 3792 6888
rect 3844 6876 3850 6928
rect 4982 6916 4988 6928
rect 4943 6888 4988 6916
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 7834 6916 7840 6928
rect 7795 6888 7840 6916
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 8754 6916 8760 6928
rect 8496 6888 8760 6916
rect 2976 6820 4200 6848
rect 2976 6792 3004 6820
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2501 6783 2559 6789
rect 2087 6752 2176 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2148 6644 2176 6752
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2958 6780 2964 6792
rect 2547 6752 2964 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 3200 6752 3433 6780
rect 3200 6740 3206 6752
rect 3421 6749 3433 6752
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3786 6780 3792 6792
rect 3651 6752 3792 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4172 6789 4200 6820
rect 4430 6808 4436 6860
rect 4488 6848 4494 6860
rect 4617 6851 4675 6857
rect 4617 6848 4629 6851
rect 4488 6820 4629 6848
rect 4488 6808 4494 6820
rect 4617 6817 4629 6820
rect 4663 6848 4675 6851
rect 5166 6848 5172 6860
rect 4663 6820 5172 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8496 6848 8524 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9677 6919 9735 6925
rect 9677 6916 9689 6919
rect 9088 6888 9689 6916
rect 9088 6876 9094 6888
rect 9677 6885 9689 6888
rect 9723 6885 9735 6919
rect 9677 6879 9735 6885
rect 9766 6876 9772 6928
rect 9824 6876 9830 6928
rect 8251 6820 8524 6848
rect 8573 6851 8631 6857
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 9122 6848 9128 6860
rect 8619 6820 9128 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 9784 6848 9812 6876
rect 9600 6820 9812 6848
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3936 6752 4077 6780
rect 3936 6740 3942 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 4893 6783 4951 6789
rect 4893 6749 4905 6783
rect 4939 6749 4951 6783
rect 5074 6780 5080 6792
rect 5035 6752 5080 6780
rect 4893 6743 4951 6749
rect 2685 6715 2743 6721
rect 2685 6681 2697 6715
rect 2731 6712 2743 6715
rect 3053 6715 3111 6721
rect 3053 6712 3065 6715
rect 2731 6684 3065 6712
rect 2731 6681 2743 6684
rect 2685 6675 2743 6681
rect 3053 6681 3065 6684
rect 3099 6681 3111 6715
rect 4706 6712 4712 6724
rect 3053 6675 3111 6681
rect 3252 6684 4712 6712
rect 2774 6644 2780 6656
rect 2148 6616 2780 6644
rect 2774 6604 2780 6616
rect 2832 6644 2838 6656
rect 3252 6653 3280 6684
rect 4706 6672 4712 6684
rect 4764 6672 4770 6724
rect 3237 6647 3295 6653
rect 2832 6616 2925 6644
rect 2832 6604 2838 6616
rect 3237 6613 3249 6647
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3878 6644 3884 6656
rect 3752 6616 3884 6644
rect 3752 6604 3758 6616
rect 3878 6604 3884 6616
rect 3936 6644 3942 6656
rect 3973 6647 4031 6653
rect 3973 6644 3985 6647
rect 3936 6616 3985 6644
rect 3936 6604 3942 6616
rect 3973 6613 3985 6616
rect 4019 6613 4031 6647
rect 4816 6644 4844 6743
rect 4908 6712 4936 6743
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 5442 6780 5448 6792
rect 5316 6752 5448 6780
rect 5316 6740 5322 6752
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 7466 6780 7472 6792
rect 7423 6752 7472 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 9600 6789 9628 6820
rect 9876 6789 9904 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10965 6987 11023 6993
rect 10965 6953 10977 6987
rect 11011 6984 11023 6987
rect 11054 6984 11060 6996
rect 11011 6956 11060 6984
rect 11011 6953 11023 6956
rect 10965 6947 11023 6953
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10226 6848 10232 6860
rect 10008 6820 10232 6848
rect 10008 6808 10014 6820
rect 10226 6808 10232 6820
rect 10284 6848 10290 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 10284 6820 10333 6848
rect 10284 6808 10290 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 11701 6851 11759 6857
rect 11701 6817 11713 6851
rect 11747 6848 11759 6851
rect 11882 6848 11888 6860
rect 11747 6820 11888 6848
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6780 8539 6783
rect 8665 6783 8723 6789
rect 8527 6752 8616 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 5718 6712 5724 6724
rect 4908 6684 5724 6712
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 6454 6672 6460 6724
rect 6512 6672 6518 6724
rect 7834 6672 7840 6724
rect 7892 6712 7898 6724
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 7892 6684 7941 6712
rect 7892 6672 7898 6684
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 8404 6712 8432 6743
rect 8588 6712 8616 6752
rect 8665 6749 8677 6783
rect 8711 6780 8723 6783
rect 9585 6783 9643 6789
rect 9585 6780 9597 6783
rect 8711 6752 9597 6780
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 9585 6749 9597 6752
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6780 10195 6783
rect 11146 6780 11152 6792
rect 10183 6752 11152 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 9784 6712 9812 6743
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 12894 6780 12900 6792
rect 12855 6752 12900 6780
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 10042 6712 10048 6724
rect 8404 6684 8524 6712
rect 8588 6684 10048 6712
rect 7929 6675 7987 6681
rect 4890 6644 4896 6656
rect 4816 6616 4896 6644
rect 3973 6607 4031 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7374 6644 7380 6656
rect 7239 6616 7380 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 8496 6644 8524 6684
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 11330 6712 11336 6724
rect 11072 6684 11336 6712
rect 9030 6644 9036 6656
rect 8496 6616 9036 6644
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 10376 6616 10517 6644
rect 10376 6604 10382 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10505 6607 10563 6613
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 11072 6653 11100 6684
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 13354 6672 13360 6724
rect 13412 6712 13418 6724
rect 13541 6715 13599 6721
rect 13541 6712 13553 6715
rect 13412 6684 13553 6712
rect 13412 6672 13418 6684
rect 13541 6681 13553 6684
rect 13587 6681 13599 6715
rect 13541 6675 13599 6681
rect 11057 6647 11115 6653
rect 10652 6616 10697 6644
rect 10652 6604 10658 6616
rect 11057 6613 11069 6647
rect 11103 6613 11115 6647
rect 11422 6644 11428 6656
rect 11383 6616 11428 6644
rect 11057 6607 11115 6613
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11572 6616 11617 6644
rect 11572 6604 11578 6616
rect 1104 6554 13892 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 13892 6554
rect 1104 6480 13892 6502
rect 3970 6440 3976 6452
rect 3528 6412 3976 6440
rect 2314 6332 2320 6384
rect 2372 6332 2378 6384
rect 3528 6372 3556 6412
rect 3970 6400 3976 6412
rect 4028 6440 4034 6452
rect 5626 6440 5632 6452
rect 4028 6412 5120 6440
rect 4028 6400 4034 6412
rect 3436 6344 3556 6372
rect 3436 6313 3464 6344
rect 3786 6332 3792 6384
rect 3844 6372 3850 6384
rect 3844 6344 5028 6372
rect 3844 6332 3850 6344
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3602 6304 3608 6316
rect 3563 6276 3608 6304
rect 3421 6267 3479 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 3927 6276 4016 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 1719 6208 3709 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3988 6168 4016 6276
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 4120 6276 4261 6304
rect 4120 6264 4126 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 4706 6304 4712 6316
rect 4663 6276 4712 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 4540 6236 4568 6267
rect 4706 6264 4712 6276
rect 4764 6264 4770 6316
rect 4540 6208 4660 6236
rect 4632 6180 4660 6208
rect 4798 6196 4804 6248
rect 4856 6196 4862 6248
rect 4430 6168 4436 6180
rect 3988 6140 4436 6168
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 4614 6128 4620 6180
rect 4672 6128 4678 6180
rect 4816 6168 4844 6196
rect 4724 6140 4844 6168
rect 5000 6168 5028 6344
rect 5092 6313 5120 6412
rect 5368 6412 5632 6440
rect 5368 6381 5396 6412
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 5902 6440 5908 6452
rect 5767 6412 5908 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6052 6412 6745 6440
rect 6052 6400 6058 6412
rect 6733 6409 6745 6412
rect 6779 6440 6791 6443
rect 6779 6412 7972 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 5353 6375 5411 6381
rect 5353 6341 5365 6375
rect 5399 6341 5411 6375
rect 5353 6335 5411 6341
rect 5445 6375 5503 6381
rect 5445 6341 5457 6375
rect 5491 6372 5503 6375
rect 6086 6372 6092 6384
rect 5491 6344 6092 6372
rect 5491 6341 5503 6344
rect 5445 6335 5503 6341
rect 6086 6332 6092 6344
rect 6144 6332 6150 6384
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 6564 6344 7849 6372
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 5225 6307 5283 6313
rect 5225 6273 5237 6307
rect 5271 6304 5283 6307
rect 5583 6307 5641 6313
rect 5271 6273 5304 6304
rect 5225 6267 5304 6273
rect 5583 6273 5595 6307
rect 5629 6304 5641 6307
rect 5810 6304 5816 6316
rect 5629 6276 5816 6304
rect 5629 6273 5641 6276
rect 5583 6267 5641 6273
rect 5276 6236 5304 6267
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 5997 6307 6055 6313
rect 5997 6304 6009 6307
rect 5960 6276 6009 6304
rect 5960 6264 5966 6276
rect 5997 6273 6009 6276
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6564 6236 6592 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 7944 6372 7972 6412
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 8076 6412 8401 6440
rect 8076 6400 8082 6412
rect 8389 6409 8401 6412
rect 8435 6440 8447 6443
rect 8938 6440 8944 6452
rect 8435 6412 8944 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 10226 6440 10232 6452
rect 9088 6412 10232 6440
rect 9088 6400 9094 6412
rect 10152 6381 10180 6412
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 10594 6440 10600 6452
rect 10428 6412 10600 6440
rect 9953 6375 10011 6381
rect 9953 6372 9965 6375
rect 7944 6344 9965 6372
rect 7837 6335 7895 6341
rect 9953 6341 9965 6344
rect 9999 6341 10011 6375
rect 9953 6335 10011 6341
rect 10137 6375 10195 6381
rect 10137 6341 10149 6375
rect 10183 6372 10195 6375
rect 10183 6344 10217 6372
rect 10183 6341 10195 6344
rect 10137 6335 10195 6341
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6696 6276 6837 6304
rect 6696 6264 6702 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 7282 6304 7288 6316
rect 7243 6276 7288 6304
rect 6825 6267 6883 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7432 6276 7481 6304
rect 7432 6264 7438 6276
rect 7469 6273 7481 6276
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 5276 6208 6592 6236
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 7760 6236 7788 6267
rect 8018 6264 8024 6316
rect 8076 6304 8082 6316
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 8076 6276 8217 6304
rect 8076 6264 8082 6276
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8846 6304 8852 6316
rect 8807 6276 8852 6304
rect 8205 6267 8263 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9398 6304 9404 6316
rect 9263 6276 9404 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 10318 6304 10324 6316
rect 10279 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10428 6313 10456 6412
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11514 6440 11520 6452
rect 11379 6412 11520 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 10778 6372 10784 6384
rect 10739 6344 10784 6372
rect 10778 6332 10784 6344
rect 10836 6332 10842 6384
rect 10870 6332 10876 6384
rect 10928 6372 10934 6384
rect 11149 6375 11207 6381
rect 11149 6372 11161 6375
rect 10928 6344 11161 6372
rect 10928 6332 10934 6344
rect 11149 6341 11161 6344
rect 11195 6372 11207 6375
rect 11882 6372 11888 6384
rect 11195 6344 11888 6372
rect 11195 6341 11207 6344
rect 11149 6335 11207 6341
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 12529 6375 12587 6381
rect 12529 6341 12541 6375
rect 12575 6372 12587 6375
rect 12894 6372 12900 6384
rect 12575 6344 12900 6372
rect 12575 6341 12587 6344
rect 12529 6335 12587 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 13081 6375 13139 6381
rect 13081 6341 13093 6375
rect 13127 6372 13139 6375
rect 13354 6372 13360 6384
rect 13127 6344 13360 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 11609 6307 11667 6313
rect 11609 6273 11621 6307
rect 11655 6304 11667 6307
rect 11698 6304 11704 6316
rect 11655 6276 11704 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 9030 6236 9036 6248
rect 7064 6208 7109 6236
rect 7208 6208 7788 6236
rect 8991 6208 9036 6236
rect 7064 6196 7070 6208
rect 5994 6168 6000 6180
rect 5000 6140 6000 6168
rect 3142 6100 3148 6112
rect 3103 6072 3148 6100
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 3878 6060 3884 6112
rect 3936 6100 3942 6112
rect 4341 6103 4399 6109
rect 4341 6100 4353 6103
rect 3936 6072 4353 6100
rect 3936 6060 3942 6072
rect 4341 6069 4353 6072
rect 4387 6100 4399 6103
rect 4724 6100 4752 6140
rect 5994 6128 6000 6140
rect 6052 6128 6058 6180
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 7208 6168 7236 6208
rect 9030 6196 9036 6208
rect 9088 6196 9094 6248
rect 10428 6236 10456 6267
rect 9140 6208 10456 6236
rect 9140 6168 9168 6208
rect 6512 6140 7236 6168
rect 7392 6140 9168 6168
rect 9493 6171 9551 6177
rect 6512 6128 6518 6140
rect 4387 6072 4752 6100
rect 4801 6103 4859 6109
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 5350 6100 5356 6112
rect 4847 6072 5356 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6362 6100 6368 6112
rect 6323 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7392 6100 7420 6140
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 10502 6168 10508 6180
rect 9539 6140 10508 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 7558 6100 7564 6112
rect 6972 6072 7420 6100
rect 7519 6072 7564 6100
rect 6972 6060 6978 6072
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 8021 6103 8079 6109
rect 8021 6100 8033 6103
rect 7892 6072 8033 6100
rect 7892 6060 7898 6072
rect 8021 6069 8033 6072
rect 8067 6069 8079 6103
rect 8021 6063 8079 6069
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8628 6072 8953 6100
rect 8628 6060 8634 6072
rect 8941 6069 8953 6072
rect 8987 6069 8999 6103
rect 9122 6100 9128 6112
rect 9083 6072 9128 6100
rect 8941 6063 8999 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9398 6100 9404 6112
rect 9272 6072 9404 6100
rect 9272 6060 9278 6072
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10612 6100 10640 6267
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 12066 6264 12072 6316
rect 12124 6304 12130 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 12124 6276 12265 6304
rect 12124 6264 12130 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12032 6208 12633 6236
rect 12032 6196 12038 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 12860 6208 13185 6236
rect 12860 6196 12866 6208
rect 13173 6205 13185 6208
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 10870 6100 10876 6112
rect 10284 6072 10640 6100
rect 10831 6072 10876 6100
rect 10284 6060 10290 6072
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 13446 6100 13452 6112
rect 13407 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 1104 6010 13892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 13892 6010
rect 1104 5936 13892 5958
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 3602 5896 3608 5908
rect 3283 5868 3608 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 4617 5899 4675 5905
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 4706 5896 4712 5908
rect 4663 5868 4712 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5896 4859 5899
rect 4982 5896 4988 5908
rect 4847 5868 4988 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5626 5896 5632 5908
rect 5215 5868 5632 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6641 5899 6699 5905
rect 6641 5896 6653 5899
rect 5736 5868 6653 5896
rect 2774 5828 2780 5840
rect 2148 5800 2780 5828
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 2148 5701 2176 5800
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 3513 5831 3571 5837
rect 3513 5797 3525 5831
rect 3559 5828 3571 5831
rect 4062 5828 4068 5840
rect 3559 5800 4068 5828
rect 3559 5797 3571 5800
rect 3513 5791 3571 5797
rect 4062 5788 4068 5800
rect 4120 5828 4126 5840
rect 4120 5800 4568 5828
rect 4120 5788 4126 5800
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5729 3019 5763
rect 3878 5760 3884 5772
rect 3839 5732 3884 5760
rect 2961 5723 3019 5729
rect 2133 5695 2191 5701
rect 2133 5692 2145 5695
rect 1820 5664 2145 5692
rect 1820 5652 1826 5664
rect 2133 5661 2145 5664
rect 2179 5661 2191 5695
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2133 5655 2191 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 2976 5624 3004 5723
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 4540 5769 4568 5800
rect 4890 5788 4896 5840
rect 4948 5828 4954 5840
rect 5736 5828 5764 5868
rect 6641 5865 6653 5868
rect 6687 5896 6699 5899
rect 7006 5896 7012 5908
rect 6687 5868 7012 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7282 5896 7288 5908
rect 7243 5868 7288 5896
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 9490 5896 9496 5908
rect 7616 5868 9168 5896
rect 9451 5868 9496 5896
rect 7616 5856 7622 5868
rect 4948 5800 5764 5828
rect 4948 5788 4954 5800
rect 5810 5788 5816 5840
rect 5868 5828 5874 5840
rect 6181 5831 6239 5837
rect 6181 5828 6193 5831
rect 5868 5800 6193 5828
rect 5868 5788 5874 5800
rect 6181 5797 6193 5800
rect 6227 5828 6239 5831
rect 6454 5828 6460 5840
rect 6227 5800 6460 5828
rect 6227 5797 6239 5800
rect 6181 5791 6239 5797
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 6914 5828 6920 5840
rect 6875 5800 6920 5828
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 5718 5760 5724 5772
rect 5675 5732 5724 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3421 5695 3479 5701
rect 3421 5692 3433 5695
rect 3200 5664 3433 5692
rect 3200 5652 3206 5664
rect 3421 5661 3433 5664
rect 3467 5692 3479 5695
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3467 5664 3985 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4356 5624 4384 5723
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 5994 5720 6000 5772
rect 6052 5760 6058 5772
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 6052 5732 6377 5760
rect 6052 5720 6058 5732
rect 6365 5729 6377 5732
rect 6411 5760 6423 5763
rect 7300 5760 7328 5856
rect 7469 5831 7527 5837
rect 7469 5797 7481 5831
rect 7515 5828 7527 5831
rect 7650 5828 7656 5840
rect 7515 5800 7656 5828
rect 7515 5797 7527 5800
rect 7469 5791 7527 5797
rect 7650 5788 7656 5800
rect 7708 5788 7714 5840
rect 8128 5837 8156 5868
rect 8113 5831 8171 5837
rect 8113 5797 8125 5831
rect 8159 5797 8171 5831
rect 8113 5791 8171 5797
rect 8665 5831 8723 5837
rect 8665 5797 8677 5831
rect 8711 5828 8723 5831
rect 8757 5831 8815 5837
rect 8757 5828 8769 5831
rect 8711 5800 8769 5828
rect 8711 5797 8723 5800
rect 8665 5791 8723 5797
rect 8757 5797 8769 5800
rect 8803 5828 8815 5831
rect 8938 5828 8944 5840
rect 8803 5800 8944 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 9033 5831 9091 5837
rect 9033 5797 9045 5831
rect 9079 5797 9091 5831
rect 9033 5791 9091 5797
rect 6411 5732 7328 5760
rect 6411 5729 6423 5732
rect 6365 5723 6423 5729
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7800 5732 8217 5760
rect 7800 5720 7806 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 9048 5760 9076 5791
rect 8205 5723 8263 5729
rect 8312 5732 9076 5760
rect 9140 5760 9168 5868
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 9861 5899 9919 5905
rect 9732 5868 9777 5896
rect 9732 5856 9738 5868
rect 9861 5865 9873 5899
rect 9907 5896 9919 5899
rect 10410 5896 10416 5908
rect 9907 5868 9941 5896
rect 10371 5868 10416 5896
rect 9907 5865 9919 5868
rect 9861 5859 9919 5865
rect 9876 5828 9904 5859
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 12802 5896 12808 5908
rect 10520 5868 11192 5896
rect 10042 5828 10048 5840
rect 9646 5800 10048 5828
rect 9646 5760 9674 5800
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10520 5828 10548 5868
rect 10284 5800 10548 5828
rect 10284 5788 10290 5800
rect 10594 5788 10600 5840
rect 10652 5828 10658 5840
rect 10778 5828 10784 5840
rect 10652 5800 10784 5828
rect 10652 5788 10658 5800
rect 10778 5788 10784 5800
rect 10836 5828 10842 5840
rect 10836 5800 11008 5828
rect 10836 5788 10842 5800
rect 10980 5769 11008 5800
rect 10965 5763 11023 5769
rect 9140 5732 9674 5760
rect 9876 5732 10916 5760
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 5537 5695 5595 5701
rect 4479 5664 5488 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 4614 5624 4620 5636
rect 2976 5596 4620 5624
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 2409 5559 2467 5565
rect 2409 5556 2421 5559
rect 1820 5528 2421 5556
rect 1820 5516 1826 5528
rect 2409 5525 2421 5528
rect 2455 5525 2467 5559
rect 2409 5519 2467 5525
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 5258 5556 5264 5568
rect 3384 5528 5264 5556
rect 3384 5516 3390 5528
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 5460 5556 5488 5664
rect 5537 5661 5549 5695
rect 5583 5692 5595 5695
rect 6178 5692 6184 5704
rect 5583 5664 6040 5692
rect 6139 5664 6184 5692
rect 5583 5661 5595 5664
rect 5537 5655 5595 5661
rect 5810 5624 5816 5636
rect 5771 5596 5816 5624
rect 5810 5584 5816 5596
rect 5868 5584 5874 5636
rect 6012 5624 6040 5664
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 6549 5695 6607 5701
rect 6549 5694 6561 5695
rect 6472 5692 6561 5694
rect 6328 5666 6561 5692
rect 6328 5664 6500 5666
rect 6328 5652 6334 5664
rect 6549 5661 6561 5666
rect 6595 5661 6607 5695
rect 7190 5692 7196 5704
rect 6549 5655 6607 5661
rect 6656 5664 7196 5692
rect 6656 5624 6684 5664
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7282 5652 7288 5704
rect 7340 5692 7346 5704
rect 8312 5701 8340 5732
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 7340 5664 7389 5692
rect 7340 5652 7346 5664
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8662 5692 8668 5704
rect 8527 5664 8668 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 6012 5596 6684 5624
rect 6914 5584 6920 5636
rect 6972 5584 6978 5636
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 8036 5624 8064 5655
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9214 5692 9220 5704
rect 8904 5664 9220 5692
rect 8904 5652 8910 5664
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9876 5701 9904 5732
rect 9861 5695 9919 5701
rect 9861 5692 9873 5695
rect 9364 5664 9873 5692
rect 9364 5652 9370 5664
rect 9861 5661 9873 5664
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5692 10103 5695
rect 10226 5692 10232 5704
rect 10091 5664 10232 5692
rect 10091 5661 10103 5664
rect 10045 5655 10103 5661
rect 9493 5627 9551 5633
rect 9493 5624 9505 5627
rect 7064 5596 9505 5624
rect 7064 5584 7070 5596
rect 6932 5556 6960 5584
rect 9048 5568 9076 5596
rect 9493 5593 9505 5596
rect 9539 5624 9551 5627
rect 10060 5624 10088 5655
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10410 5692 10416 5704
rect 10367 5664 10416 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10888 5692 10916 5732
rect 10965 5729 10977 5763
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 11054 5692 11060 5704
rect 10888 5664 11060 5692
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11164 5692 11192 5868
rect 11532 5868 12434 5896
rect 12763 5868 12808 5896
rect 11532 5837 11560 5868
rect 11517 5831 11575 5837
rect 11517 5797 11529 5831
rect 11563 5797 11575 5831
rect 11517 5791 11575 5797
rect 12066 5788 12072 5840
rect 12124 5828 12130 5840
rect 12161 5831 12219 5837
rect 12161 5828 12173 5831
rect 12124 5800 12173 5828
rect 12124 5788 12130 5800
rect 12161 5797 12173 5800
rect 12207 5797 12219 5831
rect 12406 5828 12434 5868
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 13587 5868 14013 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14001 5859 14059 5865
rect 13170 5828 13176 5840
rect 12406 5800 13176 5828
rect 12161 5791 12219 5797
rect 12176 5760 12204 5791
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 12176 5732 12434 5760
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 11164 5664 11253 5692
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5661 11483 5695
rect 11698 5692 11704 5704
rect 11659 5664 11704 5692
rect 11425 5655 11483 5661
rect 11440 5624 11468 5655
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 9539 5596 10088 5624
rect 10244 5596 11468 5624
rect 12253 5627 12311 5633
rect 9539 5593 9551 5596
rect 9493 5587 9551 5593
rect 7834 5556 7840 5568
rect 5460 5528 6960 5556
rect 7795 5528 7840 5556
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 8110 5516 8116 5568
rect 8168 5556 8174 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8168 5528 8769 5556
rect 8168 5516 8174 5528
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 9030 5516 9036 5568
rect 9088 5516 9094 5568
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 10244 5565 10272 5596
rect 12253 5593 12265 5627
rect 12299 5593 12311 5627
rect 12406 5624 12434 5732
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5692 12679 5695
rect 12894 5692 12900 5704
rect 12667 5664 12900 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 12406 5596 12725 5624
rect 12253 5587 12311 5593
rect 12713 5593 12725 5596
rect 12759 5593 12771 5627
rect 13170 5624 13176 5636
rect 13131 5596 13176 5624
rect 12713 5587 12771 5593
rect 10229 5559 10287 5565
rect 10229 5556 10241 5559
rect 10008 5528 10241 5556
rect 10008 5516 10014 5528
rect 10229 5525 10241 5528
rect 10275 5525 10287 5559
rect 10778 5556 10784 5568
rect 10739 5528 10784 5556
rect 10229 5519 10287 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 10870 5516 10876 5568
rect 10928 5556 10934 5568
rect 12268 5556 12296 5587
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 12437 5559 12495 5565
rect 12437 5556 12449 5559
rect 10928 5528 10973 5556
rect 12268 5528 12449 5556
rect 10928 5516 10934 5528
rect 12437 5525 12449 5528
rect 12483 5525 12495 5559
rect 12986 5556 12992 5568
rect 12947 5528 12992 5556
rect 12437 5519 12495 5525
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 1104 5466 13892 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 13892 5466
rect 1104 5392 13892 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 2866 5352 2872 5364
rect 1535 5324 2872 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3881 5355 3939 5361
rect 3881 5321 3893 5355
rect 3927 5352 3939 5355
rect 4706 5352 4712 5364
rect 3927 5324 4712 5352
rect 3927 5321 3939 5324
rect 3881 5315 3939 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 5718 5352 5724 5364
rect 5583 5324 5724 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6178 5312 6184 5364
rect 6236 5312 6242 5364
rect 7650 5352 7656 5364
rect 6288 5324 7656 5352
rect 1946 5244 1952 5296
rect 2004 5244 2010 5296
rect 2884 5284 2912 5312
rect 5626 5284 5632 5296
rect 2884 5256 3832 5284
rect 3804 5225 3832 5256
rect 4172 5256 4936 5284
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4172 5225 4200 5256
rect 4908 5225 4936 5256
rect 5000 5256 5632 5284
rect 5000 5225 5028 5256
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 6196 5284 6224 5312
rect 5736 5256 6224 5284
rect 4157 5219 4215 5225
rect 4157 5216 4169 5219
rect 4120 5188 4169 5216
rect 4120 5176 4126 5188
rect 4157 5185 4169 5188
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 2958 5148 2964 5160
rect 2919 5120 2964 5148
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 3326 5148 3332 5160
rect 3283 5120 3332 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 4356 5148 4384 5179
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 5316 5188 5365 5216
rect 5316 5176 5322 5188
rect 5353 5185 5365 5188
rect 5399 5216 5411 5219
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5399 5188 5457 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 5445 5185 5457 5188
rect 5491 5216 5503 5219
rect 5736 5216 5764 5256
rect 5994 5216 6000 5228
rect 5491 5188 5764 5216
rect 5955 5188 6000 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6288 5216 6316 5324
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 7834 5352 7840 5364
rect 7795 5324 7840 5352
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 8662 5352 8668 5364
rect 8623 5324 8668 5352
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9214 5352 9220 5364
rect 8864 5324 9220 5352
rect 6457 5287 6515 5293
rect 6457 5253 6469 5287
rect 6503 5284 6515 5287
rect 6546 5284 6552 5296
rect 6503 5256 6552 5284
rect 6503 5253 6515 5256
rect 6457 5247 6515 5253
rect 6546 5244 6552 5256
rect 6604 5244 6610 5296
rect 7009 5287 7067 5293
rect 7009 5253 7021 5287
rect 7055 5284 7067 5287
rect 7282 5284 7288 5296
rect 7055 5256 7288 5284
rect 7055 5253 7067 5256
rect 7009 5247 7067 5253
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 7392 5256 7604 5284
rect 6227 5188 6316 5216
rect 6641 5219 6699 5225
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7190 5216 7196 5228
rect 6871 5188 7196 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 5074 5148 5080 5160
rect 4356 5120 5080 5148
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5148 5227 5151
rect 6086 5148 6092 5160
rect 5215 5120 6092 5148
rect 5215 5117 5227 5120
rect 5169 5111 5227 5117
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6656 5148 6684 5179
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7392 5225 7420 5256
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 7466 5176 7472 5228
rect 7524 5176 7530 5228
rect 6512 5120 7328 5148
rect 6512 5108 6518 5120
rect 4525 5083 4583 5089
rect 4525 5049 4537 5083
rect 4571 5080 4583 5083
rect 5810 5080 5816 5092
rect 4571 5052 5816 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6638 5080 6644 5092
rect 5951 5052 6644 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 4709 5015 4767 5021
rect 4709 4981 4721 5015
rect 4755 5012 4767 5015
rect 4890 5012 4896 5024
rect 4755 4984 4896 5012
rect 4755 4981 4767 4984
rect 4709 4975 4767 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 7300 5021 7328 5120
rect 7484 5089 7512 5176
rect 7576 5148 7604 5256
rect 8864 5216 8892 5324
rect 9214 5312 9220 5324
rect 9272 5352 9278 5364
rect 10778 5352 10784 5364
rect 9272 5324 10784 5352
rect 9272 5312 9278 5324
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11698 5352 11704 5364
rect 11379 5324 11704 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 10962 5284 10968 5296
rect 9732 5256 9777 5284
rect 9732 5244 9738 5256
rect 8920 5219 8978 5225
rect 8920 5216 8932 5219
rect 7760 5188 8248 5216
rect 8864 5188 8932 5216
rect 7650 5148 7656 5160
rect 7576 5120 7656 5148
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 7469 5083 7527 5089
rect 7469 5049 7481 5083
rect 7515 5049 7527 5083
rect 7469 5043 7527 5049
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7760 5012 7788 5188
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 8110 5148 8116 5160
rect 8071 5120 8116 5148
rect 7929 5111 7987 5117
rect 7944 5080 7972 5111
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 8220 5148 8248 5188
rect 8920 5185 8932 5188
rect 8966 5185 8978 5219
rect 8920 5179 8978 5185
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9490 5216 9496 5228
rect 9447 5188 9496 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 9490 5176 9496 5188
rect 9548 5216 9554 5228
rect 9861 5219 9919 5225
rect 9548 5206 9812 5216
rect 9861 5206 9873 5219
rect 9548 5188 9873 5206
rect 9548 5176 9554 5188
rect 9784 5185 9873 5188
rect 9907 5185 9919 5219
rect 10134 5210 10140 5262
rect 10192 5210 10198 5262
rect 10923 5256 10968 5284
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 11112 5256 11744 5284
rect 11112 5244 11118 5256
rect 9784 5179 9919 5185
rect 10136 5185 10148 5210
rect 10182 5185 10194 5210
rect 10136 5179 10194 5185
rect 9784 5178 9904 5179
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 10778 5216 10784 5228
rect 10376 5188 10784 5216
rect 10376 5186 10456 5188
rect 10376 5176 10382 5186
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 11146 5216 11152 5228
rect 10919 5188 11152 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 11514 5216 11520 5228
rect 11475 5188 11520 5216
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 11716 5225 11744 5256
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12710 5216 12716 5228
rect 12023 5188 12716 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13446 5216 13452 5228
rect 13407 5188 13452 5216
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 9217 5151 9275 5157
rect 9217 5148 9229 5151
rect 8220 5120 9229 5148
rect 9217 5117 9229 5120
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 8481 5083 8539 5089
rect 8481 5080 8493 5083
rect 7944 5052 8493 5080
rect 8481 5049 8493 5052
rect 8527 5080 8539 5083
rect 8846 5080 8852 5092
rect 8527 5052 8852 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 8846 5040 8852 5052
rect 8904 5040 8910 5092
rect 8938 5040 8944 5092
rect 8996 5080 9002 5092
rect 9125 5083 9183 5089
rect 9125 5080 9137 5083
rect 8996 5052 9137 5080
rect 8996 5040 9002 5052
rect 9125 5049 9137 5052
rect 9171 5049 9183 5083
rect 9232 5080 9260 5111
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 9674 5148 9680 5160
rect 9640 5120 9680 5148
rect 9640 5108 9646 5120
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 10091 5120 10456 5148
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 10428 5092 10456 5120
rect 10594 5108 10600 5160
rect 10652 5148 10658 5160
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 10652 5120 10701 5148
rect 10652 5108 10658 5120
rect 10689 5117 10701 5120
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 9953 5083 10011 5089
rect 9953 5080 9965 5083
rect 9232 5052 9965 5080
rect 9125 5043 9183 5049
rect 9953 5049 9965 5052
rect 9999 5049 10011 5083
rect 9953 5043 10011 5049
rect 10134 5040 10140 5092
rect 10192 5040 10198 5092
rect 10410 5040 10416 5092
rect 10468 5040 10474 5092
rect 11146 5080 11152 5092
rect 10888 5052 11152 5080
rect 7331 4984 7788 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 7984 4984 9045 5012
rect 7984 4972 7990 4984
rect 9033 4981 9045 4984
rect 9079 4981 9091 5015
rect 9033 4975 9091 4981
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 9766 5012 9772 5024
rect 9640 4984 9772 5012
rect 9640 4972 9646 4984
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10152 5012 10180 5040
rect 10226 5012 10232 5024
rect 10152 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 10505 5015 10563 5021
rect 10505 4981 10517 5015
rect 10551 5012 10563 5015
rect 10888 5012 10916 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 13078 5040 13084 5092
rect 13136 5080 13142 5092
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 13136 5052 13277 5080
rect 13136 5040 13142 5052
rect 13265 5049 13277 5052
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 10551 4984 10916 5012
rect 10551 4981 10563 4984
rect 10505 4975 10563 4981
rect 10962 4972 10968 5024
rect 11020 5012 11026 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11020 4984 11805 5012
rect 11020 4972 11026 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 11793 4975 11851 4981
rect 1104 4922 13892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 13892 4922
rect 1104 4848 13892 4870
rect 1946 4768 1952 4820
rect 2004 4808 2010 4820
rect 2041 4811 2099 4817
rect 2041 4808 2053 4811
rect 2004 4780 2053 4808
rect 2004 4768 2010 4780
rect 2041 4777 2053 4780
rect 2087 4777 2099 4811
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2041 4771 2099 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4120 4780 4629 4808
rect 4120 4768 4126 4780
rect 4356 4752 4384 4780
rect 4617 4777 4629 4780
rect 4663 4777 4675 4811
rect 4617 4771 4675 4777
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 6457 4811 6515 4817
rect 6457 4808 6469 4811
rect 5132 4780 6469 4808
rect 5132 4768 5138 4780
rect 6457 4777 6469 4780
rect 6503 4777 6515 4811
rect 6457 4771 6515 4777
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7926 4808 7932 4820
rect 7064 4780 7932 4808
rect 7064 4768 7070 4780
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8021 4811 8079 4817
rect 8021 4777 8033 4811
rect 8067 4808 8079 4811
rect 8938 4808 8944 4820
rect 8067 4780 8944 4808
rect 8067 4777 8079 4780
rect 8021 4771 8079 4777
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9214 4808 9220 4820
rect 9175 4780 9220 4808
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 10962 4808 10968 4820
rect 10652 4780 10968 4808
rect 10652 4768 10658 4780
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 4338 4700 4344 4752
rect 4396 4700 4402 4752
rect 5902 4740 5908 4752
rect 5000 4712 5908 4740
rect 2682 4672 2688 4684
rect 2332 4644 2688 4672
rect 2332 4613 2360 4644
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 3050 4672 3056 4684
rect 3011 4644 3056 4672
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4641 3571 4675
rect 3513 4635 3571 4641
rect 1857 4607 1915 4613
rect 1857 4604 1869 4607
rect 1780 4576 1869 4604
rect 1780 4480 1808 4576
rect 1857 4573 1869 4576
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2866 4604 2872 4616
rect 2639 4576 2872 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3418 4604 3424 4616
rect 3379 4576 3424 4604
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3528 4604 3556 4635
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4229 4675 4287 4681
rect 4229 4672 4241 4675
rect 4120 4644 4241 4672
rect 4120 4632 4126 4644
rect 4229 4641 4241 4644
rect 4275 4672 4287 4675
rect 4275 4644 4483 4672
rect 4275 4641 4287 4644
rect 4229 4635 4287 4641
rect 4455 4604 4483 4644
rect 4522 4632 4528 4684
rect 4580 4672 4586 4684
rect 4580 4644 4625 4672
rect 4580 4632 4586 4644
rect 5000 4613 5028 4712
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 5997 4743 6055 4749
rect 5997 4709 6009 4743
rect 6043 4740 6055 4743
rect 7098 4740 7104 4752
rect 6043 4712 7104 4740
rect 6043 4709 6055 4712
rect 5997 4703 6055 4709
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 7650 4700 7656 4752
rect 7708 4740 7714 4752
rect 7837 4743 7895 4749
rect 7837 4740 7849 4743
rect 7708 4712 7849 4740
rect 7708 4700 7714 4712
rect 7837 4709 7849 4712
rect 7883 4709 7895 4743
rect 8294 4740 8300 4752
rect 7837 4703 7895 4709
rect 7944 4712 8300 4740
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 3528 4576 4108 4604
rect 4455 4576 4997 4604
rect 3786 4536 3792 4548
rect 3747 4508 3792 4536
rect 3786 4496 3792 4508
rect 3844 4496 3850 4548
rect 3970 4536 3976 4548
rect 3931 4508 3976 4536
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 4080 4536 4108 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 5092 4604 5120 4635
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 6638 4672 6644 4684
rect 5224 4644 5580 4672
rect 6599 4644 6644 4672
rect 5224 4632 5230 4644
rect 5258 4604 5264 4616
rect 5092 4576 5264 4604
rect 4985 4567 5043 4573
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5442 4604 5448 4616
rect 5403 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5552 4604 5580 4644
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 7006 4632 7012 4684
rect 7064 4632 7070 4684
rect 7944 4672 7972 4712
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8389 4743 8447 4749
rect 8389 4709 8401 4743
rect 8435 4740 8447 4743
rect 9398 4740 9404 4752
rect 8435 4712 9404 4740
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 9493 4743 9551 4749
rect 9493 4709 9505 4743
rect 9539 4740 9551 4743
rect 10410 4740 10416 4752
rect 9539 4712 10416 4740
rect 9539 4709 9551 4712
rect 9493 4703 9551 4709
rect 10410 4700 10416 4712
rect 10468 4740 10474 4752
rect 11514 4740 11520 4752
rect 10468 4712 11520 4740
rect 10468 4700 10474 4712
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 13078 4740 13084 4752
rect 13039 4712 13084 4740
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 8662 4672 8668 4684
rect 7392 4644 7972 4672
rect 8220 4644 8668 4672
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5552 4576 5641 4604
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 6178 4604 6184 4616
rect 5951 4576 6184 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4604 6331 4607
rect 6454 4604 6460 4616
rect 6319 4576 6460 4604
rect 6319 4573 6331 4576
rect 6273 4567 6331 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6730 4604 6736 4616
rect 6691 4576 6736 4604
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 7024 4604 7052 4632
rect 7392 4613 7420 4644
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 7024 4576 7113 4604
rect 6917 4567 6975 4573
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4573 7435 4607
rect 7742 4604 7748 4616
rect 7703 4576 7748 4604
rect 7377 4567 7435 4573
rect 5994 4536 6000 4548
rect 4080 4508 6000 4536
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 6840 4536 6868 4567
rect 6696 4508 6868 4536
rect 6696 4496 6702 4508
rect 1762 4468 1768 4480
rect 1723 4440 1768 4468
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 2225 4471 2283 4477
rect 2225 4437 2237 4471
rect 2271 4468 2283 4471
rect 2958 4468 2964 4480
rect 2271 4440 2964 4468
rect 2271 4437 2283 4440
rect 2225 4431 2283 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 4246 4468 4252 4480
rect 3292 4440 4252 4468
rect 3292 4428 3298 4440
rect 4246 4428 4252 4440
rect 4304 4468 4310 4480
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 4304 4440 4353 4468
rect 4304 4428 4310 4440
rect 4341 4437 4353 4440
rect 4387 4437 4399 4471
rect 4341 4431 4399 4437
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4468 4491 4471
rect 5810 4468 5816 4480
rect 4479 4440 5816 4468
rect 4479 4437 4491 4440
rect 4433 4431 4491 4437
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 6932 4468 6960 4567
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 8134 4607 8192 4613
rect 8134 4573 8146 4607
rect 8180 4604 8192 4607
rect 8220 4604 8248 4644
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 10244 4644 10456 4672
rect 8180 4576 8248 4604
rect 8180 4573 8192 4576
rect 8134 4567 8192 4573
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8352 4576 8585 4604
rect 8352 4564 8358 4576
rect 8573 4573 8585 4576
rect 8619 4604 8631 4607
rect 8754 4604 8760 4616
rect 8619 4576 8760 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9401 4607 9459 4613
rect 9401 4606 9413 4607
rect 9324 4604 9413 4606
rect 9088 4578 9413 4604
rect 9088 4576 9352 4578
rect 9088 4564 9094 4576
rect 9401 4573 9413 4578
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 7006 4496 7012 4548
rect 7064 4536 7070 4548
rect 7193 4539 7251 4545
rect 7193 4536 7205 4539
rect 7064 4508 7205 4536
rect 7064 4496 7070 4508
rect 7193 4505 7205 4508
rect 7239 4505 7251 4539
rect 7558 4536 7564 4548
rect 7519 4508 7564 4536
rect 7193 4499 7251 4505
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 7760 4536 7788 4564
rect 8665 4539 8723 4545
rect 8665 4536 8677 4539
rect 7760 4508 8677 4536
rect 8665 4505 8677 4508
rect 8711 4536 8723 4539
rect 9600 4536 9628 4635
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 9766 4604 9772 4616
rect 9723 4576 9772 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 9950 4604 9956 4616
rect 9907 4576 9956 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10244 4613 10272 4644
rect 10428 4616 10456 4644
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 10873 4675 10931 4681
rect 10873 4672 10885 4675
rect 10652 4644 10885 4672
rect 10652 4632 10658 4644
rect 10873 4641 10885 4644
rect 10919 4641 10931 4675
rect 10873 4635 10931 4641
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 12621 4675 12679 4681
rect 11379 4644 12204 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 10336 4536 10364 4567
rect 10410 4564 10416 4616
rect 10468 4564 10474 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 10778 4604 10784 4616
rect 10735 4576 10784 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 8711 4508 9628 4536
rect 9876 4508 10364 4536
rect 8711 4505 8723 4508
rect 8665 4499 8723 4505
rect 9490 4468 9496 4480
rect 6144 4440 9496 4468
rect 6144 4428 6150 4440
rect 9490 4428 9496 4440
rect 9548 4468 9554 4480
rect 9876 4468 9904 4508
rect 10042 4468 10048 4480
rect 9548 4440 9904 4468
rect 10003 4440 10048 4468
rect 9548 4428 9554 4440
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10520 4468 10548 4567
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 10888 4604 10916 4635
rect 12176 4613 12204 4644
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12710 4672 12716 4684
rect 12667 4644 12716 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 13170 4672 13176 4684
rect 13131 4644 13176 4672
rect 13170 4632 13176 4644
rect 13228 4632 13234 4684
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 10888 4576 11529 4604
rect 11517 4573 11529 4576
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 13446 4604 13452 4616
rect 12483 4576 13452 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 11425 4539 11483 4545
rect 11425 4505 11437 4539
rect 11471 4505 11483 4539
rect 12176 4536 12204 4567
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 12986 4536 12992 4548
rect 12176 4508 12992 4536
rect 11425 4499 11483 4505
rect 10284 4440 10548 4468
rect 10284 4428 10290 4440
rect 10686 4428 10692 4480
rect 10744 4468 10750 4480
rect 10962 4468 10968 4480
rect 10744 4440 10968 4468
rect 10744 4428 10750 4440
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11440 4468 11468 4499
rect 12986 4496 12992 4508
rect 13044 4496 13050 4548
rect 13265 4471 13323 4477
rect 13265 4468 13277 4471
rect 11440 4440 13277 4468
rect 13265 4437 13277 4440
rect 13311 4437 13323 4471
rect 13265 4431 13323 4437
rect 1104 4378 13892 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 13892 4378
rect 1104 4304 13892 4326
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 3234 4264 3240 4276
rect 2740 4236 3240 4264
rect 2740 4224 2746 4236
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 3970 4264 3976 4276
rect 3344 4236 3976 4264
rect 3344 4205 3372 4236
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4522 4264 4528 4276
rect 4304 4236 4528 4264
rect 4304 4224 4310 4236
rect 4522 4224 4528 4236
rect 4580 4264 4586 4276
rect 4982 4264 4988 4276
rect 4580 4236 4988 4264
rect 4580 4224 4586 4236
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 5169 4267 5227 4273
rect 5169 4233 5181 4267
rect 5215 4264 5227 4267
rect 5442 4264 5448 4276
rect 5215 4236 5448 4264
rect 5215 4233 5227 4236
rect 5169 4227 5227 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 5718 4264 5724 4276
rect 5675 4236 5724 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 6089 4267 6147 4273
rect 6089 4233 6101 4267
rect 6135 4264 6147 4267
rect 6730 4264 6736 4276
rect 6135 4236 6736 4264
rect 6135 4233 6147 4236
rect 6089 4227 6147 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 7650 4264 7656 4276
rect 7024 4236 7656 4264
rect 7024 4208 7052 4236
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 8481 4267 8539 4273
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 8662 4264 8668 4276
rect 8527 4236 8668 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 8662 4224 8668 4236
rect 8720 4224 8726 4276
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 9272 4236 10456 4264
rect 9272 4224 9278 4236
rect 10428 4208 10456 4236
rect 3329 4199 3387 4205
rect 3329 4165 3341 4199
rect 3375 4165 3387 4199
rect 5074 4196 5080 4208
rect 3329 4159 3387 4165
rect 4080 4168 5080 4196
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 2225 4131 2283 4137
rect 2225 4128 2237 4131
rect 1820 4100 2237 4128
rect 1820 4088 1826 4100
rect 2225 4097 2237 4100
rect 2271 4128 2283 4131
rect 3050 4128 3056 4140
rect 2271 4100 2636 4128
rect 3011 4100 3056 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2608 4001 2636 4100
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 2958 4069 2964 4072
rect 2941 4063 2964 4069
rect 2941 4029 2953 4063
rect 3016 4060 3022 4072
rect 3344 4060 3372 4159
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4080 4128 4108 4168
rect 5074 4156 5080 4168
rect 5132 4156 5138 4208
rect 7006 4196 7012 4208
rect 5552 4168 7012 4196
rect 4019 4100 4108 4128
rect 4157 4131 4215 4137
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4157 4097 4169 4131
rect 4203 4128 4215 4131
rect 4338 4128 4344 4140
rect 4203 4100 4344 4128
rect 4203 4097 4215 4100
rect 4157 4091 4215 4097
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4128 4491 4131
rect 4522 4128 4528 4140
rect 4479 4100 4528 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4614 4088 4620 4140
rect 4672 4128 4678 4140
rect 4798 4128 4804 4140
rect 4672 4100 4717 4128
rect 4759 4100 4804 4128
rect 4672 4088 4678 4100
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5552 4137 5580 4168
rect 7006 4156 7012 4168
rect 7064 4156 7070 4208
rect 7558 4156 7564 4208
rect 7616 4196 7622 4208
rect 9677 4199 9735 4205
rect 7616 4168 9628 4196
rect 7616 4156 7622 4168
rect 5537 4131 5595 4137
rect 4948 4100 4993 4128
rect 4948 4088 4954 4100
rect 5537 4097 5549 4131
rect 5583 4097 5595 4131
rect 5994 4128 6000 4140
rect 5955 4100 6000 4128
rect 5537 4091 5595 4097
rect 3016 4032 3372 4060
rect 2941 4023 2964 4029
rect 2958 4020 2964 4023
rect 3016 4020 3022 4032
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 5552 4060 5580 4091
rect 5994 4088 6000 4100
rect 6052 4128 6058 4140
rect 6052 4100 6408 4128
rect 6052 4088 6058 4100
rect 3476 4032 5580 4060
rect 3476 4020 3482 4032
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 6380 4069 6408 4100
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6512 4100 6745 4128
rect 6512 4088 6518 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7248 4100 7389 4128
rect 7248 4088 7254 4100
rect 7377 4097 7389 4100
rect 7423 4128 7435 4131
rect 7742 4128 7748 4140
rect 7423 4100 7748 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5684 4032 5733 4060
rect 5684 4020 5690 4032
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 6365 4063 6423 4069
rect 6365 4029 6377 4063
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 6822 4060 6828 4072
rect 6687 4032 6828 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 2593 3995 2651 4001
rect 2593 3961 2605 3995
rect 2639 3992 2651 3995
rect 3142 3992 3148 4004
rect 2639 3964 3148 3992
rect 2639 3961 2651 3964
rect 2593 3955 2651 3961
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 4430 3992 4436 4004
rect 4111 3964 4436 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 4430 3952 4436 3964
rect 4488 3952 4494 4004
rect 4614 3992 4620 4004
rect 4575 3964 4620 3992
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 6178 3952 6184 4004
rect 6236 3992 6242 4004
rect 6656 3992 6684 4023
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 7156 4032 7297 4060
rect 7156 4020 7162 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 6236 3964 6684 3992
rect 6236 3952 6242 3964
rect 2406 3924 2412 3936
rect 2367 3896 2412 3924
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2832 3896 2877 3924
rect 2832 3884 2838 3896
rect 4706 3884 4712 3936
rect 4764 3924 4770 3936
rect 4985 3927 5043 3933
rect 4985 3924 4997 3927
rect 4764 3896 4997 3924
rect 4764 3884 4770 3896
rect 4985 3893 4997 3896
rect 5031 3893 5043 3927
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 4985 3887 5043 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7650 3924 7656 3936
rect 7611 3896 7656 3924
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 7852 3924 7880 4091
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8168 4100 8953 4128
rect 8168 4088 8174 4100
rect 8312 4069 8340 4100
rect 8941 4097 8953 4100
rect 8987 4128 8999 4131
rect 9030 4128 9036 4140
rect 8987 4100 9036 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 9490 4128 9496 4140
rect 9451 4100 9496 4128
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 9600 4137 9628 4168
rect 9677 4165 9689 4199
rect 9723 4165 9735 4199
rect 9677 4159 9735 4165
rect 9861 4199 9919 4205
rect 9861 4165 9873 4199
rect 9907 4196 9919 4199
rect 10134 4196 10140 4208
rect 9907 4168 10140 4196
rect 9907 4165 9919 4168
rect 9861 4159 9919 4165
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4097 9643 4131
rect 9692 4128 9720 4159
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 10321 4199 10379 4205
rect 10321 4165 10333 4199
rect 10367 4165 10379 4199
rect 10321 4159 10379 4165
rect 9950 4128 9956 4140
rect 9692 4100 9956 4128
rect 9585 4091 9643 4097
rect 9950 4088 9956 4100
rect 10008 4128 10014 4140
rect 10226 4128 10232 4140
rect 10008 4100 10232 4128
rect 10008 4088 10014 4100
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10336 4128 10364 4159
rect 10410 4156 10416 4208
rect 10468 4196 10474 4208
rect 10505 4199 10563 4205
rect 10505 4196 10517 4199
rect 10468 4168 10517 4196
rect 10468 4156 10474 4168
rect 10505 4165 10517 4168
rect 10551 4165 10563 4199
rect 10505 4159 10563 4165
rect 13078 4156 13084 4208
rect 13136 4196 13142 4208
rect 13265 4199 13323 4205
rect 13265 4196 13277 4199
rect 13136 4168 13277 4196
rect 13136 4156 13142 4168
rect 13265 4165 13277 4168
rect 13311 4165 13323 4199
rect 13265 4159 13323 4165
rect 10336 4100 10456 4128
rect 10428 4072 10456 4100
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 11054 4128 11060 4140
rect 10744 4100 11060 4128
rect 10744 4088 10750 4100
rect 11054 4088 11060 4100
rect 11112 4128 11118 4140
rect 11241 4131 11299 4137
rect 11241 4128 11253 4131
rect 11112 4100 11253 4128
rect 11112 4088 11118 4100
rect 11241 4097 11253 4100
rect 11287 4128 11299 4131
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11287 4100 11529 4128
rect 11287 4097 11299 4100
rect 11241 4091 11299 4097
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12802 4128 12808 4140
rect 11931 4100 12480 4128
rect 12763 4100 12808 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4029 8355 4063
rect 8297 4023 8355 4029
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 8570 4060 8576 4072
rect 8435 4032 8576 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 8570 4020 8576 4032
rect 8628 4060 8634 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8628 4032 9137 4060
rect 8628 4020 8634 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10410 4060 10416 4072
rect 9732 4032 10416 4060
rect 9732 4020 9738 4032
rect 10410 4020 10416 4032
rect 10468 4060 10474 4072
rect 10468 4032 10561 4060
rect 10468 4020 10474 4032
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 12032 4032 12173 4060
rect 12032 4020 12038 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 8849 3995 8907 4001
rect 8849 3961 8861 3995
rect 8895 3992 8907 3995
rect 10594 3992 10600 4004
rect 8895 3964 10600 3992
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10689 3995 10747 4001
rect 10689 3961 10701 3995
rect 10735 3992 10747 3995
rect 11422 3992 11428 4004
rect 10735 3964 11428 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 7800 3896 7941 3924
rect 7800 3884 7806 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 9858 3924 9864 3936
rect 9819 3896 9864 3924
rect 7929 3887 7987 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 11054 3924 11060 3936
rect 10091 3896 11060 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 12066 3924 12072 3936
rect 12027 3896 12072 3924
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 12452 3924 12480 4100
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4060 12771 4063
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12759 4032 12909 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3992 12679 3995
rect 13262 3992 13268 4004
rect 12667 3964 13268 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 13262 3952 13268 3964
rect 13320 3952 13326 4004
rect 13170 3924 13176 3936
rect 12452 3896 13176 3924
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 1104 3834 13892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 13892 3834
rect 1104 3760 13892 3782
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 3418 3720 3424 3732
rect 3283 3692 3424 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4157 3723 4215 3729
rect 4157 3689 4169 3723
rect 4203 3720 4215 3723
rect 4203 3692 4476 3720
rect 4203 3689 4215 3692
rect 4157 3683 4215 3689
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3584 1823 3587
rect 2774 3584 2780 3596
rect 1811 3556 2780 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4028 3556 4384 3584
rect 4028 3544 4034 3556
rect 1486 3516 1492 3528
rect 1447 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 4356 3525 4384 3556
rect 4448 3525 4476 3692
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4856 3692 4997 3720
rect 4856 3680 4862 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 4985 3683 5043 3689
rect 6546 3680 6552 3732
rect 6604 3720 6610 3732
rect 6604 3692 9628 3720
rect 6604 3680 6610 3692
rect 4890 3612 4896 3664
rect 4948 3612 4954 3664
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 9600 3652 9628 3692
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 11146 3720 11152 3732
rect 9732 3692 9777 3720
rect 10060 3692 11152 3720
rect 9732 3680 9738 3692
rect 10060 3652 10088 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 8812 3624 9168 3652
rect 9600 3624 10088 3652
rect 8812 3612 8818 3624
rect 4908 3584 4936 3612
rect 4540 3556 4936 3584
rect 5169 3587 5227 3593
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4434 3519 4492 3525
rect 4434 3485 4446 3519
rect 4480 3485 4492 3519
rect 4434 3479 4492 3485
rect 2406 3408 2412 3460
rect 2464 3408 2470 3460
rect 4264 3380 4292 3479
rect 4540 3448 4568 3556
rect 5169 3553 5181 3587
rect 5215 3553 5227 3587
rect 5169 3547 5227 3553
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 5718 3584 5724 3596
rect 5491 3556 5724 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 4706 3516 4712 3528
rect 4667 3488 4712 3516
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 4845 3519 4903 3525
rect 4845 3485 4857 3519
rect 4891 3516 4903 3519
rect 5184 3516 5212 3547
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 7006 3584 7012 3596
rect 6595 3556 7012 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3584 8079 3587
rect 8772 3584 8800 3612
rect 9030 3584 9036 3596
rect 8067 3556 8800 3584
rect 8991 3556 9036 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 4891 3488 5212 3516
rect 5537 3519 5595 3525
rect 4891 3485 4903 3488
rect 4845 3479 4903 3485
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 4617 3451 4675 3457
rect 4617 3448 4629 3451
rect 4540 3420 4629 3448
rect 4617 3417 4629 3420
rect 4663 3417 4675 3451
rect 4617 3411 4675 3417
rect 4862 3380 4890 3479
rect 5552 3448 5580 3479
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 6144 3488 6285 3516
rect 6144 3476 6150 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8501 3519 8559 3525
rect 8501 3516 8513 3519
rect 8352 3488 8513 3516
rect 8352 3476 8358 3488
rect 8501 3485 8513 3488
rect 8547 3485 8559 3519
rect 8501 3479 8559 3485
rect 5718 3448 5724 3460
rect 5552 3420 5724 3448
rect 5718 3408 5724 3420
rect 5776 3448 5782 3460
rect 6178 3448 6184 3460
rect 5776 3420 6184 3448
rect 5776 3408 5782 3420
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 8110 3408 8116 3460
rect 8168 3448 8174 3460
rect 8205 3451 8263 3457
rect 8205 3448 8217 3451
rect 8168 3420 8217 3448
rect 8168 3408 8174 3420
rect 8205 3417 8217 3420
rect 8251 3417 8263 3451
rect 8205 3411 8263 3417
rect 8389 3451 8447 3457
rect 8389 3417 8401 3451
rect 8435 3448 8447 3451
rect 8588 3448 8616 3556
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9140 3584 9168 3624
rect 10134 3612 10140 3664
rect 10192 3661 10198 3664
rect 10192 3652 10199 3661
rect 10192 3624 10237 3652
rect 10192 3615 10199 3624
rect 10192 3612 10198 3615
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 10505 3655 10563 3661
rect 10505 3652 10517 3655
rect 10468 3624 10517 3652
rect 10468 3612 10474 3624
rect 10505 3621 10517 3624
rect 10551 3621 10563 3655
rect 13262 3652 13268 3664
rect 13223 3624 13268 3652
rect 10505 3615 10563 3621
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 9490 3584 9496 3596
rect 9140 3556 9496 3584
rect 9490 3544 9496 3556
rect 9548 3584 9554 3596
rect 10229 3587 10287 3593
rect 10229 3584 10241 3587
rect 9548 3556 10241 3584
rect 9548 3544 9554 3556
rect 10229 3553 10241 3556
rect 10275 3553 10287 3587
rect 10229 3547 10287 3553
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8757 3519 8815 3525
rect 8757 3516 8769 3519
rect 8720 3488 8769 3516
rect 8720 3476 8726 3488
rect 8757 3485 8769 3488
rect 8803 3516 8815 3519
rect 9950 3516 9956 3528
rect 8803 3488 9956 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 9950 3476 9956 3488
rect 10008 3516 10014 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 10008 3488 10057 3516
rect 10008 3476 10014 3488
rect 10045 3485 10057 3488
rect 10091 3516 10103 3519
rect 10334 3519 10392 3525
rect 10091 3488 10272 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 10134 3448 10140 3460
rect 8435 3420 8616 3448
rect 8680 3420 10140 3448
rect 8435 3417 8447 3420
rect 8389 3411 8447 3417
rect 4264 3352 4890 3380
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 7524 3352 8585 3380
rect 7524 3340 7530 3352
rect 8573 3349 8585 3352
rect 8619 3380 8631 3383
rect 8680 3380 8708 3420
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 10244 3448 10272 3488
rect 10334 3485 10346 3519
rect 10380 3516 10392 3519
rect 10428 3516 10456 3612
rect 11882 3584 11888 3596
rect 11716 3556 11888 3584
rect 10380 3488 10456 3516
rect 10965 3519 11023 3525
rect 10380 3485 10392 3488
rect 10334 3479 10392 3485
rect 10965 3485 10977 3519
rect 11011 3516 11023 3519
rect 11146 3516 11152 3528
rect 11011 3488 11152 3516
rect 11011 3485 11023 3488
rect 10965 3479 11023 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11716 3525 11744 3556
rect 11882 3544 11888 3556
rect 11940 3584 11946 3596
rect 12802 3584 12808 3596
rect 11940 3556 12808 3584
rect 11940 3544 11946 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3485 11759 3519
rect 11974 3516 11980 3528
rect 11935 3488 11980 3516
rect 11701 3479 11759 3485
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 13170 3516 13176 3528
rect 13131 3488 13176 3516
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 10594 3448 10600 3460
rect 10244 3420 10600 3448
rect 10594 3408 10600 3420
rect 10652 3448 10658 3460
rect 10689 3451 10747 3457
rect 10689 3448 10701 3451
rect 10652 3420 10701 3448
rect 10652 3408 10658 3420
rect 10689 3417 10701 3420
rect 10735 3417 10747 3451
rect 10689 3411 10747 3417
rect 10873 3451 10931 3457
rect 10873 3417 10885 3451
rect 10919 3417 10931 3451
rect 10873 3411 10931 3417
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3448 11943 3451
rect 13188 3448 13216 3476
rect 11931 3420 13216 3448
rect 11931 3417 11943 3420
rect 11885 3411 11943 3417
rect 8619 3352 8708 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 9180 3352 9229 3380
rect 9180 3340 9186 3352
rect 9217 3349 9229 3352
rect 9263 3349 9275 3383
rect 9217 3343 9275 3349
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9364 3352 9409 3380
rect 9364 3340 9370 3352
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9732 3352 9873 3380
rect 9732 3340 9738 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 9861 3343 9919 3349
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 10888 3380 10916 3411
rect 10376 3352 10916 3380
rect 10376 3340 10382 3352
rect 1104 3290 13892 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 13892 3290
rect 1104 3216 13892 3238
rect 1578 3176 1584 3188
rect 1539 3148 1584 3176
rect 1578 3136 1584 3148
rect 1636 3136 1642 3188
rect 3326 3176 3332 3188
rect 2148 3148 3332 3176
rect 2148 3108 2176 3148
rect 3326 3136 3332 3148
rect 3384 3176 3390 3188
rect 3789 3179 3847 3185
rect 3384 3148 3643 3176
rect 3384 3136 3390 3148
rect 2056 3080 2176 3108
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 2056 3049 2084 3080
rect 3050 3068 3056 3120
rect 3108 3068 3114 3120
rect 3615 3108 3643 3148
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 4062 3176 4068 3188
rect 3835 3148 4068 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4614 3136 4620 3188
rect 4672 3136 4678 3188
rect 4982 3136 4988 3188
rect 5040 3176 5046 3188
rect 8021 3179 8079 3185
rect 5040 3148 7788 3176
rect 5040 3136 5046 3148
rect 4249 3111 4307 3117
rect 3615 3080 3924 3108
rect 3896 3052 3924 3080
rect 4249 3077 4261 3111
rect 4295 3108 4307 3111
rect 4632 3108 4660 3136
rect 4295 3080 4660 3108
rect 4295 3077 4307 3080
rect 4249 3071 4307 3077
rect 4890 3068 4896 3120
rect 4948 3068 4954 3120
rect 7760 3108 7788 3148
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8110 3176 8116 3188
rect 8067 3148 8116 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8220 3148 8769 3176
rect 8220 3108 8248 3148
rect 8757 3145 8769 3148
rect 8803 3176 8815 3179
rect 9122 3176 9128 3188
rect 8803 3148 9128 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9306 3176 9312 3188
rect 9267 3148 9312 3176
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 9640 3148 9996 3176
rect 9640 3136 9646 3148
rect 7760 3080 8248 3108
rect 8665 3111 8723 3117
rect 8665 3077 8677 3111
rect 8711 3108 8723 3111
rect 9858 3108 9864 3120
rect 8711 3080 9864 3108
rect 8711 3077 8723 3080
rect 8665 3071 8723 3077
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1544 3012 1777 3040
rect 1544 3000 1550 3012
rect 1765 3009 1777 3012
rect 1811 3040 1823 3043
rect 2041 3043 2099 3049
rect 2041 3040 2053 3043
rect 1811 3012 2053 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 2041 3009 2053 3012
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3936 3012 3985 3040
rect 3936 3000 3942 3012
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 3973 3003 4031 3009
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6880 3012 7021 3040
rect 6880 3000 6886 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8018 3040 8024 3052
rect 7607 3012 8024 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2972 2375 2975
rect 3786 2972 3792 2984
rect 2363 2944 3792 2972
rect 2363 2941 2375 2944
rect 2317 2935 2375 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 6917 2975 6975 2981
rect 4080 2944 5856 2972
rect 4080 2904 4108 2944
rect 5718 2904 5724 2916
rect 3712 2876 4108 2904
rect 5679 2876 5724 2904
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 3712 2836 3740 2876
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 992 2808 3740 2836
rect 5828 2836 5856 2944
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 6963 2944 7113 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 7101 2941 7113 2944
rect 7147 2941 7159 2975
rect 7101 2935 7159 2941
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 7190 2904 7196 2916
rect 6871 2876 7196 2904
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 7190 2864 7196 2876
rect 7248 2904 7254 2916
rect 7392 2904 7420 3003
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8680 3040 8708 3071
rect 9858 3068 9864 3080
rect 9916 3068 9922 3120
rect 9968 3117 9996 3148
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 12032 3148 12173 3176
rect 12032 3136 12038 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 9953 3111 10011 3117
rect 9953 3077 9965 3111
rect 9999 3077 10011 3111
rect 10134 3108 10140 3120
rect 10095 3080 10140 3108
rect 9953 3071 10011 3077
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 9030 3040 9036 3052
rect 8159 3012 8708 3040
rect 8991 3012 9036 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 10336 3049 10364 3136
rect 10686 3108 10692 3120
rect 10612 3080 10692 3108
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 9456 3012 9505 3040
rect 9456 3000 9462 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 8297 2975 8355 2981
rect 8297 2941 8309 2975
rect 8343 2972 8355 2975
rect 8386 2972 8392 2984
rect 8343 2944 8392 2972
rect 8343 2941 8355 2944
rect 8297 2935 8355 2941
rect 8386 2932 8392 2944
rect 8444 2972 8450 2984
rect 9048 2972 9076 3000
rect 9582 2972 9588 2984
rect 9640 2981 9646 2984
rect 8444 2944 9076 2972
rect 9547 2944 9588 2972
rect 8444 2932 8450 2944
rect 9582 2932 9588 2944
rect 9640 2935 9647 2981
rect 9784 2972 9812 3003
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10612 3040 10640 3080
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 10778 3040 10784 3052
rect 10468 3012 10640 3040
rect 10739 3012 10784 3040
rect 10468 3000 10474 3012
rect 10612 2981 10640 3012
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11164 3040 11192 3136
rect 12066 3108 12072 3120
rect 12027 3080 12072 3108
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11164 3012 11529 3040
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11940 3012 11989 3040
rect 11940 3000 11946 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 11977 3003 12035 3009
rect 12406 3012 12541 3040
rect 10597 2975 10655 2981
rect 9784 2944 10364 2972
rect 9640 2932 9646 2935
rect 7248 2876 7420 2904
rect 7248 2864 7254 2876
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 9677 2907 9735 2913
rect 9677 2904 9689 2907
rect 9548 2876 9689 2904
rect 9548 2864 9554 2876
rect 9677 2873 9689 2876
rect 9723 2873 9735 2907
rect 9677 2867 9735 2873
rect 7282 2836 7288 2848
rect 5828 2808 7288 2836
rect 992 2796 998 2808
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 7558 2796 7564 2848
rect 7616 2836 7622 2848
rect 7653 2839 7711 2845
rect 7653 2836 7665 2839
rect 7616 2808 7665 2836
rect 7616 2796 7622 2808
rect 7653 2805 7665 2808
rect 7699 2805 7711 2839
rect 10336 2836 10364 2944
rect 10597 2941 10609 2975
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10735 2944 11253 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 10410 2864 10416 2916
rect 10468 2904 10474 2916
rect 10704 2904 10732 2935
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 12406 2972 12434 3012
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 11480 2944 12434 2972
rect 12621 2975 12679 2981
rect 11480 2932 11486 2944
rect 12621 2941 12633 2975
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 10468 2876 10732 2904
rect 10468 2864 10474 2876
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 12636 2904 12664 2935
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13173 2975 13231 2981
rect 13173 2972 13185 2975
rect 12768 2944 13185 2972
rect 12768 2932 12774 2944
rect 13173 2941 13185 2944
rect 13219 2941 13231 2975
rect 13173 2935 13231 2941
rect 12124 2876 12434 2904
rect 12636 2876 13308 2904
rect 12124 2864 12130 2876
rect 11054 2836 11060 2848
rect 10336 2808 11060 2836
rect 7653 2799 7711 2805
rect 11054 2796 11060 2808
rect 11112 2836 11118 2848
rect 11698 2836 11704 2848
rect 11112 2808 11704 2836
rect 11112 2796 11118 2808
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 12406 2836 12434 2876
rect 12989 2839 13047 2845
rect 12989 2836 13001 2839
rect 12406 2808 13001 2836
rect 12989 2805 13001 2808
rect 13035 2805 13047 2839
rect 13280 2836 13308 2876
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 13280 2808 13461 2836
rect 12989 2799 13047 2805
rect 13449 2805 13461 2808
rect 13495 2836 13507 2839
rect 14001 2839 14059 2845
rect 14001 2836 14013 2839
rect 13495 2808 14013 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 14001 2805 14013 2808
rect 14047 2805 14059 2839
rect 14001 2799 14059 2805
rect 1104 2746 13892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 13892 2746
rect 1104 2672 13892 2694
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 4028 2604 4077 2632
rect 4028 2592 4034 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4890 2632 4896 2644
rect 4851 2604 4896 2632
rect 4065 2595 4123 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 7742 2632 7748 2644
rect 5123 2604 7748 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4614 2496 4620 2508
rect 4571 2468 4620 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3142 2428 3148 2440
rect 2915 2400 3148 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3142 2388 3148 2400
rect 3200 2428 3206 2440
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 3200 2400 3249 2428
rect 3200 2388 3206 2400
rect 3237 2397 3249 2400
rect 3283 2428 3295 2431
rect 3605 2431 3663 2437
rect 3605 2428 3617 2431
rect 3283 2400 3617 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3605 2397 3617 2400
rect 3651 2428 3663 2431
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3651 2400 3801 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 4430 2428 4436 2440
rect 4391 2400 4436 2428
rect 3789 2391 3847 2397
rect 3804 2360 3832 2391
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5092 2428 5120 2595
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2632 8450 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 8444 2604 8493 2632
rect 8444 2592 8450 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 10778 2632 10784 2644
rect 10735 2604 10784 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 7190 2564 7196 2576
rect 7151 2536 7196 2564
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 8404 2564 8432 2592
rect 10318 2564 10324 2576
rect 7484 2536 10324 2564
rect 4755 2400 5120 2428
rect 5629 2431 5687 2437
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 6362 2428 6368 2440
rect 5767 2400 6368 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 4724 2360 4752 2391
rect 3804 2332 4752 2360
rect 5644 2360 5672 2391
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7484 2437 7512 2536
rect 7742 2496 7748 2508
rect 7703 2468 7748 2496
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 9508 2505 9536 2536
rect 10318 2524 10324 2536
rect 10376 2564 10382 2576
rect 10965 2567 11023 2573
rect 10965 2564 10977 2567
rect 10376 2536 10977 2564
rect 10376 2524 10382 2536
rect 10704 2508 10732 2536
rect 10965 2533 10977 2536
rect 11011 2564 11023 2567
rect 11241 2567 11299 2573
rect 11241 2564 11253 2567
rect 11011 2536 11253 2564
rect 11011 2533 11023 2536
rect 10965 2527 11023 2533
rect 11241 2533 11253 2536
rect 11287 2564 11299 2567
rect 11425 2567 11483 2573
rect 11425 2564 11437 2567
rect 11287 2536 11437 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11425 2533 11437 2536
rect 11471 2564 11483 2567
rect 12710 2564 12716 2576
rect 11471 2536 12716 2564
rect 11471 2533 11483 2536
rect 11425 2527 11483 2533
rect 9493 2499 9551 2505
rect 9493 2465 9505 2499
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 10686 2456 10692 2508
rect 10744 2456 10750 2508
rect 11900 2505 11928 2536
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 11885 2499 11943 2505
rect 11885 2465 11897 2499
rect 11931 2465 11943 2499
rect 12066 2496 12072 2508
rect 12027 2468 12072 2496
rect 11885 2459 11943 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7650 2428 7656 2440
rect 7611 2400 7656 2428
rect 7469 2391 7527 2397
rect 7650 2388 7656 2400
rect 7708 2428 7714 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7708 2400 7849 2428
rect 7708 2388 7714 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 8168 2400 8217 2428
rect 8168 2388 8174 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9674 2428 9680 2440
rect 9355 2400 9680 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 9858 2428 9864 2440
rect 9815 2400 9864 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10594 2428 10600 2440
rect 10551 2400 10600 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 11020 2400 11621 2428
rect 11020 2388 11026 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 12161 2431 12219 2437
rect 12161 2428 12173 2431
rect 11756 2400 12173 2428
rect 11756 2388 11762 2400
rect 12161 2397 12173 2400
rect 12207 2397 12219 2431
rect 12161 2391 12219 2397
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 7742 2360 7748 2372
rect 5644 2332 7748 2360
rect 7742 2320 7748 2332
rect 7800 2360 7806 2372
rect 10226 2360 10232 2372
rect 7800 2332 8248 2360
rect 10187 2332 10232 2360
rect 7800 2320 7806 2332
rect 3970 2292 3976 2304
rect 3931 2264 3976 2292
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 6454 2292 6460 2304
rect 5491 2264 6460 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 8220 2301 8248 2332
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 10318 2320 10324 2372
rect 10376 2360 10382 2372
rect 10376 2332 10421 2360
rect 10376 2320 10382 2332
rect 12636 2304 12664 2391
rect 13262 2388 13268 2440
rect 13320 2428 13326 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 13320 2400 13461 2428
rect 13320 2388 13326 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13078 2360 13084 2372
rect 13039 2332 13084 2360
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 13170 2320 13176 2372
rect 13228 2360 13234 2372
rect 13228 2332 13273 2360
rect 13228 2320 13234 2332
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2261 8263 2295
rect 8938 2292 8944 2304
rect 8899 2264 8944 2292
rect 8205 2255 8263 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 9401 2295 9459 2301
rect 9401 2261 9413 2295
rect 9447 2292 9459 2295
rect 10870 2292 10876 2304
rect 9447 2264 10876 2292
rect 9447 2261 9459 2264
rect 9401 2255 9459 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 12529 2295 12587 2301
rect 12529 2261 12541 2295
rect 12575 2292 12587 2295
rect 12618 2292 12624 2304
rect 12575 2264 12624 2292
rect 12575 2261 12587 2264
rect 12529 2255 12587 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 1104 2202 13892 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 13892 2202
rect 1104 2128 13892 2150
rect 3145 2091 3203 2097
rect 3145 2057 3157 2091
rect 3191 2057 3203 2091
rect 3145 2051 3203 2057
rect 2222 1980 2228 2032
rect 2280 1980 2286 2032
rect 3160 2020 3188 2051
rect 4430 2048 4436 2100
rect 4488 2088 4494 2100
rect 5077 2091 5135 2097
rect 5077 2088 5089 2091
rect 4488 2060 5089 2088
rect 4488 2048 4494 2060
rect 5077 2057 5089 2060
rect 5123 2088 5135 2091
rect 5350 2088 5356 2100
rect 5123 2060 5356 2088
rect 5123 2057 5135 2060
rect 5077 2051 5135 2057
rect 5350 2048 5356 2060
rect 5408 2048 5414 2100
rect 10594 2048 10600 2100
rect 10652 2088 10658 2100
rect 10965 2091 11023 2097
rect 10965 2088 10977 2091
rect 10652 2060 10977 2088
rect 10652 2048 10658 2060
rect 10965 2057 10977 2060
rect 11011 2057 11023 2091
rect 10965 2051 11023 2057
rect 11333 2091 11391 2097
rect 11333 2057 11345 2091
rect 11379 2057 11391 2091
rect 13170 2088 13176 2100
rect 13131 2060 13176 2088
rect 11333 2051 11391 2057
rect 3605 2023 3663 2029
rect 3605 2020 3617 2023
rect 3160 1992 3617 2020
rect 3605 1989 3617 1992
rect 3651 1989 3663 2023
rect 3605 1983 3663 1989
rect 5997 2023 6055 2029
rect 5997 1989 6009 2023
rect 6043 2020 6055 2023
rect 6822 2020 6828 2032
rect 6043 1992 6828 2020
rect 6043 1989 6055 1992
rect 5997 1983 6055 1989
rect 6822 1980 6828 1992
rect 6880 1980 6886 2032
rect 7190 1980 7196 2032
rect 7248 2020 7254 2032
rect 7561 2023 7619 2029
rect 7561 2020 7573 2023
rect 7248 1992 7573 2020
rect 7248 1980 7254 1992
rect 7561 1989 7573 1992
rect 7607 1989 7619 2023
rect 7742 2020 7748 2032
rect 7703 1992 7748 2020
rect 7561 1983 7619 1989
rect 7742 1980 7748 1992
rect 7800 1980 7806 2032
rect 10505 2023 10563 2029
rect 10505 2020 10517 2023
rect 9416 1992 10517 2020
rect 1394 1952 1400 1964
rect 1355 1924 1400 1952
rect 1394 1912 1400 1924
rect 1452 1912 1458 1964
rect 4706 1912 4712 1964
rect 4764 1912 4770 1964
rect 5261 1955 5319 1961
rect 5261 1921 5273 1955
rect 5307 1952 5319 1955
rect 5810 1952 5816 1964
rect 5307 1924 5816 1952
rect 5307 1921 5319 1924
rect 5261 1915 5319 1921
rect 5810 1912 5816 1924
rect 5868 1912 5874 1964
rect 6181 1955 6239 1961
rect 6181 1921 6193 1955
rect 6227 1921 6239 1955
rect 6454 1952 6460 1964
rect 6415 1924 6460 1952
rect 6181 1915 6239 1921
rect 1673 1887 1731 1893
rect 1673 1853 1685 1887
rect 1719 1884 1731 1887
rect 3234 1884 3240 1896
rect 1719 1856 3240 1884
rect 1719 1853 1731 1856
rect 1673 1847 1731 1853
rect 3234 1844 3240 1856
rect 3292 1844 3298 1896
rect 3329 1887 3387 1893
rect 3329 1853 3341 1887
rect 3375 1884 3387 1887
rect 3694 1884 3700 1896
rect 3375 1856 3700 1884
rect 3375 1853 3387 1856
rect 3329 1847 3387 1853
rect 3694 1844 3700 1856
rect 3752 1844 3758 1896
rect 6196 1884 6224 1915
rect 6454 1912 6460 1924
rect 6512 1912 6518 1964
rect 7208 1884 7236 1980
rect 6196 1856 7236 1884
rect 7760 1816 7788 1980
rect 7926 1952 7932 1964
rect 7887 1924 7932 1952
rect 7926 1912 7932 1924
rect 7984 1912 7990 1964
rect 9416 1961 9444 1992
rect 10505 1989 10517 1992
rect 10551 2020 10563 2023
rect 10870 2020 10876 2032
rect 10551 1992 10876 2020
rect 10551 1989 10563 1992
rect 10505 1983 10563 1989
rect 10870 1980 10876 1992
rect 10928 1980 10934 2032
rect 9401 1955 9459 1961
rect 9401 1921 9413 1955
rect 9447 1921 9459 1955
rect 9401 1915 9459 1921
rect 9585 1955 9643 1961
rect 9585 1921 9597 1955
rect 9631 1952 9643 1955
rect 9858 1952 9864 1964
rect 9631 1924 9864 1952
rect 9631 1921 9643 1924
rect 9585 1915 9643 1921
rect 9858 1912 9864 1924
rect 9916 1912 9922 1964
rect 10226 1952 10232 1964
rect 10187 1924 10232 1952
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
rect 11348 1952 11376 2051
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 12710 1980 12716 2032
rect 12768 2020 12774 2032
rect 13449 2023 13507 2029
rect 13449 2020 13461 2023
rect 12768 1992 13461 2020
rect 12768 1980 12774 1992
rect 13449 1989 13461 1992
rect 13495 1989 13507 2023
rect 13449 1983 13507 1989
rect 11514 1952 11520 1964
rect 11348 1924 11520 1952
rect 11514 1912 11520 1924
rect 11572 1912 11578 1964
rect 12989 1955 13047 1961
rect 12989 1921 13001 1955
rect 13035 1952 13047 1955
rect 13354 1952 13360 1964
rect 13035 1924 13360 1952
rect 13035 1921 13047 1924
rect 12989 1915 13047 1921
rect 13354 1912 13360 1924
rect 13412 1912 13418 1964
rect 10686 1884 10692 1896
rect 10647 1856 10692 1884
rect 10686 1844 10692 1856
rect 10744 1844 10750 1896
rect 10873 1887 10931 1893
rect 10873 1853 10885 1887
rect 10919 1853 10931 1887
rect 10873 1847 10931 1853
rect 9217 1819 9275 1825
rect 9217 1816 9229 1819
rect 7760 1788 9229 1816
rect 9217 1785 9229 1788
rect 9263 1816 9275 1819
rect 9398 1816 9404 1828
rect 9263 1788 9404 1816
rect 9263 1785 9275 1788
rect 9217 1779 9275 1785
rect 9398 1776 9404 1788
rect 9456 1776 9462 1828
rect 10888 1816 10916 1847
rect 10962 1816 10968 1828
rect 10888 1788 10968 1816
rect 10962 1776 10968 1788
rect 11020 1776 11026 1828
rect 12805 1819 12863 1825
rect 12805 1785 12817 1819
rect 12851 1785 12863 1819
rect 12805 1779 12863 1785
rect 5626 1708 5632 1760
rect 5684 1748 5690 1760
rect 6086 1748 6092 1760
rect 5684 1720 6092 1748
rect 5684 1708 5690 1720
rect 6086 1708 6092 1720
rect 6144 1748 6150 1760
rect 6457 1751 6515 1757
rect 6457 1748 6469 1751
rect 6144 1720 6469 1748
rect 6144 1708 6150 1720
rect 6457 1717 6469 1720
rect 6503 1717 6515 1751
rect 6457 1711 6515 1717
rect 10870 1708 10876 1760
rect 10928 1748 10934 1760
rect 12820 1748 12848 1779
rect 10928 1720 12848 1748
rect 10928 1708 10934 1720
rect 1104 1658 13892 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 13892 1658
rect 1104 1584 13892 1606
rect 2222 1544 2228 1556
rect 2183 1516 2228 1544
rect 2222 1504 2228 1516
rect 2280 1504 2286 1556
rect 3142 1544 3148 1556
rect 3103 1516 3148 1544
rect 3142 1504 3148 1516
rect 3200 1504 3206 1556
rect 7837 1547 7895 1553
rect 7837 1513 7849 1547
rect 7883 1544 7895 1547
rect 7926 1544 7932 1556
rect 7883 1516 7932 1544
rect 7883 1513 7895 1516
rect 7837 1507 7895 1513
rect 7926 1504 7932 1516
rect 7984 1504 7990 1556
rect 9858 1544 9864 1556
rect 9819 1516 9864 1544
rect 9858 1504 9864 1516
rect 9916 1504 9922 1556
rect 10318 1504 10324 1556
rect 10376 1544 10382 1556
rect 10689 1547 10747 1553
rect 10689 1544 10701 1547
rect 10376 1516 10701 1544
rect 10376 1504 10382 1516
rect 10689 1513 10701 1516
rect 10735 1513 10747 1547
rect 10689 1507 10747 1513
rect 3160 1408 3188 1504
rect 6822 1476 6828 1488
rect 6783 1448 6828 1476
rect 6822 1436 6828 1448
rect 6880 1436 6886 1488
rect 9398 1476 9404 1488
rect 9359 1448 9404 1476
rect 9398 1436 9404 1448
rect 9456 1436 9462 1488
rect 4706 1408 4712 1420
rect 2884 1380 3188 1408
rect 4172 1380 4712 1408
rect 2884 1349 2912 1380
rect 2041 1343 2099 1349
rect 2041 1309 2053 1343
rect 2087 1340 2099 1343
rect 2409 1343 2467 1349
rect 2409 1340 2421 1343
rect 2087 1312 2421 1340
rect 2087 1309 2099 1312
rect 2041 1303 2099 1309
rect 2409 1309 2421 1312
rect 2455 1340 2467 1343
rect 2869 1343 2927 1349
rect 2869 1340 2881 1343
rect 2455 1312 2881 1340
rect 2455 1309 2467 1312
rect 2409 1303 2467 1309
rect 2869 1309 2881 1312
rect 2915 1309 2927 1343
rect 3234 1340 3240 1352
rect 2869 1303 2927 1309
rect 2976 1312 3240 1340
rect 2774 1232 2780 1284
rect 2832 1272 2838 1284
rect 2976 1272 3004 1312
rect 3234 1300 3240 1312
rect 3292 1340 3298 1352
rect 3329 1343 3387 1349
rect 3329 1340 3341 1343
rect 3292 1312 3341 1340
rect 3292 1300 3298 1312
rect 3329 1309 3341 1312
rect 3375 1309 3387 1343
rect 4172 1340 4200 1380
rect 4706 1368 4712 1380
rect 4764 1368 4770 1420
rect 5350 1408 5356 1420
rect 5311 1380 5356 1408
rect 5350 1368 5356 1380
rect 5408 1368 5414 1420
rect 5626 1408 5632 1420
rect 5587 1380 5632 1408
rect 5626 1368 5632 1380
rect 5684 1368 5690 1420
rect 7558 1408 7564 1420
rect 6886 1380 7564 1408
rect 3329 1303 3387 1309
rect 3528 1312 4200 1340
rect 3528 1272 3556 1312
rect 5810 1300 5816 1352
rect 5868 1340 5874 1352
rect 6365 1343 6423 1349
rect 6365 1340 6377 1343
rect 5868 1312 6377 1340
rect 5868 1300 5874 1312
rect 6365 1309 6377 1312
rect 6411 1340 6423 1343
rect 6886 1340 6914 1380
rect 7558 1368 7564 1380
rect 7616 1368 7622 1420
rect 8110 1368 8116 1420
rect 8168 1408 8174 1420
rect 8205 1411 8263 1417
rect 8205 1408 8217 1411
rect 8168 1380 8217 1408
rect 8168 1368 8174 1380
rect 8205 1377 8217 1380
rect 8251 1377 8263 1411
rect 8938 1408 8944 1420
rect 8899 1380 8944 1408
rect 8205 1371 8263 1377
rect 8938 1368 8944 1380
rect 8996 1368 9002 1420
rect 10505 1411 10563 1417
rect 10505 1377 10517 1411
rect 10551 1408 10563 1411
rect 10686 1408 10692 1420
rect 10551 1380 10692 1408
rect 10551 1377 10563 1380
rect 10505 1371 10563 1377
rect 10686 1368 10692 1380
rect 10744 1408 10750 1420
rect 11149 1411 11207 1417
rect 11149 1408 11161 1411
rect 10744 1380 11161 1408
rect 10744 1368 10750 1380
rect 11149 1377 11161 1380
rect 11195 1377 11207 1411
rect 11514 1408 11520 1420
rect 11475 1380 11520 1408
rect 11149 1371 11207 1377
rect 11514 1368 11520 1380
rect 11572 1368 11578 1420
rect 7190 1340 7196 1352
rect 6411 1312 6914 1340
rect 7151 1312 7196 1340
rect 6411 1309 6423 1312
rect 6365 1303 6423 1309
rect 7190 1300 7196 1312
rect 7248 1300 7254 1352
rect 7282 1300 7288 1352
rect 7340 1340 7346 1352
rect 7469 1343 7527 1349
rect 7340 1312 7385 1340
rect 7340 1300 7346 1312
rect 7469 1309 7481 1343
rect 7515 1309 7527 1343
rect 7469 1303 7527 1309
rect 2832 1244 3004 1272
rect 3068 1244 3556 1272
rect 2832 1232 2838 1244
rect 3068 1213 3096 1244
rect 3970 1232 3976 1284
rect 4028 1272 4034 1284
rect 6917 1275 6975 1281
rect 4028 1244 4186 1272
rect 4028 1232 4034 1244
rect 6917 1241 6929 1275
rect 6963 1241 6975 1275
rect 6917 1235 6975 1241
rect 3053 1207 3111 1213
rect 3053 1173 3065 1207
rect 3099 1173 3111 1207
rect 3053 1167 3111 1173
rect 3881 1207 3939 1213
rect 3881 1173 3893 1207
rect 3927 1204 3939 1207
rect 4614 1204 4620 1216
rect 3927 1176 4620 1204
rect 3927 1173 3939 1176
rect 3881 1167 3939 1173
rect 4614 1164 4620 1176
rect 4672 1164 4678 1216
rect 6932 1204 6960 1235
rect 7009 1207 7067 1213
rect 7009 1204 7021 1207
rect 6932 1176 7021 1204
rect 7009 1173 7021 1176
rect 7055 1173 7067 1207
rect 7484 1204 7512 1303
rect 7650 1300 7656 1352
rect 7708 1340 7714 1352
rect 7929 1343 7987 1349
rect 7929 1340 7941 1343
rect 7708 1312 7941 1340
rect 7708 1300 7714 1312
rect 7929 1309 7941 1312
rect 7975 1309 7987 1343
rect 8665 1343 8723 1349
rect 8665 1340 8677 1343
rect 7929 1303 7987 1309
rect 8036 1312 8677 1340
rect 7558 1232 7564 1284
rect 7616 1272 7622 1284
rect 8036 1272 8064 1312
rect 8665 1309 8677 1312
rect 8711 1309 8723 1343
rect 8665 1303 8723 1309
rect 7616 1244 8064 1272
rect 8113 1275 8171 1281
rect 7616 1232 7622 1244
rect 8113 1241 8125 1275
rect 8159 1272 8171 1275
rect 8956 1272 8984 1368
rect 9769 1343 9827 1349
rect 9769 1309 9781 1343
rect 9815 1340 9827 1343
rect 10226 1340 10232 1352
rect 9815 1312 10232 1340
rect 9815 1309 9827 1312
rect 9769 1303 9827 1309
rect 10226 1300 10232 1312
rect 10284 1300 10290 1352
rect 10870 1340 10876 1352
rect 10831 1312 10876 1340
rect 10870 1300 10876 1312
rect 10928 1340 10934 1352
rect 11977 1343 12035 1349
rect 11977 1340 11989 1343
rect 10928 1312 11989 1340
rect 10928 1300 10934 1312
rect 11977 1309 11989 1312
rect 12023 1309 12035 1343
rect 11977 1303 12035 1309
rect 12437 1343 12495 1349
rect 12437 1309 12449 1343
rect 12483 1340 12495 1343
rect 12618 1340 12624 1352
rect 12483 1312 12624 1340
rect 12483 1309 12495 1312
rect 12437 1303 12495 1309
rect 12618 1300 12624 1312
rect 12676 1300 12682 1352
rect 13078 1340 13084 1352
rect 13039 1312 13084 1340
rect 13078 1300 13084 1312
rect 13136 1300 13142 1352
rect 13354 1340 13360 1352
rect 13315 1312 13360 1340
rect 13354 1300 13360 1312
rect 13412 1300 13418 1352
rect 8159 1244 8984 1272
rect 9493 1275 9551 1281
rect 8159 1241 8171 1244
rect 8113 1235 8171 1241
rect 9493 1241 9505 1275
rect 9539 1272 9551 1275
rect 9585 1275 9643 1281
rect 9585 1272 9597 1275
rect 9539 1244 9597 1272
rect 9539 1241 9551 1244
rect 9493 1235 9551 1241
rect 9585 1241 9597 1244
rect 9631 1241 9643 1275
rect 9585 1235 9643 1241
rect 10321 1275 10379 1281
rect 10321 1241 10333 1275
rect 10367 1272 10379 1275
rect 11057 1275 11115 1281
rect 11057 1272 11069 1275
rect 10367 1244 11069 1272
rect 10367 1241 10379 1244
rect 10321 1235 10379 1241
rect 11057 1241 11069 1244
rect 11103 1272 11115 1275
rect 12069 1275 12127 1281
rect 11103 1244 11836 1272
rect 11103 1241 11115 1244
rect 11057 1235 11115 1241
rect 8573 1207 8631 1213
rect 8573 1204 8585 1207
rect 7484 1176 8585 1204
rect 7009 1167 7067 1173
rect 8573 1173 8585 1176
rect 8619 1204 8631 1207
rect 9674 1204 9680 1216
rect 8619 1176 9680 1204
rect 8619 1173 8631 1176
rect 8573 1167 8631 1173
rect 9674 1164 9680 1176
rect 9732 1164 9738 1216
rect 10042 1164 10048 1216
rect 10100 1204 10106 1216
rect 10229 1207 10287 1213
rect 10229 1204 10241 1207
rect 10100 1176 10241 1204
rect 10100 1164 10106 1176
rect 10229 1173 10241 1176
rect 10275 1173 10287 1207
rect 11808 1204 11836 1244
rect 12069 1241 12081 1275
rect 12115 1272 12127 1275
rect 12161 1275 12219 1281
rect 12161 1272 12173 1275
rect 12115 1244 12173 1272
rect 12115 1241 12127 1244
rect 12069 1235 12127 1241
rect 12161 1241 12173 1244
rect 12207 1241 12219 1275
rect 12161 1235 12219 1241
rect 12345 1275 12403 1281
rect 12345 1241 12357 1275
rect 12391 1272 12403 1275
rect 13096 1272 13124 1300
rect 12391 1244 13124 1272
rect 12391 1241 12403 1244
rect 12345 1235 12403 1241
rect 13998 1204 14004 1216
rect 11808 1176 14004 1204
rect 10229 1167 10287 1173
rect 13998 1164 14004 1176
rect 14056 1164 14062 1216
rect 1104 1114 13892 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 13892 1114
rect 1104 1040 13892 1062
rect 9674 960 9680 1012
rect 9732 1000 9738 1012
rect 10778 1000 10784 1012
rect 9732 972 10784 1000
rect 9732 960 9738 972
rect 10778 960 10784 972
rect 10836 960 10842 1012
rect 13906 484 13912 536
rect 13964 524 13970 536
rect 14001 527 14059 533
rect 14001 524 14013 527
rect 13964 496 14013 524
rect 13964 484 13970 496
rect 14001 493 14013 496
rect 14047 493 14059 527
rect 14001 487 14059 493
<< via1 >>
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 3424 13268 3476 13320
rect 5540 13472 5592 13524
rect 6920 13447 6972 13456
rect 6920 13413 6929 13447
rect 6929 13413 6963 13447
rect 6963 13413 6972 13447
rect 6920 13404 6972 13413
rect 8208 13472 8260 13524
rect 9772 13404 9824 13456
rect 5908 13336 5960 13388
rect 6000 13268 6052 13320
rect 6828 13336 6880 13388
rect 5172 13200 5224 13252
rect 6552 13243 6604 13252
rect 6552 13209 6561 13243
rect 6561 13209 6595 13243
rect 6595 13209 6604 13243
rect 6552 13200 6604 13209
rect 6828 13200 6880 13252
rect 3332 13175 3384 13184
rect 3332 13141 3341 13175
rect 3341 13141 3375 13175
rect 3375 13141 3384 13175
rect 3332 13132 3384 13141
rect 5356 13175 5408 13184
rect 5356 13141 5365 13175
rect 5365 13141 5399 13175
rect 5399 13141 5408 13175
rect 5356 13132 5408 13141
rect 7932 13268 7984 13320
rect 7012 13132 7064 13184
rect 7564 13132 7616 13184
rect 8576 13132 8628 13184
rect 9496 13132 9548 13184
rect 11336 13268 11388 13320
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 12532 13243 12584 13252
rect 12532 13209 12541 13243
rect 12541 13209 12575 13243
rect 12575 13209 12584 13243
rect 12532 13200 12584 13209
rect 12624 13243 12676 13252
rect 12624 13209 12633 13243
rect 12633 13209 12667 13243
rect 12667 13209 12676 13243
rect 13176 13243 13228 13252
rect 12624 13200 12676 13209
rect 13176 13209 13185 13243
rect 13185 13209 13219 13243
rect 13219 13209 13228 13243
rect 13176 13200 13228 13209
rect 13360 13200 13412 13252
rect 10048 13175 10100 13184
rect 10048 13141 10057 13175
rect 10057 13141 10091 13175
rect 10091 13141 10100 13175
rect 10048 13132 10100 13141
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 2504 12928 2556 12980
rect 3332 12860 3384 12912
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 4712 12928 4764 12980
rect 6000 12971 6052 12980
rect 5540 12860 5592 12912
rect 6000 12937 6009 12971
rect 6009 12937 6043 12971
rect 6043 12937 6052 12971
rect 6000 12928 6052 12937
rect 6828 12928 6880 12980
rect 7932 12928 7984 12980
rect 6552 12860 6604 12912
rect 6920 12860 6972 12912
rect 8116 12792 8168 12844
rect 11336 12903 11388 12912
rect 11336 12869 11345 12903
rect 11345 12869 11379 12903
rect 11379 12869 11388 12903
rect 11336 12860 11388 12869
rect 8576 12792 8628 12844
rect 9128 12792 9180 12844
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 11244 12835 11296 12844
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 12072 12928 12124 12980
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 4620 12724 4672 12776
rect 10048 12724 10100 12776
rect 8392 12656 8444 12708
rect 9220 12656 9272 12708
rect 12532 12656 12584 12708
rect 12992 12699 13044 12708
rect 12992 12665 13001 12699
rect 13001 12665 13035 12699
rect 13035 12665 13044 12699
rect 12992 12656 13044 12665
rect 10048 12588 10100 12640
rect 10876 12588 10928 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 4620 12427 4672 12436
rect 4620 12393 4629 12427
rect 4629 12393 4663 12427
rect 4663 12393 4672 12427
rect 4620 12384 4672 12393
rect 5908 12384 5960 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 10876 12384 10928 12436
rect 12624 12384 12676 12436
rect 3516 12316 3568 12368
rect 2964 12180 3016 12232
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 2688 12112 2740 12164
rect 4620 12180 4672 12232
rect 9312 12316 9364 12368
rect 5356 12291 5408 12300
rect 5356 12257 5365 12291
rect 5365 12257 5399 12291
rect 5399 12257 5408 12291
rect 5356 12248 5408 12257
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 1400 12044 1452 12096
rect 2504 12044 2556 12096
rect 3148 12087 3200 12096
rect 3148 12053 3157 12087
rect 3157 12053 3191 12087
rect 3191 12053 3200 12087
rect 3148 12044 3200 12053
rect 3884 12044 3936 12096
rect 5080 12112 5132 12164
rect 5540 12180 5592 12232
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 7196 12180 7248 12232
rect 8392 12223 8444 12232
rect 6736 12112 6788 12164
rect 8392 12189 8400 12223
rect 8400 12189 8434 12223
rect 8434 12189 8444 12223
rect 8392 12180 8444 12189
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 9220 12223 9272 12232
rect 6000 12044 6052 12096
rect 8668 12112 8720 12164
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 8760 12044 8812 12096
rect 11336 12248 11388 12300
rect 10324 12223 10376 12232
rect 9404 12112 9456 12164
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 12716 12316 12768 12368
rect 13176 12248 13228 12300
rect 9680 12112 9732 12164
rect 10140 12112 10192 12164
rect 12900 12112 12952 12164
rect 9956 12087 10008 12096
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 11152 12044 11204 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 2688 11840 2740 11892
rect 3884 11772 3936 11824
rect 5080 11840 5132 11892
rect 6736 11883 6788 11892
rect 2872 11704 2924 11756
rect 1492 11679 1544 11688
rect 1492 11645 1501 11679
rect 1501 11645 1535 11679
rect 1535 11645 1544 11679
rect 1492 11636 1544 11645
rect 2504 11636 2556 11688
rect 3792 11636 3844 11688
rect 5540 11704 5592 11756
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 6736 11849 6745 11883
rect 6745 11849 6779 11883
rect 6779 11849 6788 11883
rect 6736 11840 6788 11849
rect 8576 11840 8628 11892
rect 9772 11840 9824 11892
rect 11244 11840 11296 11892
rect 6552 11704 6604 11756
rect 6736 11636 6788 11688
rect 7196 11704 7248 11756
rect 8760 11704 8812 11756
rect 9312 11815 9364 11824
rect 9312 11781 9321 11815
rect 9321 11781 9355 11815
rect 9355 11781 9364 11815
rect 9312 11772 9364 11781
rect 7380 11636 7432 11688
rect 8024 11636 8076 11688
rect 8668 11636 8720 11688
rect 9680 11636 9732 11688
rect 10048 11772 10100 11824
rect 11152 11815 11204 11824
rect 11152 11781 11161 11815
rect 11161 11781 11195 11815
rect 11195 11781 11204 11815
rect 11152 11772 11204 11781
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10876 11704 10928 11756
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 11244 11704 11296 11756
rect 12992 11772 13044 11824
rect 10048 11636 10100 11645
rect 10324 11636 10376 11688
rect 11336 11636 11388 11688
rect 11888 11636 11940 11688
rect 12900 11679 12952 11688
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 12900 11636 12952 11645
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 5080 11500 5132 11552
rect 5264 11500 5316 11552
rect 5356 11500 5408 11552
rect 6828 11500 6880 11552
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 9128 11568 9180 11620
rect 12992 11568 13044 11620
rect 9312 11500 9364 11552
rect 10232 11500 10284 11552
rect 10876 11500 10928 11552
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 2596 11228 2648 11280
rect 4620 11296 4672 11348
rect 3792 11271 3844 11280
rect 3792 11237 3801 11271
rect 3801 11237 3835 11271
rect 3835 11237 3844 11271
rect 3792 11228 3844 11237
rect 3884 11228 3936 11280
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 7196 11296 7248 11348
rect 4804 11160 4856 11212
rect 6920 11228 6972 11280
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 11244 11228 11296 11280
rect 12992 11228 13044 11280
rect 8668 11160 8720 11212
rect 9312 11203 9364 11212
rect 3240 11092 3292 11144
rect 3516 11092 3568 11144
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 3976 11092 4028 11144
rect 3884 11024 3936 11076
rect 4160 11095 4168 11122
rect 4168 11095 4202 11122
rect 4202 11095 4212 11122
rect 4160 11070 4212 11095
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 4896 11067 4948 11076
rect 4896 11033 4923 11067
rect 4923 11033 4948 11067
rect 5080 11067 5132 11076
rect 4896 11024 4948 11033
rect 5080 11033 5089 11067
rect 5089 11033 5123 11067
rect 5123 11033 5132 11067
rect 5080 11024 5132 11033
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 6092 11135 6144 11144
rect 5908 11092 5960 11101
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 6828 11092 6880 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7104 11024 7156 11076
rect 7380 11092 7432 11144
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 9312 11160 9364 11169
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 9404 11092 9456 11144
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 9312 11024 9364 11076
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 3148 10999 3200 11008
rect 3148 10965 3157 10999
rect 3157 10965 3191 10999
rect 3191 10965 3200 10999
rect 3148 10956 3200 10965
rect 3976 10956 4028 11008
rect 4160 10956 4212 11008
rect 5540 10956 5592 11008
rect 5724 10956 5776 11008
rect 6460 10956 6512 11008
rect 8116 10956 8168 11008
rect 9404 10956 9456 11008
rect 9588 10999 9640 11008
rect 9588 10965 9597 10999
rect 9597 10965 9631 10999
rect 9631 10965 9640 10999
rect 9588 10956 9640 10965
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 4896 10752 4948 10804
rect 9220 10752 9272 10804
rect 9404 10752 9456 10804
rect 9680 10752 9732 10804
rect 9864 10752 9916 10804
rect 2320 10684 2372 10736
rect 3608 10684 3660 10736
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 4804 10684 4856 10736
rect 5632 10727 5684 10736
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 5632 10693 5641 10727
rect 5641 10693 5675 10727
rect 5675 10693 5684 10727
rect 5632 10684 5684 10693
rect 6092 10684 6144 10736
rect 6552 10684 6604 10736
rect 7196 10727 7248 10736
rect 4160 10616 4212 10625
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 3792 10548 3844 10557
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 5540 10616 5592 10668
rect 6644 10616 6696 10668
rect 7196 10693 7205 10727
rect 7205 10693 7239 10727
rect 7239 10693 7248 10727
rect 7196 10684 7248 10693
rect 7288 10616 7340 10668
rect 6828 10591 6880 10600
rect 4620 10548 4672 10557
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 10140 10752 10192 10804
rect 11888 10752 11940 10804
rect 12900 10752 12952 10804
rect 11244 10727 11296 10736
rect 8116 10659 8168 10668
rect 8116 10625 8125 10659
rect 8125 10625 8159 10659
rect 8159 10625 8168 10659
rect 8116 10616 8168 10625
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 8668 10616 8720 10668
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 10232 10616 10284 10668
rect 11244 10693 11253 10727
rect 11253 10693 11287 10727
rect 11287 10693 11296 10727
rect 11244 10684 11296 10693
rect 13084 10684 13136 10736
rect 13268 10684 13320 10736
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 12624 10616 12676 10668
rect 7104 10548 7156 10557
rect 8852 10591 8904 10600
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 5264 10480 5316 10532
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 9956 10548 10008 10600
rect 9404 10480 9456 10532
rect 4712 10412 4764 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5356 10412 5408 10464
rect 5724 10412 5776 10464
rect 8668 10412 8720 10464
rect 10416 10412 10468 10464
rect 11704 10455 11756 10464
rect 11704 10421 11713 10455
rect 11713 10421 11747 10455
rect 11747 10421 11756 10455
rect 11704 10412 11756 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 1676 10208 1728 10260
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2872 10208 2924 10260
rect 4620 10208 4672 10260
rect 3424 10072 3476 10124
rect 2872 10004 2924 10056
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 4344 10140 4396 10192
rect 5356 10208 5408 10260
rect 5448 10208 5500 10260
rect 6920 10251 6972 10260
rect 6368 10183 6420 10192
rect 6368 10149 6377 10183
rect 6377 10149 6411 10183
rect 6411 10149 6420 10183
rect 6368 10140 6420 10149
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 7104 10208 7156 10260
rect 8116 10208 8168 10260
rect 8576 10208 8628 10260
rect 10048 10208 10100 10260
rect 8944 10140 8996 10192
rect 9956 10140 10008 10192
rect 10876 10208 10928 10260
rect 10416 10183 10468 10192
rect 10416 10149 10425 10183
rect 10425 10149 10459 10183
rect 10459 10149 10468 10183
rect 10416 10140 10468 10149
rect 11796 10183 11848 10192
rect 4620 10072 4672 10124
rect 2228 9936 2280 9988
rect 2964 9936 3016 9988
rect 3148 9936 3200 9988
rect 3700 10004 3752 10056
rect 4712 10047 4764 10056
rect 3792 9936 3844 9988
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5632 10072 5684 10124
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 6000 10072 6052 10124
rect 7196 10115 7248 10124
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 7196 10081 7205 10115
rect 7205 10081 7239 10115
rect 7239 10081 7248 10115
rect 7196 10072 7248 10081
rect 5816 10004 5868 10013
rect 5632 9979 5684 9988
rect 5632 9945 5641 9979
rect 5641 9945 5675 9979
rect 5675 9945 5684 9979
rect 5632 9936 5684 9945
rect 6920 10004 6972 10056
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 8576 10072 8628 10124
rect 8116 10004 8168 10056
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 8668 9936 8720 9988
rect 6276 9868 6328 9920
rect 6828 9868 6880 9920
rect 8576 9868 8628 9920
rect 11152 10004 11204 10056
rect 11796 10149 11805 10183
rect 11805 10149 11839 10183
rect 11839 10149 11848 10183
rect 11796 10140 11848 10149
rect 13084 10183 13136 10192
rect 13084 10149 13093 10183
rect 13093 10149 13127 10183
rect 13127 10149 13136 10183
rect 13084 10140 13136 10149
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 12624 10047 12676 10056
rect 11060 9936 11112 9988
rect 11520 9936 11572 9988
rect 11152 9868 11204 9920
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 13268 10004 13320 10056
rect 14188 9868 14240 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 2964 9664 3016 9716
rect 6552 9664 6604 9716
rect 6920 9664 6972 9716
rect 8852 9707 8904 9716
rect 8852 9673 8861 9707
rect 8861 9673 8895 9707
rect 8895 9673 8904 9707
rect 8852 9664 8904 9673
rect 2228 9596 2280 9648
rect 3792 9639 3844 9648
rect 3792 9605 3801 9639
rect 3801 9605 3835 9639
rect 3835 9605 3844 9639
rect 3792 9596 3844 9605
rect 3608 9571 3660 9580
rect 3608 9537 3612 9571
rect 3612 9537 3646 9571
rect 3646 9537 3660 9571
rect 3608 9528 3660 9537
rect 5540 9596 5592 9648
rect 5816 9596 5868 9648
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 3332 9460 3384 9512
rect 4712 9571 4764 9580
rect 3792 9460 3844 9512
rect 3884 9460 3936 9512
rect 4344 9503 4396 9512
rect 4344 9469 4353 9503
rect 4353 9469 4387 9503
rect 4387 9469 4396 9503
rect 4344 9460 4396 9469
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 4804 9460 4856 9512
rect 3608 9392 3660 9444
rect 5908 9528 5960 9580
rect 6368 9596 6420 9648
rect 8944 9596 8996 9648
rect 10324 9596 10376 9648
rect 11060 9639 11112 9648
rect 11060 9605 11069 9639
rect 11069 9605 11103 9639
rect 11103 9605 11112 9639
rect 11060 9596 11112 9605
rect 12992 9596 13044 9648
rect 8300 9571 8352 9580
rect 5540 9460 5592 9512
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 8576 9528 8628 9580
rect 9680 9528 9732 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 11244 9528 11296 9580
rect 12072 9528 12124 9580
rect 5448 9392 5500 9444
rect 2780 9324 2832 9376
rect 5172 9324 5224 9376
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 6828 9324 6880 9376
rect 8852 9460 8904 9512
rect 10508 9460 10560 9512
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 10876 9392 10928 9444
rect 11980 9392 12032 9444
rect 13084 9367 13136 9376
rect 13084 9333 13093 9367
rect 13093 9333 13127 9367
rect 13127 9333 13136 9367
rect 13084 9324 13136 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 4620 9120 4672 9172
rect 4988 9120 5040 9172
rect 2872 9052 2924 9104
rect 3424 9052 3476 9104
rect 1860 8916 1912 8968
rect 3332 8916 3384 8968
rect 5172 9027 5224 9036
rect 5172 8993 5181 9027
rect 5181 8993 5215 9027
rect 5215 8993 5224 9027
rect 5172 8984 5224 8993
rect 7196 9120 7248 9172
rect 8852 9120 8904 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 10324 9095 10376 9104
rect 10324 9061 10333 9095
rect 10333 9061 10367 9095
rect 10367 9061 10376 9095
rect 10324 9052 10376 9061
rect 12532 9052 12584 9104
rect 13084 8984 13136 9036
rect 7012 8916 7064 8968
rect 11244 8916 11296 8968
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 13268 8916 13320 8968
rect 5448 8848 5500 8900
rect 6184 8848 6236 8900
rect 7932 8891 7984 8900
rect 7932 8857 7941 8891
rect 7941 8857 7975 8891
rect 7975 8857 7984 8891
rect 7932 8848 7984 8857
rect 8024 8891 8076 8900
rect 8024 8857 8033 8891
rect 8033 8857 8067 8891
rect 8067 8857 8076 8891
rect 8024 8848 8076 8857
rect 12072 8848 12124 8900
rect 3332 8780 3384 8832
rect 3792 8780 3844 8832
rect 3884 8780 3936 8832
rect 4160 8780 4212 8832
rect 9404 8780 9456 8832
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 13084 8780 13136 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 3332 8576 3384 8628
rect 3424 8576 3476 8628
rect 2872 8508 2924 8560
rect 3056 8508 3108 8560
rect 3884 8508 3936 8560
rect 4896 8576 4948 8628
rect 5908 8576 5960 8628
rect 6184 8576 6236 8628
rect 7932 8576 7984 8628
rect 5816 8508 5868 8560
rect 10140 8576 10192 8628
rect 11520 8619 11572 8628
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 2780 8440 2832 8492
rect 4712 8440 4764 8492
rect 9036 8551 9088 8560
rect 9036 8517 9045 8551
rect 9045 8517 9079 8551
rect 9079 8517 9088 8551
rect 9036 8508 9088 8517
rect 10508 8551 10560 8560
rect 10508 8517 10517 8551
rect 10517 8517 10551 8551
rect 10551 8517 10560 8551
rect 10508 8508 10560 8517
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 12624 8576 12676 8628
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 10416 8440 10468 8492
rect 11428 8508 11480 8560
rect 12532 8551 12584 8560
rect 12532 8517 12541 8551
rect 12541 8517 12575 8551
rect 12575 8517 12584 8551
rect 12532 8508 12584 8517
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 1952 8304 2004 8356
rect 11980 8372 12032 8424
rect 12900 8304 12952 8356
rect 2688 8279 2740 8288
rect 2688 8245 2697 8279
rect 2697 8245 2731 8279
rect 2731 8245 2740 8279
rect 2688 8236 2740 8245
rect 2964 8236 3016 8288
rect 7748 8236 7800 8288
rect 9036 8236 9088 8288
rect 10784 8236 10836 8288
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 13176 8236 13228 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 2412 8032 2464 8084
rect 6552 8032 6604 8084
rect 1400 7896 1452 7948
rect 2964 7896 3016 7948
rect 4620 7896 4672 7948
rect 6184 7896 6236 7948
rect 7012 8032 7064 8084
rect 9036 8032 9088 8084
rect 8024 7964 8076 8016
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 1952 7760 2004 7812
rect 2688 7760 2740 7812
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 3976 7692 4028 7744
rect 5448 7760 5500 7812
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 8024 7828 8076 7880
rect 8576 7896 8628 7948
rect 8852 7828 8904 7880
rect 9036 7828 9088 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 9956 7828 10008 7880
rect 10048 7828 10100 7880
rect 9588 7760 9640 7812
rect 10876 8032 10928 8084
rect 11980 8032 12032 8084
rect 13176 8032 13228 8084
rect 11888 7964 11940 8016
rect 12624 7964 12676 8016
rect 10784 7896 10836 7948
rect 11520 7896 11572 7948
rect 13084 7896 13136 7948
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11980 7828 12032 7880
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 7932 7692 7984 7744
rect 10140 7735 10192 7744
rect 10140 7701 10149 7735
rect 10149 7701 10183 7735
rect 10183 7701 10192 7735
rect 10140 7692 10192 7701
rect 10968 7692 11020 7744
rect 12716 7692 12768 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 2964 7488 3016 7540
rect 2228 7420 2280 7472
rect 3884 7420 3936 7472
rect 3056 7352 3108 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 2320 7284 2372 7336
rect 2412 7284 2464 7336
rect 3700 7395 3752 7404
rect 3700 7361 3714 7395
rect 3714 7361 3748 7395
rect 3748 7361 3752 7395
rect 3700 7352 3752 7361
rect 4620 7395 4672 7404
rect 3792 7284 3844 7336
rect 3976 7216 4028 7268
rect 4620 7361 4628 7395
rect 4628 7361 4662 7395
rect 4662 7361 4672 7395
rect 4620 7352 4672 7361
rect 8668 7488 8720 7540
rect 9496 7488 9548 7540
rect 5724 7420 5776 7472
rect 5816 7420 5868 7472
rect 5172 7352 5224 7404
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 7012 7420 7064 7472
rect 7840 7463 7892 7472
rect 7840 7429 7849 7463
rect 7849 7429 7883 7463
rect 7883 7429 7892 7463
rect 7840 7420 7892 7429
rect 8024 7420 8076 7472
rect 4712 7327 4764 7336
rect 4712 7293 4721 7327
rect 4721 7293 4755 7327
rect 4755 7293 4764 7327
rect 4712 7284 4764 7293
rect 4620 7216 4672 7268
rect 5632 7284 5684 7336
rect 7472 7352 7524 7404
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 7380 7284 7432 7336
rect 7932 7284 7984 7336
rect 8852 7352 8904 7404
rect 9036 7420 9088 7472
rect 10140 7488 10192 7540
rect 10968 7531 11020 7540
rect 10968 7497 10977 7531
rect 10977 7497 11011 7531
rect 11011 7497 11020 7531
rect 10968 7488 11020 7497
rect 11152 7488 11204 7540
rect 11980 7488 12032 7540
rect 9404 7352 9456 7404
rect 9772 7352 9824 7404
rect 9956 7352 10008 7404
rect 8024 7216 8076 7268
rect 2780 7148 2832 7200
rect 3424 7148 3476 7200
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 6092 7148 6144 7157
rect 6460 7148 6512 7200
rect 8576 7148 8628 7200
rect 9220 7284 9272 7336
rect 11152 7352 11204 7404
rect 12808 7352 12860 7404
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 10968 7284 11020 7336
rect 11980 7284 12032 7336
rect 10140 7216 10192 7268
rect 13268 7216 13320 7268
rect 9036 7148 9088 7200
rect 11980 7191 12032 7200
rect 11980 7157 11989 7191
rect 11989 7157 12023 7191
rect 12023 7157 12032 7191
rect 11980 7148 12032 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 2228 6987 2280 6996
rect 2228 6953 2237 6987
rect 2237 6953 2271 6987
rect 2271 6953 2280 6987
rect 2228 6944 2280 6953
rect 2872 6944 2924 6996
rect 4620 6944 4672 6996
rect 5816 6944 5868 6996
rect 9312 6944 9364 6996
rect 2320 6919 2372 6928
rect 2320 6885 2329 6919
rect 2329 6885 2363 6919
rect 2363 6885 2372 6919
rect 2320 6876 2372 6885
rect 3332 6876 3384 6928
rect 3608 6876 3660 6928
rect 3792 6919 3844 6928
rect 3792 6885 3801 6919
rect 3801 6885 3835 6919
rect 3835 6885 3844 6919
rect 3792 6876 3844 6885
rect 4988 6919 5040 6928
rect 4988 6885 4997 6919
rect 4997 6885 5031 6919
rect 5031 6885 5040 6919
rect 4988 6876 5040 6885
rect 7840 6919 7892 6928
rect 7840 6885 7849 6919
rect 7849 6885 7883 6919
rect 7883 6885 7892 6919
rect 7840 6876 7892 6885
rect 2964 6740 3016 6792
rect 3148 6740 3200 6792
rect 3792 6740 3844 6792
rect 3884 6740 3936 6792
rect 4436 6808 4488 6860
rect 5172 6808 5224 6860
rect 8760 6876 8812 6928
rect 9036 6876 9088 6928
rect 9772 6876 9824 6928
rect 9128 6808 9180 6860
rect 5080 6783 5132 6792
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 4712 6672 4764 6724
rect 2780 6604 2832 6613
rect 3700 6604 3752 6656
rect 3884 6604 3936 6656
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5264 6740 5316 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 7472 6740 7524 6792
rect 10048 6944 10100 6996
rect 11060 6944 11112 6996
rect 9956 6808 10008 6860
rect 10232 6808 10284 6860
rect 11888 6808 11940 6860
rect 5724 6672 5776 6724
rect 6460 6672 6512 6724
rect 7840 6672 7892 6724
rect 11152 6740 11204 6792
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 4896 6604 4948 6656
rect 7380 6604 7432 6656
rect 10048 6672 10100 6724
rect 9036 6604 9088 6656
rect 10324 6604 10376 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 11336 6672 11388 6724
rect 13360 6672 13412 6724
rect 10600 6604 10652 6613
rect 11428 6647 11480 6656
rect 11428 6613 11437 6647
rect 11437 6613 11471 6647
rect 11471 6613 11480 6647
rect 11428 6604 11480 6613
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 2320 6332 2372 6384
rect 3976 6400 4028 6452
rect 3792 6332 3844 6384
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4712 6264 4764 6316
rect 4804 6196 4856 6248
rect 4436 6128 4488 6180
rect 4620 6128 4672 6180
rect 5632 6400 5684 6452
rect 5908 6400 5960 6452
rect 6000 6400 6052 6452
rect 6092 6332 6144 6384
rect 5816 6264 5868 6316
rect 5908 6264 5960 6316
rect 8024 6400 8076 6452
rect 8944 6400 8996 6452
rect 9036 6400 9088 6452
rect 10232 6400 10284 6452
rect 6644 6264 6696 6316
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7380 6264 7432 6316
rect 7012 6239 7064 6248
rect 7012 6205 7021 6239
rect 7021 6205 7055 6239
rect 7055 6205 7064 6239
rect 8024 6264 8076 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 9404 6264 9456 6316
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10600 6400 10652 6452
rect 11520 6400 11572 6452
rect 10784 6375 10836 6384
rect 10784 6341 10793 6375
rect 10793 6341 10827 6375
rect 10827 6341 10836 6375
rect 10784 6332 10836 6341
rect 10876 6332 10928 6384
rect 11888 6332 11940 6384
rect 12900 6332 12952 6384
rect 13360 6375 13412 6384
rect 13360 6341 13369 6375
rect 13369 6341 13403 6375
rect 13403 6341 13412 6375
rect 13360 6332 13412 6341
rect 9036 6239 9088 6248
rect 7012 6196 7064 6205
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 3884 6060 3936 6112
rect 6000 6128 6052 6180
rect 6460 6128 6512 6180
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 5356 6060 5408 6112
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 6920 6060 6972 6112
rect 10508 6128 10560 6180
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 7840 6060 7892 6112
rect 8576 6060 8628 6112
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 9220 6060 9272 6112
rect 9404 6060 9456 6112
rect 10232 6060 10284 6112
rect 11704 6264 11756 6316
rect 12072 6264 12124 6316
rect 11980 6196 12032 6248
rect 12808 6196 12860 6248
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 3608 5856 3660 5908
rect 4712 5856 4764 5908
rect 4988 5856 5040 5908
rect 5632 5856 5684 5908
rect 1768 5652 1820 5704
rect 2780 5788 2832 5840
rect 4068 5788 4120 5840
rect 3884 5763 3936 5772
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 3884 5729 3893 5763
rect 3893 5729 3927 5763
rect 3927 5729 3936 5763
rect 3884 5720 3936 5729
rect 4896 5788 4948 5840
rect 7012 5856 7064 5908
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 7564 5856 7616 5908
rect 9496 5899 9548 5908
rect 5816 5788 5868 5840
rect 6460 5788 6512 5840
rect 6920 5831 6972 5840
rect 6920 5797 6929 5831
rect 6929 5797 6963 5831
rect 6963 5797 6972 5831
rect 6920 5788 6972 5797
rect 3148 5652 3200 5704
rect 5724 5720 5776 5772
rect 6000 5720 6052 5772
rect 7656 5788 7708 5840
rect 8944 5788 8996 5840
rect 7748 5720 7800 5772
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 12808 5899 12860 5908
rect 10048 5788 10100 5840
rect 10232 5788 10284 5840
rect 10600 5788 10652 5840
rect 10784 5788 10836 5840
rect 4620 5584 4672 5636
rect 1768 5516 1820 5568
rect 3332 5516 3384 5568
rect 5264 5516 5316 5568
rect 6184 5695 6236 5704
rect 5816 5627 5868 5636
rect 5816 5593 5825 5627
rect 5825 5593 5859 5627
rect 5859 5593 5868 5627
rect 5816 5584 5868 5593
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 6276 5652 6328 5704
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 6920 5584 6972 5636
rect 7012 5584 7064 5636
rect 8668 5652 8720 5704
rect 8852 5652 8904 5704
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 10232 5652 10284 5704
rect 10416 5652 10468 5704
rect 11060 5652 11112 5704
rect 12072 5788 12124 5840
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 13176 5788 13228 5840
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 8116 5516 8168 5568
rect 9036 5516 9088 5568
rect 9956 5516 10008 5568
rect 12900 5652 12952 5704
rect 13176 5627 13228 5636
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 10876 5559 10928 5568
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 13176 5593 13185 5627
rect 13185 5593 13219 5627
rect 13219 5593 13228 5627
rect 13176 5584 13228 5593
rect 10876 5516 10928 5525
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 2872 5312 2924 5364
rect 4712 5312 4764 5364
rect 5724 5312 5776 5364
rect 6184 5312 6236 5364
rect 1952 5244 2004 5296
rect 4068 5176 4120 5228
rect 5632 5244 5684 5296
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 3332 5108 3384 5160
rect 5264 5176 5316 5228
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 7656 5312 7708 5364
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 8668 5355 8720 5364
rect 8668 5321 8677 5355
rect 8677 5321 8711 5355
rect 8711 5321 8720 5355
rect 8668 5312 8720 5321
rect 6552 5244 6604 5296
rect 7288 5244 7340 5296
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 6092 5108 6144 5160
rect 6460 5108 6512 5160
rect 7196 5176 7248 5228
rect 7472 5176 7524 5228
rect 5816 5040 5868 5092
rect 6644 5040 6696 5092
rect 4896 4972 4948 5024
rect 9220 5312 9272 5364
rect 10784 5312 10836 5364
rect 11704 5312 11756 5364
rect 9680 5287 9732 5296
rect 9680 5253 9689 5287
rect 9689 5253 9723 5287
rect 9723 5253 9732 5287
rect 10968 5287 11020 5296
rect 9680 5244 9732 5253
rect 7656 5108 7708 5160
rect 8116 5151 8168 5160
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 9496 5176 9548 5228
rect 10140 5219 10192 5262
rect 10140 5210 10148 5219
rect 10148 5210 10182 5219
rect 10182 5210 10192 5219
rect 10968 5253 10977 5287
rect 10977 5253 11011 5287
rect 11011 5253 11020 5287
rect 10968 5244 11020 5253
rect 11060 5244 11112 5296
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 10784 5176 10836 5228
rect 11152 5176 11204 5228
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 12716 5176 12768 5228
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 13452 5176 13504 5185
rect 8852 5040 8904 5092
rect 8944 5040 8996 5092
rect 9588 5108 9640 5160
rect 9680 5108 9732 5160
rect 10600 5108 10652 5160
rect 10140 5040 10192 5092
rect 10416 5040 10468 5092
rect 7932 4972 7984 5024
rect 9588 4972 9640 5024
rect 9772 4972 9824 5024
rect 10232 4972 10284 5024
rect 11152 5040 11204 5092
rect 13084 5040 13136 5092
rect 10968 4972 11020 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 1952 4768 2004 4820
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 4068 4768 4120 4820
rect 5080 4768 5132 4820
rect 7012 4768 7064 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 8944 4768 8996 4820
rect 9220 4811 9272 4820
rect 9220 4777 9229 4811
rect 9229 4777 9263 4811
rect 9263 4777 9272 4811
rect 9220 4768 9272 4777
rect 10600 4768 10652 4820
rect 10968 4768 11020 4820
rect 4344 4700 4396 4752
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 3056 4675 3108 4684
rect 3056 4641 3065 4675
rect 3065 4641 3099 4675
rect 3099 4641 3108 4675
rect 3056 4632 3108 4641
rect 2872 4564 2924 4616
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 4068 4632 4120 4684
rect 4528 4675 4580 4684
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 5908 4700 5960 4752
rect 7104 4700 7156 4752
rect 7656 4700 7708 4752
rect 3792 4539 3844 4548
rect 3792 4505 3801 4539
rect 3801 4505 3835 4539
rect 3835 4505 3844 4539
rect 3792 4496 3844 4505
rect 3976 4539 4028 4548
rect 3976 4505 3985 4539
rect 3985 4505 4019 4539
rect 4019 4505 4028 4539
rect 3976 4496 4028 4505
rect 5172 4632 5224 4684
rect 6644 4675 6696 4684
rect 5264 4564 5316 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 7012 4632 7064 4684
rect 8300 4700 8352 4752
rect 9404 4700 9456 4752
rect 10416 4743 10468 4752
rect 10416 4709 10425 4743
rect 10425 4709 10459 4743
rect 10459 4709 10468 4743
rect 10416 4700 10468 4709
rect 11520 4700 11572 4752
rect 13084 4743 13136 4752
rect 13084 4709 13093 4743
rect 13093 4709 13127 4743
rect 13127 4709 13136 4743
rect 13084 4700 13136 4709
rect 6184 4564 6236 4616
rect 6460 4564 6512 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 7748 4607 7800 4616
rect 6000 4496 6052 4548
rect 6644 4496 6696 4548
rect 1768 4471 1820 4480
rect 1768 4437 1777 4471
rect 1777 4437 1811 4471
rect 1811 4437 1820 4471
rect 1768 4428 1820 4437
rect 2964 4428 3016 4480
rect 3240 4428 3292 4480
rect 4252 4428 4304 4480
rect 5816 4428 5868 4480
rect 6092 4428 6144 4480
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 8668 4632 8720 4684
rect 8300 4564 8352 4616
rect 8760 4564 8812 4616
rect 9036 4564 9088 4616
rect 7012 4496 7064 4548
rect 7564 4539 7616 4548
rect 7564 4505 7573 4539
rect 7573 4505 7607 4539
rect 7607 4505 7616 4539
rect 7564 4496 7616 4505
rect 9772 4564 9824 4616
rect 9956 4564 10008 4616
rect 10600 4632 10652 4684
rect 10416 4564 10468 4616
rect 9496 4428 9548 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 10232 4428 10284 4480
rect 10784 4564 10836 4616
rect 12716 4632 12768 4684
rect 13176 4675 13228 4684
rect 13176 4641 13185 4675
rect 13185 4641 13219 4675
rect 13219 4641 13228 4675
rect 13176 4632 13228 4641
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 10692 4428 10744 4480
rect 10968 4428 11020 4480
rect 12992 4496 13044 4548
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 2688 4224 2740 4276
rect 3240 4224 3292 4276
rect 3976 4224 4028 4276
rect 4252 4224 4304 4276
rect 4528 4224 4580 4276
rect 4988 4224 5040 4276
rect 5448 4224 5500 4276
rect 5724 4224 5776 4276
rect 6736 4224 6788 4276
rect 7656 4224 7708 4276
rect 8668 4224 8720 4276
rect 9220 4224 9272 4276
rect 1768 4088 1820 4140
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 2964 4063 3016 4072
rect 2964 4029 2987 4063
rect 2987 4029 3016 4063
rect 5080 4156 5132 4208
rect 4344 4088 4396 4140
rect 4528 4088 4580 4140
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4804 4131 4856 4140
rect 4620 4088 4672 4097
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 7012 4156 7064 4208
rect 7564 4156 7616 4208
rect 4896 4088 4948 4097
rect 6000 4131 6052 4140
rect 2964 4020 3016 4029
rect 3424 4063 3476 4072
rect 3424 4029 3433 4063
rect 3433 4029 3467 4063
rect 3467 4029 3476 4063
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 3424 4020 3476 4029
rect 5632 4020 5684 4072
rect 6460 4088 6512 4140
rect 7196 4088 7248 4140
rect 7748 4088 7800 4140
rect 3148 3952 3200 4004
rect 4436 3952 4488 4004
rect 4620 3995 4672 4004
rect 4620 3961 4629 3995
rect 4629 3961 4663 3995
rect 4663 3961 4672 3995
rect 4620 3952 4672 3961
rect 6184 3952 6236 4004
rect 6828 4020 6880 4072
rect 7104 4020 7156 4072
rect 2412 3927 2464 3936
rect 2412 3893 2421 3927
rect 2421 3893 2455 3927
rect 2455 3893 2464 3927
rect 2412 3884 2464 3893
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 4712 3884 4764 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 7748 3884 7800 3936
rect 8116 4088 8168 4140
rect 9036 4088 9088 4140
rect 9496 4131 9548 4140
rect 9496 4097 9505 4131
rect 9505 4097 9539 4131
rect 9539 4097 9548 4131
rect 9496 4088 9548 4097
rect 10140 4156 10192 4208
rect 9956 4088 10008 4140
rect 10232 4088 10284 4140
rect 10416 4156 10468 4208
rect 13084 4156 13136 4208
rect 10692 4088 10744 4140
rect 11060 4088 11112 4140
rect 12808 4131 12860 4140
rect 8576 4020 8628 4072
rect 9680 4020 9732 4072
rect 10416 4020 10468 4072
rect 11980 4020 12032 4072
rect 10600 3952 10652 4004
rect 11428 3952 11480 4004
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 9864 3884 9916 3893
rect 11060 3884 11112 3936
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 13268 3952 13320 4004
rect 13176 3927 13228 3936
rect 13176 3893 13185 3927
rect 13185 3893 13219 3927
rect 13219 3893 13228 3927
rect 13176 3884 13228 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 3424 3680 3476 3732
rect 2780 3544 2832 3596
rect 3976 3544 4028 3596
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 4804 3680 4856 3732
rect 6552 3680 6604 3732
rect 4896 3612 4948 3664
rect 8760 3612 8812 3664
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 11152 3680 11204 3732
rect 2412 3408 2464 3460
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 5724 3544 5776 3596
rect 7012 3544 7064 3596
rect 9036 3587 9088 3596
rect 6092 3476 6144 3528
rect 7656 3476 7708 3528
rect 8300 3476 8352 3528
rect 5724 3408 5776 3460
rect 6184 3408 6236 3460
rect 8116 3408 8168 3460
rect 9036 3553 9045 3587
rect 9045 3553 9079 3587
rect 9079 3553 9088 3587
rect 9036 3544 9088 3553
rect 10140 3655 10192 3664
rect 10140 3621 10153 3655
rect 10153 3621 10187 3655
rect 10187 3621 10192 3655
rect 10140 3612 10192 3621
rect 10416 3612 10468 3664
rect 13268 3655 13320 3664
rect 13268 3621 13277 3655
rect 13277 3621 13311 3655
rect 13311 3621 13320 3655
rect 13268 3612 13320 3621
rect 9496 3544 9548 3596
rect 8668 3476 8720 3528
rect 9956 3476 10008 3528
rect 7472 3340 7524 3392
rect 10140 3408 10192 3460
rect 11152 3476 11204 3528
rect 11888 3544 11940 3596
rect 12808 3544 12860 3596
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 10600 3408 10652 3460
rect 9128 3340 9180 3392
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9680 3340 9732 3392
rect 10324 3340 10376 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 1584 3179 1636 3188
rect 1584 3145 1593 3179
rect 1593 3145 1627 3179
rect 1627 3145 1636 3179
rect 1584 3136 1636 3145
rect 3332 3136 3384 3188
rect 1492 3000 1544 3052
rect 3056 3068 3108 3120
rect 4068 3136 4120 3188
rect 4620 3136 4672 3188
rect 4988 3136 5040 3188
rect 4896 3068 4948 3120
rect 8116 3136 8168 3188
rect 9128 3136 9180 3188
rect 9312 3179 9364 3188
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 9588 3136 9640 3188
rect 3884 3000 3936 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 6828 3000 6880 3052
rect 3792 2932 3844 2984
rect 5724 2907 5776 2916
rect 940 2796 992 2848
rect 5724 2873 5733 2907
rect 5733 2873 5767 2907
rect 5767 2873 5776 2907
rect 5724 2864 5776 2873
rect 7196 2864 7248 2916
rect 8024 3000 8076 3052
rect 9864 3068 9916 3120
rect 10324 3136 10376 3188
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 11980 3136 12032 3188
rect 10140 3111 10192 3120
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 10140 3068 10192 3077
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9404 3000 9456 3052
rect 8392 2932 8444 2984
rect 9588 2975 9640 2984
rect 9588 2941 9601 2975
rect 9601 2941 9635 2975
rect 9635 2941 9640 2975
rect 9588 2932 9640 2941
rect 10416 3000 10468 3052
rect 10692 3068 10744 3120
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 12072 3111 12124 3120
rect 12072 3077 12081 3111
rect 12081 3077 12115 3111
rect 12115 3077 12124 3111
rect 12072 3068 12124 3077
rect 11888 3000 11940 3052
rect 9496 2864 9548 2916
rect 7288 2796 7340 2848
rect 7564 2796 7616 2848
rect 10416 2864 10468 2916
rect 11428 2932 11480 2984
rect 12072 2864 12124 2916
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 11060 2796 11112 2848
rect 11704 2796 11756 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 3976 2592 4028 2644
rect 4896 2635 4948 2644
rect 4896 2601 4905 2635
rect 4905 2601 4939 2635
rect 4939 2601 4948 2635
rect 4896 2592 4948 2601
rect 4620 2456 4672 2508
rect 3148 2388 3200 2440
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 7748 2592 7800 2644
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 10784 2592 10836 2644
rect 7196 2567 7248 2576
rect 7196 2533 7205 2567
rect 7205 2533 7239 2567
rect 7239 2533 7248 2567
rect 7196 2524 7248 2533
rect 6368 2388 6420 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 10324 2524 10376 2576
rect 10692 2456 10744 2508
rect 12716 2524 12768 2576
rect 12072 2499 12124 2508
rect 12072 2465 12081 2499
rect 12081 2465 12115 2499
rect 12115 2465 12124 2499
rect 12072 2456 12124 2465
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 8116 2388 8168 2440
rect 9680 2388 9732 2440
rect 9864 2388 9916 2440
rect 10600 2388 10652 2440
rect 10968 2388 11020 2440
rect 11704 2388 11756 2440
rect 7748 2320 7800 2372
rect 10232 2363 10284 2372
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 6460 2252 6512 2304
rect 10232 2329 10241 2363
rect 10241 2329 10275 2363
rect 10275 2329 10284 2363
rect 10232 2320 10284 2329
rect 10324 2363 10376 2372
rect 10324 2329 10333 2363
rect 10333 2329 10367 2363
rect 10367 2329 10376 2363
rect 10324 2320 10376 2329
rect 13268 2388 13320 2440
rect 13084 2363 13136 2372
rect 13084 2329 13093 2363
rect 13093 2329 13127 2363
rect 13127 2329 13136 2363
rect 13084 2320 13136 2329
rect 13176 2363 13228 2372
rect 13176 2329 13185 2363
rect 13185 2329 13219 2363
rect 13219 2329 13228 2363
rect 13176 2320 13228 2329
rect 8944 2295 8996 2304
rect 8944 2261 8953 2295
rect 8953 2261 8987 2295
rect 8987 2261 8996 2295
rect 8944 2252 8996 2261
rect 10876 2295 10928 2304
rect 10876 2261 10885 2295
rect 10885 2261 10919 2295
rect 10919 2261 10928 2295
rect 10876 2252 10928 2261
rect 12624 2252 12676 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 2228 1980 2280 2032
rect 4436 2048 4488 2100
rect 5356 2048 5408 2100
rect 10600 2048 10652 2100
rect 13176 2091 13228 2100
rect 6828 1980 6880 2032
rect 7196 1980 7248 2032
rect 7748 2023 7800 2032
rect 7748 1989 7757 2023
rect 7757 1989 7791 2023
rect 7791 1989 7800 2023
rect 7748 1980 7800 1989
rect 1400 1955 1452 1964
rect 1400 1921 1409 1955
rect 1409 1921 1443 1955
rect 1443 1921 1452 1955
rect 1400 1912 1452 1921
rect 4712 1912 4764 1964
rect 5816 1912 5868 1964
rect 6460 1955 6512 1964
rect 3240 1844 3292 1896
rect 3700 1844 3752 1896
rect 6460 1921 6469 1955
rect 6469 1921 6503 1955
rect 6503 1921 6512 1955
rect 6460 1912 6512 1921
rect 7932 1955 7984 1964
rect 7932 1921 7941 1955
rect 7941 1921 7975 1955
rect 7975 1921 7984 1955
rect 7932 1912 7984 1921
rect 10876 1980 10928 2032
rect 9864 1912 9916 1964
rect 10232 1955 10284 1964
rect 10232 1921 10241 1955
rect 10241 1921 10275 1955
rect 10275 1921 10284 1955
rect 10232 1912 10284 1921
rect 13176 2057 13185 2091
rect 13185 2057 13219 2091
rect 13219 2057 13228 2091
rect 13176 2048 13228 2057
rect 12716 1980 12768 2032
rect 11520 1955 11572 1964
rect 11520 1921 11529 1955
rect 11529 1921 11563 1955
rect 11563 1921 11572 1955
rect 11520 1912 11572 1921
rect 13360 1955 13412 1964
rect 13360 1921 13369 1955
rect 13369 1921 13403 1955
rect 13403 1921 13412 1955
rect 13360 1912 13412 1921
rect 10692 1887 10744 1896
rect 10692 1853 10701 1887
rect 10701 1853 10735 1887
rect 10735 1853 10744 1887
rect 10692 1844 10744 1853
rect 9404 1776 9456 1828
rect 10968 1776 11020 1828
rect 5632 1708 5684 1760
rect 6092 1708 6144 1760
rect 10876 1708 10928 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 2228 1547 2280 1556
rect 2228 1513 2237 1547
rect 2237 1513 2271 1547
rect 2271 1513 2280 1547
rect 2228 1504 2280 1513
rect 3148 1547 3200 1556
rect 3148 1513 3157 1547
rect 3157 1513 3191 1547
rect 3191 1513 3200 1547
rect 3148 1504 3200 1513
rect 7932 1504 7984 1556
rect 9864 1547 9916 1556
rect 9864 1513 9873 1547
rect 9873 1513 9907 1547
rect 9907 1513 9916 1547
rect 9864 1504 9916 1513
rect 10324 1504 10376 1556
rect 6828 1479 6880 1488
rect 6828 1445 6837 1479
rect 6837 1445 6871 1479
rect 6871 1445 6880 1479
rect 6828 1436 6880 1445
rect 9404 1479 9456 1488
rect 9404 1445 9413 1479
rect 9413 1445 9447 1479
rect 9447 1445 9456 1479
rect 9404 1436 9456 1445
rect 2780 1232 2832 1284
rect 3240 1300 3292 1352
rect 4712 1368 4764 1420
rect 5356 1411 5408 1420
rect 5356 1377 5365 1411
rect 5365 1377 5399 1411
rect 5399 1377 5408 1411
rect 5356 1368 5408 1377
rect 5632 1411 5684 1420
rect 5632 1377 5641 1411
rect 5641 1377 5675 1411
rect 5675 1377 5684 1411
rect 5632 1368 5684 1377
rect 5816 1300 5868 1352
rect 7564 1368 7616 1420
rect 8116 1368 8168 1420
rect 8944 1411 8996 1420
rect 8944 1377 8953 1411
rect 8953 1377 8987 1411
rect 8987 1377 8996 1411
rect 8944 1368 8996 1377
rect 10692 1368 10744 1420
rect 11520 1411 11572 1420
rect 11520 1377 11529 1411
rect 11529 1377 11563 1411
rect 11563 1377 11572 1411
rect 11520 1368 11572 1377
rect 7196 1343 7248 1352
rect 7196 1309 7205 1343
rect 7205 1309 7239 1343
rect 7239 1309 7248 1343
rect 7196 1300 7248 1309
rect 7288 1343 7340 1352
rect 7288 1309 7297 1343
rect 7297 1309 7331 1343
rect 7331 1309 7340 1343
rect 7288 1300 7340 1309
rect 3976 1232 4028 1284
rect 4620 1164 4672 1216
rect 7656 1343 7708 1352
rect 7656 1309 7665 1343
rect 7665 1309 7699 1343
rect 7699 1309 7708 1343
rect 7656 1300 7708 1309
rect 7564 1232 7616 1284
rect 10232 1300 10284 1352
rect 10876 1343 10928 1352
rect 10876 1309 10885 1343
rect 10885 1309 10919 1343
rect 10919 1309 10928 1343
rect 10876 1300 10928 1309
rect 12624 1300 12676 1352
rect 13084 1343 13136 1352
rect 13084 1309 13093 1343
rect 13093 1309 13127 1343
rect 13127 1309 13136 1343
rect 13084 1300 13136 1309
rect 13360 1343 13412 1352
rect 13360 1309 13369 1343
rect 13369 1309 13403 1343
rect 13403 1309 13412 1343
rect 13360 1300 13412 1309
rect 9680 1164 9732 1216
rect 10048 1164 10100 1216
rect 14004 1164 14056 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 9680 960 9732 1012
rect 10784 960 10836 1012
rect 13912 484 13964 536
<< metal2 >>
rect 754 14200 810 15000
rect 2226 14200 2282 15000
rect 3698 14200 3754 15000
rect 5170 14200 5226 15000
rect 6734 14200 6790 15000
rect 8206 14200 8262 15000
rect 9678 14200 9734 15000
rect 10874 14512 10930 14521
rect 10874 14447 10930 14456
rect 768 10577 796 14200
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 10674 1440 12038
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 11257 1532 11630
rect 1490 11248 1546 11257
rect 1490 11183 1546 11192
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 754 10568 810 10577
rect 754 10503 810 10512
rect 1412 9518 1440 10610
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 10266 1716 10542
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 2240 9994 2268 14200
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2516 12102 2544 12922
rect 3344 12918 3372 13126
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2516 11694 2544 12038
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2608 11286 2636 12718
rect 3436 12238 3464 13262
rect 3712 12434 3740 14200
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 5184 13410 5212 14200
rect 6748 13546 6776 14200
rect 5540 13524 5592 13530
rect 6748 13518 6868 13546
rect 8220 13530 8248 14200
rect 9692 13546 9720 14200
rect 5540 13466 5592 13472
rect 5184 13382 5488 13410
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4632 12442 4660 12718
rect 4620 12436 4672 12442
rect 3712 12406 4108 12434
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 2964 12232 3016 12238
rect 2884 12180 2964 12186
rect 2884 12174 3016 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2884 12158 3004 12174
rect 2700 11898 2728 12106
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2884 11762 2912 12158
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2884 11558 2912 11698
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2320 10736 2372 10742
rect 2320 10678 2372 10684
rect 2332 10266 2360 10678
rect 2884 10266 2912 11494
rect 3160 11014 3188 12038
rect 3528 11354 3556 12310
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11830 3924 12038
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3528 11150 3556 11290
rect 3804 11286 3832 11630
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3516 11144 3568 11150
rect 3608 11144 3660 11150
rect 3516 11086 3568 11092
rect 3606 11112 3608 11121
rect 3660 11112 3662 11121
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2884 10062 2912 10202
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 7954 1440 9454
rect 2240 9178 2268 9590
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 8498 1900 8910
rect 2792 8650 2820 9318
rect 2884 9110 2912 9998
rect 3160 9994 3188 10950
rect 3252 10062 3280 11086
rect 3896 11082 3924 11222
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3606 11047 3662 11056
rect 3884 11076 3936 11082
rect 3620 10742 3648 11047
rect 3884 11018 3936 11024
rect 3988 11014 4016 11086
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10130 3464 10406
rect 3804 10248 3832 10542
rect 3712 10220 3832 10248
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3712 10062 3740 10220
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 2976 9722 3004 9930
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2792 8622 3004 8650
rect 2792 8498 2820 8622
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7342 1440 7890
rect 1964 7818 1992 8298
rect 2424 8090 2452 8434
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 6254 1440 7278
rect 2240 7002 2268 7414
rect 2424 7342 2452 8026
rect 2700 7818 2728 8230
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2884 7562 2912 8502
rect 2976 8378 3004 8622
rect 3068 8566 3096 9862
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 8974 3372 9454
rect 3620 9450 3648 9522
rect 3712 9500 3740 9998
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 3804 9654 3832 9930
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3896 9518 3924 10542
rect 3792 9512 3844 9518
rect 3712 9472 3792 9500
rect 3792 9454 3844 9460
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8634 3372 8774
rect 3436 8634 3464 9046
rect 3804 8838 3832 9454
rect 4080 8922 4108 12406
rect 4620 12378 4672 12384
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4632 11354 4660 12174
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4632 11234 4660 11290
rect 4264 11206 4660 11234
rect 4264 11150 4292 11206
rect 4724 11150 4752 12922
rect 5184 12238 5212 13194
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12306 5396 13126
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5092 11898 5120 12106
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5092 11558 5120 11834
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4252 11144 4304 11150
rect 4160 11122 4212 11128
rect 4158 11112 4160 11121
rect 4212 11112 4214 11121
rect 4252 11086 4304 11092
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4158 11047 4214 11056
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4172 10674 4200 10950
rect 4816 10742 4844 11154
rect 4894 11112 4950 11121
rect 5092 11082 5120 11494
rect 4894 11047 4896 11056
rect 4948 11047 4950 11056
rect 5080 11076 5132 11082
rect 4896 11018 4948 11024
rect 5080 11018 5132 11024
rect 4908 10810 4936 11018
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4632 10266 4660 10542
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4356 9518 4384 10134
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4632 9178 4660 10066
rect 4724 10062 4752 10406
rect 4802 10160 4858 10169
rect 4802 10095 4858 10104
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4816 9908 4844 10095
rect 4724 9880 4844 9908
rect 4724 9586 4752 9880
rect 4908 9674 4936 10746
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 10044 5120 10406
rect 5184 10169 5212 12174
rect 5368 11558 5396 12242
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5276 10674 5304 11494
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5276 10538 5304 10610
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10266 5396 10406
rect 5460 10266 5488 13382
rect 5552 12918 5580 13466
rect 6840 13394 6868 13518
rect 8208 13524 8260 13530
rect 9692 13518 9904 13546
rect 8208 13466 8260 13472
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5920 12442 5948 13330
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6012 12986 6040 13262
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11762 5580 12174
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5920 11150 5948 12378
rect 6012 12102 6040 12922
rect 6564 12918 6592 13194
rect 6840 12986 6868 13194
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6932 12918 6960 13398
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11762 6040 12038
rect 6564 11762 6592 12854
rect 7024 12238 7052 13126
rect 7576 12306 7604 13126
rect 7944 12986 7972 13262
rect 8220 13240 8248 13466
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 8128 13212 8248 13240
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8128 12850 8156 13212
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 8214 13084 8522 13104
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13008 8522 13028
rect 8588 12850 8616 13126
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6748 11898 6776 12106
rect 6736 11892 6788 11898
rect 6656 11852 6736 11880
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6274 11112 6330 11121
rect 5736 11014 5764 11086
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5552 10674 5580 10950
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5170 10160 5226 10169
rect 5170 10095 5226 10104
rect 5264 10056 5316 10062
rect 5092 10024 5264 10044
rect 5448 10056 5500 10062
rect 5316 10024 5318 10033
rect 5092 10016 5262 10024
rect 5448 9998 5500 10004
rect 5262 9959 5318 9968
rect 4816 9646 4936 9674
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4080 8894 4200 8922
rect 4172 8838 4200 8894
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2976 8350 3096 8378
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7954 3004 8230
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2884 7546 3004 7562
rect 2884 7540 3016 7546
rect 2884 7534 2964 7540
rect 2964 7482 3016 7488
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2332 6934 2360 7278
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2792 6662 2820 7142
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 1400 6248 1452 6254
rect 1452 6208 1532 6236
rect 1400 6190 1452 6196
rect 1504 3534 1532 6208
rect 2332 5914 2360 6326
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2792 5846 2820 6598
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2884 5710 2912 6938
rect 2976 6798 3004 7482
rect 3068 7410 3096 8350
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3344 6934 3372 8570
rect 3436 7886 3464 8570
rect 3896 8566 3924 8774
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4724 8498 4752 9522
rect 4816 9518 4844 9646
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4908 8634 4936 9522
rect 5000 9178 5028 9522
rect 5460 9450 5488 9998
rect 5552 9654 5580 10610
rect 5644 10130 5672 10678
rect 5736 10470 5764 10950
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5814 10160 5870 10169
rect 5632 10124 5684 10130
rect 5814 10095 5870 10104
rect 5920 10112 5948 11086
rect 6104 10742 6132 11086
rect 6274 11047 6330 11056
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 6000 10124 6052 10130
rect 5632 10066 5684 10072
rect 5828 10062 5856 10095
rect 5920 10084 6000 10112
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9674 5672 9930
rect 5540 9648 5592 9654
rect 5644 9646 5764 9674
rect 5540 9590 5592 9596
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5184 9042 5212 9318
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5448 8900 5500 8906
rect 5552 8888 5580 9454
rect 5500 8860 5580 8888
rect 5448 8842 5500 8848
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 7206 3464 7822
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3896 7478 3924 7686
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3608 6928 3660 6934
rect 3712 6916 3740 7346
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3804 6934 3832 7278
rect 3660 6888 3740 6916
rect 3608 6870 3660 6876
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 6118 3188 6734
rect 3712 6662 3740 6888
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3896 6798 3924 7414
rect 3988 7274 4016 7686
rect 4632 7426 4660 7890
rect 5460 7818 5488 8842
rect 5736 7886 5764 9646
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5828 9382 5856 9590
rect 5920 9586 5948 10084
rect 6000 10066 6052 10072
rect 6288 9926 6316 11047
rect 6472 11014 6500 11290
rect 6656 11218 6684 11852
rect 6736 11834 6788 11840
rect 7208 11762 7236 12174
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10724 6500 10950
rect 6552 10736 6604 10742
rect 6472 10696 6552 10724
rect 6552 10678 6604 10684
rect 6656 10674 6684 11154
rect 6748 11150 6776 11630
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11150 6868 11494
rect 7208 11354 7236 11698
rect 8036 11694 8064 12242
rect 8404 12238 8432 12650
rect 9140 12434 9168 12786
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 8864 12406 9168 12434
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8214 11996 8522 12016
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11920 8522 11940
rect 8588 11898 8616 12174
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8680 11694 8708 12106
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 11762 8800 12038
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6840 10606 6868 11086
rect 6828 10600 6880 10606
rect 6642 10568 6698 10577
rect 6828 10542 6880 10548
rect 6642 10503 6698 10512
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6380 9654 6408 10134
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 8566 5856 9318
rect 5920 8634 5948 9522
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6196 8634 6224 8842
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 4632 7410 4844 7426
rect 4620 7404 4844 7410
rect 4672 7398 4844 7404
rect 4620 7346 4672 7352
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4632 7002 4660 7210
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3804 6390 3832 6734
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5710 3188 6054
rect 3620 5914 3648 6258
rect 3896 6236 3924 6598
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3804 6208 3924 6236
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3804 5658 3832 6208
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5778 3924 6054
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 1780 5574 1808 5646
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1780 4486 1808 5510
rect 2884 5370 2912 5646
rect 3804 5630 3924 5658
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 1952 5296 2004 5302
rect 1952 5238 2004 5244
rect 1964 4826 1992 5238
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 4146 1808 4422
rect 2700 4282 2728 4626
rect 2884 4622 2912 5306
rect 3344 5166 3372 5510
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 2976 4826 3004 5102
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 2976 4078 3004 4422
rect 3068 4146 3096 4626
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4282 3280 4422
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 1582 3768 1638 3777
rect 1582 3703 1638 3712
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1504 3058 1532 3470
rect 1596 3194 1624 3703
rect 2424 3466 2452 3878
rect 2792 3602 2820 3878
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 952 800 980 2790
rect 1400 1964 1452 1970
rect 1504 1952 1532 2994
rect 3068 2650 3096 3062
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3160 2446 3188 3946
rect 3344 3194 3372 5102
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3436 4185 3464 4558
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 3738 3464 4014
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3804 2990 3832 4490
rect 3896 3482 3924 5630
rect 3988 4554 4016 6394
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4080 5846 4108 6258
rect 4448 6186 4476 6802
rect 4724 6730 4752 7278
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4632 5642 4660 6122
rect 4724 5914 4752 6258
rect 4816 6254 4844 7398
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4724 5370 4752 5850
rect 4908 5846 4936 6598
rect 5000 5914 5028 6870
rect 5092 6798 5120 7142
rect 5184 6866 5212 7346
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4908 5250 4936 5782
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4632 5222 4936 5250
rect 4080 4826 4108 5170
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3988 4282 4016 4490
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3988 3602 4016 4218
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3896 3454 4016 3482
rect 3882 3088 3938 3097
rect 3882 3023 3884 3032
rect 3936 3023 3938 3032
rect 3884 2994 3936 3000
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 1452 1924 1532 1952
rect 1400 1906 1452 1912
rect 2240 1562 2268 1974
rect 3160 1562 3188 2382
rect 3240 1896 3292 1902
rect 3240 1838 3292 1844
rect 3700 1896 3752 1902
rect 3896 1884 3924 2994
rect 3988 2650 4016 3454
rect 4080 3194 4108 4626
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 4282 4292 4422
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4356 4146 4384 4694
rect 4528 4684 4580 4690
rect 4448 4644 4528 4672
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4448 4010 4476 4644
rect 4528 4626 4580 4632
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4540 4146 4568 4218
rect 4632 4146 4660 5222
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4146 4936 4966
rect 5092 4826 5120 5102
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3194 4660 3946
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4724 3534 4752 3878
rect 4816 3738 4844 4082
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4908 3670 4936 4082
rect 5000 4026 5028 4218
rect 5092 4214 5120 4762
rect 5184 4690 5212 6802
rect 5460 6798 5488 7754
rect 5736 7478 5764 7822
rect 5828 7478 5856 8502
rect 6564 8090 6592 9658
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5276 5574 5304 6734
rect 5644 6458 5672 7278
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 7002 5856 7142
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5184 4026 5212 4626
rect 5276 4622 5304 5170
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5368 4185 5396 6054
rect 5644 5914 5672 6394
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5644 5302 5672 5850
rect 5736 5778 5764 6666
rect 5920 6458 5948 7346
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5828 5846 5856 6258
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5736 5370 5764 5714
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4282 5488 4558
rect 5736 4282 5764 5306
rect 5828 5098 5856 5578
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5828 4486 5856 5034
rect 5920 4758 5948 6258
rect 6012 6186 6040 6394
rect 6104 6390 6132 7142
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6092 6112 6144 6118
rect 6012 6060 6092 6066
rect 6012 6054 6144 6060
rect 6012 6038 6132 6054
rect 6012 5778 6040 6038
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6196 5710 6224 7890
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6730 6500 7142
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6656 6322 6684 10503
rect 6932 10266 6960 11222
rect 7392 11150 7420 11630
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11218 8708 11494
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 7196 11144 7248 11150
rect 7380 11144 7432 11150
rect 7196 11086 7248 11092
rect 7378 11112 7380 11121
rect 7432 11112 7434 11121
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10606 7144 11018
rect 7208 10742 7236 11086
rect 7378 11047 7434 11056
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 8128 10674 8156 10950
rect 8214 10908 8522 10928
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10832 8522 10852
rect 8864 10690 8892 12406
rect 9232 12238 9260 12650
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9324 11830 9352 12310
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8956 10826 8984 11086
rect 8956 10798 9076 10826
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8772 10662 8892 10690
rect 8944 10668 8996 10674
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7116 10266 7144 10542
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9382 6868 9862
rect 6932 9722 6960 9998
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 7208 9178 7236 10066
rect 7300 10062 7328 10610
rect 8128 10266 8156 10610
rect 8588 10266 8616 10610
rect 8680 10470 8708 10610
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8128 10062 8156 10202
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 7288 10056 7340 10062
rect 8116 10056 8168 10062
rect 7288 9998 7340 10004
rect 8022 10024 8078 10033
rect 8116 9998 8168 10004
rect 8022 9959 8078 9968
rect 8036 9674 8064 9959
rect 8588 9926 8616 10066
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8214 9820 8522 9840
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9744 8522 9764
rect 8036 9646 8156 9674
rect 8128 9602 8156 9646
rect 8128 9586 8340 9602
rect 8588 9586 8616 9862
rect 8128 9580 8352 9586
rect 8128 9574 8300 9580
rect 8300 9522 8352 9528
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7024 8498 7052 8910
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7944 8634 7972 8842
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7024 8090 7052 8434
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7760 7954 7788 8230
rect 8036 8022 8064 8842
rect 8214 8732 8522 8752
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8656 8522 8676
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7024 7478 7052 7686
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 6662 7420 7278
rect 7484 6798 7512 7346
rect 7852 6934 7880 7414
rect 7944 7342 7972 7686
rect 8036 7478 8064 7822
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8036 7274 8064 7414
rect 8128 7410 8156 8434
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8214 7644 8522 7664
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7568 8522 7588
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7010 6488 7066 6497
rect 7010 6423 7066 6432
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6274 6216 6330 6225
rect 6274 6151 6330 6160
rect 6460 6180 6512 6186
rect 6288 5710 6316 6151
rect 6460 6122 6512 6128
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6196 5370 6224 5646
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5354 4176 5410 4185
rect 5354 4111 5410 4120
rect 5630 4176 5686 4185
rect 5630 4111 5686 4120
rect 5644 4078 5672 4111
rect 5000 3998 5212 4026
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 5736 3602 5764 4218
rect 5920 4049 5948 4694
rect 6012 4672 6040 5170
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6104 5001 6132 5102
rect 6090 4992 6146 5001
rect 6090 4927 6146 4936
rect 6012 4644 6132 4672
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6012 4146 6040 4490
rect 6104 4486 6132 4644
rect 6196 4622 6224 5306
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5906 4040 5962 4049
rect 6196 4010 6224 4558
rect 5906 3975 5962 3984
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6288 3641 6316 5646
rect 6274 3632 6330 3641
rect 5724 3596 5776 3602
rect 6274 3567 6330 3576
rect 5724 3538 5776 3544
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4908 2650 4936 3062
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3752 1856 3924 1884
rect 3700 1838 3752 1844
rect 2228 1556 2280 1562
rect 2228 1498 2280 1504
rect 3148 1556 3200 1562
rect 3148 1498 3200 1504
rect 3252 1358 3280 1838
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 3988 1290 4016 2246
rect 4448 2106 4476 2382
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 4214 1660 4522 1680
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1584 4522 1604
rect 2780 1284 2832 1290
rect 2780 1226 2832 1232
rect 3976 1284 4028 1290
rect 3976 1226 4028 1232
rect 2792 800 2820 1226
rect 4632 1222 4660 2450
rect 4712 1964 4764 1970
rect 4712 1906 4764 1912
rect 4724 1426 4752 1906
rect 4712 1420 4764 1426
rect 4712 1362 4764 1368
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 4632 870 4752 898
rect 4632 800 4660 870
rect 938 0 994 800
rect 2778 0 2834 800
rect 4618 0 4674 800
rect 4724 762 4752 870
rect 5000 762 5028 3130
rect 5736 2922 5764 3402
rect 6104 3097 6132 3470
rect 6184 3460 6236 3466
rect 6288 3448 6316 3567
rect 6236 3420 6316 3448
rect 6184 3402 6236 3408
rect 6090 3088 6146 3097
rect 6380 3058 6408 6054
rect 6472 5846 6500 6122
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6656 5386 6684 6258
rect 7024 6254 7052 6423
rect 7392 6322 7420 6598
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5846 6960 6054
rect 7300 5914 7328 6258
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6932 5642 6960 5782
rect 7024 5642 7052 5850
rect 7196 5704 7248 5710
rect 7194 5672 7196 5681
rect 7288 5704 7340 5710
rect 7248 5672 7250 5681
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 7012 5636 7064 5642
rect 7288 5646 7340 5652
rect 7194 5607 7250 5616
rect 7012 5578 7064 5584
rect 6564 5358 6684 5386
rect 6564 5302 6592 5358
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6472 4622 6500 5102
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6656 4690 6684 5034
rect 7024 4826 7052 5578
rect 7300 5302 7328 5646
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 6644 4684 6696 4690
rect 7012 4684 7064 4690
rect 6644 4626 6696 4632
rect 6840 4644 7012 4672
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6472 4146 6500 4558
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6656 4185 6684 4490
rect 6748 4282 6776 4558
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6642 4176 6698 4185
rect 6460 4140 6512 4146
rect 6642 4111 6698 4120
rect 6460 4082 6512 4088
rect 6840 4078 6868 4644
rect 7012 4626 7064 4632
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7024 4214 7052 4490
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 7116 4078 7144 4694
rect 7208 4146 7236 5170
rect 7392 5114 7420 6258
rect 7484 5234 7512 6734
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7852 6118 7880 6666
rect 8022 6488 8078 6497
rect 8022 6423 8024 6432
rect 8076 6423 8078 6432
rect 8024 6394 8076 6400
rect 8128 6338 8156 7346
rect 8588 7206 8616 7890
rect 8680 7546 8708 9930
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8214 6556 8522 6576
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6480 8522 6500
rect 8036 6322 8156 6338
rect 8024 6316 8156 6322
rect 8076 6310 8156 6316
rect 8024 6258 8076 6264
rect 7564 6112 7616 6118
rect 7840 6112 7892 6118
rect 7564 6054 7616 6060
rect 7654 6080 7710 6089
rect 7576 5914 7604 6054
rect 7840 6054 7892 6060
rect 7654 6015 7710 6024
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7668 5846 7696 6015
rect 7656 5840 7708 5846
rect 7656 5782 7708 5788
rect 7668 5370 7696 5782
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7656 5160 7708 5166
rect 7562 5128 7618 5137
rect 7392 5086 7512 5114
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6090 3023 6146 3032
rect 6368 3052 6420 3058
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5368 1426 5396 2042
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 5632 1760 5684 1766
rect 5632 1702 5684 1708
rect 5644 1426 5672 1702
rect 5356 1420 5408 1426
rect 5356 1362 5408 1368
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5828 1358 5856 1906
rect 6104 1766 6132 3023
rect 6368 2994 6420 3000
rect 6380 2446 6408 2994
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 1970 6500 2246
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 6092 1760 6144 1766
rect 6092 1702 6144 1708
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 6564 800 6592 3674
rect 7024 3602 7052 3878
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7484 3398 7512 5086
rect 7656 5102 7708 5108
rect 7562 5063 7618 5072
rect 7576 4554 7604 5063
rect 7668 4758 7696 5102
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7576 4214 7604 4490
rect 7668 4282 7696 4694
rect 7760 4622 7788 5714
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7852 5370 7880 5510
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4826 7972 4966
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7760 4146 7788 4558
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7668 3534 7696 3878
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6840 2038 6868 2994
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7208 2582 7236 2858
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7208 2038 7236 2382
rect 6828 2032 6880 2038
rect 6828 1974 6880 1980
rect 7196 2032 7248 2038
rect 7196 1974 7248 1980
rect 6840 1494 6868 1974
rect 6828 1488 6880 1494
rect 6828 1430 6880 1436
rect 7208 1358 7236 1974
rect 7300 1358 7328 2790
rect 7576 1426 7604 2790
rect 7760 2650 7788 3878
rect 8036 3058 8064 6258
rect 8588 6118 8616 7142
rect 8772 6934 8800 10662
rect 8944 10610 8996 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 9722 8892 10542
rect 8956 10198 8984 10610
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8944 10056 8996 10062
rect 9048 10044 9076 10798
rect 9140 10062 9168 11562
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11218 9352 11494
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9416 11150 9444 12106
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9232 10810 9260 11086
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 8996 10016 9076 10044
rect 9128 10056 9180 10062
rect 8944 9998 8996 10004
rect 9128 9998 9180 10004
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8956 9654 8984 9998
rect 9324 9674 9352 11018
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10810 9444 10950
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9416 10062 9444 10474
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9232 9646 9352 9674
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8864 9178 8892 9454
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9048 8566 9076 8978
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9048 8294 9076 8502
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8090 9076 8230
rect 9036 8084 9088 8090
rect 8956 8044 9036 8072
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 7410 8892 7822
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8864 6322 8892 7346
rect 8956 6458 8984 8044
rect 9036 8026 9088 8032
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9048 7478 9076 7822
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 9232 7342 9260 9646
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 7886 9444 8774
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6934 9076 7142
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 9048 6662 9076 6870
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6458 9076 6598
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5953 8616 6054
rect 8574 5944 8630 5953
rect 8574 5879 8630 5888
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 5166 8156 5510
rect 8214 5468 8522 5488
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5392 8522 5412
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8128 4146 8156 5102
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8312 4622 8340 4694
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8214 4380 8522 4400
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4304 8522 4324
rect 8588 4264 8616 5879
rect 8864 5710 8892 6258
rect 8956 5846 8984 6394
rect 9048 6254 9076 6394
rect 9036 6248 9088 6254
rect 9034 6216 9036 6225
rect 9088 6216 9090 6225
rect 9034 6151 9090 6160
rect 9140 6118 9168 6802
rect 9232 6118 9260 7278
rect 9324 7002 9352 7822
rect 9416 7410 9444 7822
rect 9508 7546 9536 13126
rect 9784 12850 9812 13398
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11694 9720 12106
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9784 11150 9812 11834
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9678 10976 9734 10985
rect 9600 7818 9628 10950
rect 9678 10911 9734 10920
rect 9692 10810 9720 10911
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 9178 9720 9522
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9784 7410 9812 11086
rect 9876 10810 9904 13518
rect 10506 13424 10562 13433
rect 10506 13359 10562 13368
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12782 10088 13126
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10138 12744 10194 12753
rect 10060 12646 10088 12718
rect 10138 12679 10194 12688
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11937 9996 12038
rect 9954 11928 10010 11937
rect 9954 11863 10010 11872
rect 10060 11830 10088 12582
rect 10152 12442 10180 12679
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10152 12170 10180 12378
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10048 11824 10100 11830
rect 9968 11772 10048 11778
rect 9968 11766 10100 11772
rect 9968 11750 10088 11766
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9968 10606 9996 11750
rect 10336 11694 10364 12174
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10198 9996 10542
rect 10060 10266 10088 11630
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 11150 10272 11494
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10152 10810 10180 11018
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10244 10674 10272 11086
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10428 10198 10456 10406
rect 9956 10192 10008 10198
rect 10416 10192 10468 10198
rect 9956 10134 10008 10140
rect 10414 10160 10416 10169
rect 10468 10160 10470 10169
rect 10414 10095 10470 10104
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10152 8634 10180 9522
rect 10336 9110 10364 9590
rect 10520 9518 10548 13359
rect 10888 12646 10916 14447
rect 11242 14200 11298 15000
rect 12714 14200 12770 15000
rect 14186 14200 14242 15000
rect 11256 13410 11284 14200
rect 12214 13628 12522 13648
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13552 12522 13572
rect 12728 13410 12756 14200
rect 11256 13382 11468 13410
rect 12728 13382 12848 13410
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10888 12442 10916 12582
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 11072 12238 11100 13126
rect 11348 12918 11376 13262
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11256 12238 11284 12786
rect 11348 12306 11376 12854
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11072 11762 11100 12174
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11830 11192 12038
rect 11256 11898 11284 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 10888 11558 10916 11698
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 11256 11286 11284 11698
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11256 10742 11284 11222
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10888 9450 10916 10202
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9654 11100 9930
rect 11164 9926 11192 9998
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10690 9072 10746 9081
rect 10690 9007 10746 9016
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10520 8566 10548 8774
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9968 7410 9996 7822
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9128 6112 9180 6118
rect 9126 6080 9128 6089
rect 9220 6112 9272 6118
rect 9180 6080 9182 6089
rect 9220 6054 9272 6060
rect 9126 6015 9182 6024
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 9324 5710 9352 6938
rect 9416 6322 9444 7346
rect 9784 6934 9812 7346
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5760 9444 6054
rect 9494 5944 9550 5953
rect 9494 5879 9496 5888
rect 9548 5879 9550 5888
rect 9678 5944 9734 5953
rect 9678 5879 9680 5888
rect 9496 5850 9548 5856
rect 9732 5879 9734 5888
rect 9680 5850 9732 5856
rect 9586 5808 9642 5817
rect 9416 5732 9536 5760
rect 9586 5743 9642 5752
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8852 5704 8904 5710
rect 9220 5704 9272 5710
rect 8852 5646 8904 5652
rect 9218 5672 9220 5681
rect 9312 5704 9364 5710
rect 9272 5672 9274 5681
rect 8680 5370 8708 5646
rect 9312 5646 9364 5652
rect 9402 5672 9458 5681
rect 9218 5607 9274 5616
rect 9036 5568 9088 5574
rect 8758 5536 8814 5545
rect 9036 5510 9088 5516
rect 8758 5471 8814 5480
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8680 4690 8708 5306
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4282 8708 4626
rect 8772 4622 8800 5471
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8312 4236 8616 4264
rect 8668 4276 8720 4282
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8312 4049 8340 4236
rect 8668 4218 8720 4224
rect 8576 4072 8628 4078
rect 8298 4040 8354 4049
rect 8576 4014 8628 4020
rect 8298 3975 8354 3984
rect 8312 3534 8340 3975
rect 8300 3528 8352 3534
rect 8298 3496 8300 3505
rect 8352 3496 8354 3505
rect 8116 3460 8168 3466
rect 8298 3431 8354 3440
rect 8116 3402 8168 3408
rect 8128 3194 8156 3402
rect 8214 3292 8522 3312
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3216 8522 3236
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8404 2650 8432 2926
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 7760 2514 7788 2586
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7668 1358 7696 2382
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7760 2038 7788 2314
rect 7748 2032 7800 2038
rect 7748 1974 7800 1980
rect 7932 1964 7984 1970
rect 7932 1906 7984 1912
rect 7944 1562 7972 1906
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 8128 1426 8156 2382
rect 8214 2204 8522 2224
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2128 8522 2148
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 7288 1352 7340 1358
rect 7656 1352 7708 1358
rect 7340 1300 7604 1306
rect 7288 1294 7604 1300
rect 7656 1294 7708 1300
rect 7300 1290 7604 1294
rect 7300 1284 7616 1290
rect 7300 1278 7564 1284
rect 7564 1226 7616 1232
rect 8214 1116 8522 1136
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1040 8522 1060
rect 8588 898 8616 4014
rect 8772 3670 8800 4558
rect 8864 4049 8892 5034
rect 8956 4865 8984 5034
rect 8942 4856 8998 4865
rect 8942 4791 8944 4800
rect 8996 4791 8998 4800
rect 8944 4762 8996 4768
rect 9048 4622 9076 5510
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 4826 9260 5306
rect 9324 5137 9352 5646
rect 9402 5607 9458 5616
rect 9310 5128 9366 5137
rect 9310 5063 9366 5072
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9416 4758 9444 5607
rect 9508 5545 9536 5732
rect 9600 5658 9628 5743
rect 9784 5658 9812 6870
rect 9968 6866 9996 7346
rect 10060 7002 10088 7822
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 7546 10180 7686
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10152 6882 10180 7210
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 10060 6854 10180 6882
rect 10232 6860 10284 6866
rect 10060 6730 10088 6854
rect 10232 6802 10284 6808
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10060 5846 10088 6666
rect 10244 6458 10272 6802
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10336 6322 10364 6598
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5846 10272 6054
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 9600 5630 9812 5658
rect 9956 5568 10008 5574
rect 9494 5536 9550 5545
rect 9956 5510 10008 5516
rect 9494 5471 9550 5480
rect 9508 5234 9536 5471
rect 9678 5298 9734 5307
rect 9968 5250 9996 5510
rect 9496 5228 9548 5234
rect 9678 5233 9734 5242
rect 9876 5222 9996 5250
rect 9876 5216 9904 5222
rect 9496 5170 9548 5176
rect 9784 5188 9904 5216
rect 9588 5160 9640 5166
rect 9586 5128 9588 5137
rect 9680 5160 9732 5166
rect 9640 5128 9642 5137
rect 9784 5148 9812 5188
rect 9732 5120 9812 5148
rect 9680 5102 9732 5108
rect 9586 5063 9642 5072
rect 9588 5024 9640 5030
rect 9586 4992 9588 5001
rect 9772 5024 9824 5030
rect 9640 4992 9642 5001
rect 9586 4927 9642 4936
rect 9770 4992 9772 5001
rect 10060 5001 10088 5782
rect 10244 5710 10272 5782
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5262 10192 5268
rect 10336 5234 10364 6258
rect 10428 5914 10456 8434
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6458 10640 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10140 5204 10192 5210
rect 10324 5228 10376 5234
rect 10152 5098 10180 5204
rect 10324 5170 10376 5176
rect 10428 5098 10456 5646
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10232 5024 10284 5030
rect 9824 4992 9826 5001
rect 9770 4927 9826 4936
rect 10046 4992 10102 5001
rect 10102 4950 10180 4978
rect 10232 4966 10284 4972
rect 10046 4927 10102 4936
rect 10060 4867 10088 4927
rect 9954 4856 10010 4865
rect 9954 4791 10010 4800
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9770 4720 9826 4729
rect 9770 4655 9826 4664
rect 9784 4622 9812 4655
rect 9968 4622 9996 4791
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9496 4480 9548 4486
rect 9218 4448 9274 4457
rect 10048 4480 10100 4486
rect 9496 4422 9548 4428
rect 9586 4448 9642 4457
rect 9218 4383 9274 4392
rect 9232 4282 9260 4383
rect 9402 4312 9458 4321
rect 9220 4276 9272 4282
rect 9402 4247 9458 4256
rect 9220 4218 9272 4224
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 8850 4040 8906 4049
rect 8850 3975 8906 3984
rect 8760 3664 8812 3670
rect 8666 3632 8722 3641
rect 8760 3606 8812 3612
rect 9048 3602 9076 4082
rect 8666 3567 8722 3576
rect 9036 3596 9088 3602
rect 8680 3534 8708 3567
rect 9036 3538 9088 3544
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 9048 3058 9076 3538
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9140 3194 9168 3334
rect 9324 3194 9352 3334
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9416 3058 9444 4247
rect 9508 4146 9536 4422
rect 9642 4406 9720 4434
rect 10048 4422 10100 4428
rect 9586 4383 9642 4392
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9692 4078 9720 4406
rect 9862 4176 9918 4185
rect 9862 4111 9918 4120
rect 9956 4140 10008 4146
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9876 3942 9904 4111
rect 9956 4082 10008 4088
rect 9864 3936 9916 3942
rect 9678 3904 9734 3913
rect 9864 3878 9916 3884
rect 9678 3839 9734 3848
rect 9692 3738 9720 3839
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9508 2922 9536 3538
rect 9968 3534 9996 4082
rect 9956 3528 10008 3534
rect 9586 3496 9642 3505
rect 9956 3470 10008 3476
rect 9586 3431 9642 3440
rect 9600 3194 9628 3431
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9600 2990 9628 3130
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9692 2446 9720 3334
rect 9864 3120 9916 3126
rect 9862 3088 9864 3097
rect 9916 3088 9918 3097
rect 9862 3023 9918 3032
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 1426 8984 2246
rect 9876 1970 9904 2382
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 9404 1828 9456 1834
rect 9404 1770 9456 1776
rect 9416 1494 9444 1770
rect 9876 1562 9904 1906
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 9404 1488 9456 1494
rect 9404 1430 9456 1436
rect 8944 1420 8996 1426
rect 8944 1362 8996 1368
rect 10060 1222 10088 4422
rect 10152 4214 10180 4950
rect 10244 4486 10272 4966
rect 10428 4758 10456 5034
rect 10416 4752 10468 4758
rect 10336 4712 10416 4740
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10152 3670 10180 4150
rect 10244 4146 10272 4422
rect 10336 4185 10364 4712
rect 10416 4694 10468 4700
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10428 4214 10456 4558
rect 10416 4208 10468 4214
rect 10322 4176 10378 4185
rect 10232 4140 10284 4146
rect 10416 4150 10468 4156
rect 10322 4111 10378 4120
rect 10232 4082 10284 4088
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 10152 3126 10180 3402
rect 10336 3398 10364 4111
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3670 10456 4014
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10336 3194 10364 3334
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10336 3058 10456 3074
rect 10336 3052 10468 3058
rect 10336 3046 10416 3052
rect 10336 2582 10364 3046
rect 10416 2994 10468 3000
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10244 1970 10272 2314
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 10244 1358 10272 1906
rect 10336 1562 10364 2314
rect 10324 1556 10376 1562
rect 10324 1498 10376 1504
rect 10232 1352 10284 1358
rect 10232 1294 10284 1300
rect 9680 1216 9732 1222
rect 9680 1158 9732 1164
rect 10048 1216 10100 1222
rect 10428 1170 10456 2858
rect 10520 2122 10548 6122
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10612 5166 10640 5782
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10612 4826 10640 5102
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 4010 10640 4626
rect 10704 4486 10732 9007
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7954 10824 8230
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10796 6390 10824 7890
rect 10888 7324 10916 8026
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7546 11008 7686
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10968 7336 11020 7342
rect 10888 7296 10968 7324
rect 10968 7278 11020 7284
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10888 6202 10916 6326
rect 10796 6174 10916 6202
rect 10796 5846 10824 6174
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10888 5574 10916 6054
rect 10980 5681 11008 7278
rect 11072 7002 11100 7822
rect 11164 7546 11192 9862
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11256 8974 11284 9522
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11164 6798 11192 7346
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 5704 11112 5710
rect 10966 5672 11022 5681
rect 11060 5646 11112 5652
rect 10966 5607 11022 5616
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10966 5536 11022 5545
rect 10796 5370 10824 5510
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10796 4978 10824 5170
rect 10888 5137 10916 5510
rect 10966 5471 11022 5480
rect 10980 5302 11008 5471
rect 11072 5302 11100 5646
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10874 5128 10930 5137
rect 10980 5114 11008 5238
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 10980 5086 11100 5114
rect 11164 5098 11192 5170
rect 10874 5063 10930 5072
rect 10968 5024 11020 5030
rect 10796 4972 10968 4978
rect 10796 4966 11020 4972
rect 10796 4950 11008 4966
rect 10796 4622 10824 4950
rect 11072 4865 11100 5086
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11058 4856 11114 4865
rect 10968 4820 11020 4826
rect 11058 4791 11114 4800
rect 10968 4762 11020 4768
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10980 4570 11008 4762
rect 10980 4542 11100 4570
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10612 2446 10640 3402
rect 10704 3126 10732 4082
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10796 2650 10824 2994
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10980 2530 11008 4422
rect 11072 4146 11100 4542
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 2854 11100 3878
rect 11164 3738 11192 5034
rect 11256 3913 11284 8910
rect 11348 6730 11376 11630
rect 11440 8566 11468 13382
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12084 12986 12112 13262
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12544 12714 12572 13194
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12214 12540 12522 12560
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12464 12522 12484
rect 12636 12442 12664 13194
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12728 12374 12756 13262
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11900 11150 11928 11630
rect 12214 11452 12522 11472
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11376 12522 11396
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11532 10674 11560 11086
rect 11900 10810 11928 11086
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 11532 9994 11560 10610
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 10130 11744 10406
rect 11808 10198 11836 10610
rect 12214 10364 12522 10384
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10288 12522 10308
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 12636 10062 12664 10610
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11532 8634 11560 8910
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11532 7954 11560 8570
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11900 8022 11928 8434
rect 11992 8430 12020 9386
rect 12084 8906 12112 9522
rect 12214 9276 12522 9296
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9200 12522 9220
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12544 8566 12572 9046
rect 12636 8634 12664 9998
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 8974 12756 9454
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12544 8378 12572 8502
rect 11992 8090 12020 8366
rect 12544 8350 12664 8378
rect 12214 8188 12522 8208
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8112 12522 8132
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11992 7886 12020 8026
rect 12636 8022 12664 8350
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11992 7546 12020 7822
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11992 7342 12020 7482
rect 11980 7336 12032 7342
rect 11900 7296 11980 7324
rect 11900 6866 11928 7296
rect 11980 7278 12032 7284
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11428 6656 11480 6662
rect 11520 6656 11572 6662
rect 11428 6598 11480 6604
rect 11518 6624 11520 6633
rect 11572 6624 11574 6633
rect 11440 5817 11468 6598
rect 11518 6559 11574 6568
rect 11532 6458 11560 6559
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11900 6390 11928 6802
rect 11992 6798 12020 7142
rect 12214 7100 12522 7120
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7024 12522 7044
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11426 5808 11482 5817
rect 11426 5743 11482 5752
rect 11716 5710 11744 6258
rect 11992 6254 12020 6734
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 12084 5846 12112 6258
rect 12214 6012 12522 6032
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5936 12522 5956
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11716 5370 11744 5646
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 12728 5234 12756 7686
rect 12820 7410 12848 13382
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 12170 12940 12786
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 13004 11830 13032 12650
rect 13188 12306 13216 13194
rect 13372 12986 13400 13194
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 10810 12940 11630
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 13004 11286 13032 11562
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13004 9654 13032 11222
rect 13188 11150 13216 11494
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13188 10826 13216 11086
rect 13188 10798 13308 10826
rect 13280 10742 13308 10798
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13096 10198 13124 10678
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13280 10062 13308 10678
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 14200 9926 14228 14200
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9042 13124 9318
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12912 6798 12940 8298
rect 13096 7954 13124 8774
rect 13280 8430 13308 8910
rect 13268 8424 13320 8430
rect 13266 8392 13268 8401
rect 13320 8392 13322 8401
rect 13266 8327 13322 8336
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 8090 13216 8230
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 14002 7440 14058 7449
rect 13176 7404 13228 7410
rect 14002 7375 14004 7384
rect 13176 7346 13228 7352
rect 14056 7375 14058 7384
rect 14004 7346 14056 7352
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12912 6390 12940 6734
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5914 12848 6190
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12912 5710 12940 6326
rect 13188 5846 13216 7346
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13280 5914 13308 7210
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13372 6390 13400 6666
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 11532 4758 11560 5170
rect 12214 4924 12522 4944
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4848 12522 4868
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 12728 4690 12756 5170
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 13004 4554 13032 5510
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 13096 4758 13124 5034
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 13096 4214 13124 4694
rect 13188 4690 13216 5578
rect 13464 5234 13492 6054
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13464 4622 13492 5170
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11242 3904 11298 3913
rect 11242 3839 11298 3848
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11164 3194 11192 3470
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11440 2990 11468 3946
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11900 3058 11928 3538
rect 11992 3534 12020 4014
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 3194 12020 3470
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12084 3126 12112 3878
rect 12214 3836 12522 3856
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3760 12522 3780
rect 12820 3602 12848 4082
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 13188 3534 13216 3878
rect 13280 3670 13308 3946
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10796 2502 11008 2530
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10520 2106 10640 2122
rect 10520 2100 10652 2106
rect 10520 2094 10600 2100
rect 10600 2042 10652 2048
rect 10704 1902 10732 2450
rect 10692 1896 10744 1902
rect 10692 1838 10744 1844
rect 10704 1426 10732 1838
rect 10692 1420 10744 1426
rect 10692 1362 10744 1368
rect 10048 1158 10100 1164
rect 9692 1018 9720 1158
rect 10244 1142 10456 1170
rect 9680 1012 9732 1018
rect 9680 954 9732 960
rect 8404 870 8616 898
rect 8404 800 8432 870
rect 10244 800 10272 1142
rect 10796 1018 10824 2502
rect 11716 2446 11744 2790
rect 12084 2514 12112 2858
rect 12214 2748 12522 2768
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2672 12522 2692
rect 12728 2582 12756 2926
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10888 2145 10916 2246
rect 10874 2136 10930 2145
rect 10874 2071 10930 2080
rect 10876 2032 10928 2038
rect 10876 1974 10928 1980
rect 10888 1766 10916 1974
rect 10980 1834 11008 2382
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 10968 1828 11020 1834
rect 10968 1770 11020 1776
rect 10876 1760 10928 1766
rect 10876 1702 10928 1708
rect 10888 1358 10916 1702
rect 10876 1352 10928 1358
rect 10980 1329 11008 1770
rect 11532 1426 11560 1906
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 10876 1294 10928 1300
rect 10966 1320 11022 1329
rect 12084 1306 12112 2450
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12214 1660 12522 1680
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1584 12522 1604
rect 12636 1358 12664 2246
rect 12728 2038 12756 2518
rect 13280 2446 13308 3606
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 12716 2032 12768 2038
rect 12716 1974 12768 1980
rect 13096 1358 13124 2314
rect 13188 2106 13216 2314
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13372 1970 13400 2246
rect 13360 1964 13412 1970
rect 13360 1906 13412 1912
rect 13372 1358 13400 1906
rect 12624 1352 12676 1358
rect 12084 1278 12204 1306
rect 12624 1294 12676 1300
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 10966 1255 11022 1264
rect 10784 1012 10836 1018
rect 10784 954 10836 960
rect 12176 800 12204 1278
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 14016 800 14044 1158
rect 4724 734 5028 762
rect 6550 0 6606 800
rect 8390 0 8446 800
rect 10230 0 10286 800
rect 12162 0 12218 800
rect 13912 536 13964 542
rect 13910 504 13912 513
rect 13964 504 13966 513
rect 13910 439 13966 448
rect 14002 0 14058 800
<< via2 >>
rect 10874 14456 10930 14512
rect 1490 11192 1546 11248
rect 754 10512 810 10568
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3606 11092 3608 11112
rect 3608 11092 3660 11112
rect 3660 11092 3662 11112
rect 3606 11056 3662 11092
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4158 11070 4160 11112
rect 4160 11070 4212 11112
rect 4212 11070 4214 11112
rect 4158 11056 4214 11070
rect 4894 11076 4950 11112
rect 4894 11056 4896 11076
rect 4896 11056 4948 11076
rect 4948 11056 4950 11076
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4802 10104 4858 10160
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 5170 10104 5226 10160
rect 5262 10004 5264 10024
rect 5264 10004 5316 10024
rect 5316 10004 5318 10024
rect 5262 9968 5318 10004
rect 5814 10104 5870 10160
rect 6274 11056 6330 11112
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 6642 10512 6698 10568
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1582 3712 1638 3768
rect 3422 4120 3478 4176
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3882 3052 3938 3088
rect 3882 3032 3884 3052
rect 3884 3032 3936 3052
rect 3936 3032 3938 3052
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 7378 11092 7380 11112
rect 7380 11092 7432 11112
rect 7432 11092 7434 11112
rect 7378 11056 7434 11092
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8022 9968 8078 10024
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 7010 6432 7066 6488
rect 6274 6160 6330 6216
rect 5354 4120 5410 4176
rect 5630 4120 5686 4176
rect 6090 4936 6146 4992
rect 5906 3984 5962 4040
rect 6274 3576 6330 3632
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 6090 3032 6146 3088
rect 7194 5652 7196 5672
rect 7196 5652 7248 5672
rect 7248 5652 7250 5672
rect 7194 5616 7250 5652
rect 6642 4120 6698 4176
rect 8022 6452 8078 6488
rect 8022 6432 8024 6452
rect 8024 6432 8076 6452
rect 8076 6432 8078 6452
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 7654 6024 7710 6080
rect 7562 5072 7618 5128
rect 8574 5888 8630 5944
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 9034 6196 9036 6216
rect 9036 6196 9088 6216
rect 9088 6196 9090 6216
rect 9034 6160 9090 6196
rect 9678 10920 9734 10976
rect 10506 13368 10562 13424
rect 10138 12688 10194 12744
rect 9954 11872 10010 11928
rect 10414 10140 10416 10160
rect 10416 10140 10468 10160
rect 10468 10140 10470 10160
rect 10414 10104 10470 10140
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 10690 9016 10746 9072
rect 9126 6060 9128 6080
rect 9128 6060 9180 6080
rect 9180 6060 9182 6080
rect 9126 6024 9182 6060
rect 9494 5908 9550 5944
rect 9494 5888 9496 5908
rect 9496 5888 9548 5908
rect 9548 5888 9550 5908
rect 9678 5908 9734 5944
rect 9678 5888 9680 5908
rect 9680 5888 9732 5908
rect 9732 5888 9734 5908
rect 9586 5752 9642 5808
rect 9218 5652 9220 5672
rect 9220 5652 9272 5672
rect 9272 5652 9274 5672
rect 9218 5616 9274 5652
rect 8758 5480 8814 5536
rect 8298 3984 8354 4040
rect 8298 3476 8300 3496
rect 8300 3476 8352 3496
rect 8352 3476 8354 3496
rect 8298 3440 8354 3476
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 8942 4820 8998 4856
rect 8942 4800 8944 4820
rect 8944 4800 8996 4820
rect 8996 4800 8998 4820
rect 9402 5616 9458 5672
rect 9310 5072 9366 5128
rect 9494 5480 9550 5536
rect 9678 5296 9734 5298
rect 9678 5244 9680 5296
rect 9680 5244 9732 5296
rect 9732 5244 9734 5296
rect 9678 5242 9734 5244
rect 9586 5108 9588 5128
rect 9588 5108 9640 5128
rect 9640 5108 9642 5128
rect 9586 5072 9642 5108
rect 9586 4972 9588 4992
rect 9588 4972 9640 4992
rect 9640 4972 9642 4992
rect 9586 4936 9642 4972
rect 9770 4972 9772 4992
rect 9772 4972 9824 4992
rect 9824 4972 9826 4992
rect 9770 4936 9826 4972
rect 10046 4936 10102 4992
rect 9954 4800 10010 4856
rect 9770 4664 9826 4720
rect 9218 4392 9274 4448
rect 9402 4256 9458 4312
rect 8850 3984 8906 4040
rect 8666 3576 8722 3632
rect 9586 4392 9642 4448
rect 9862 4120 9918 4176
rect 9678 3848 9734 3904
rect 9586 3440 9642 3496
rect 9862 3068 9864 3088
rect 9864 3068 9916 3088
rect 9916 3068 9918 3088
rect 9862 3032 9918 3068
rect 10322 4120 10378 4176
rect 10966 5616 11022 5672
rect 10966 5480 11022 5536
rect 10874 5072 10930 5128
rect 11058 4800 11114 4856
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 11518 6604 11520 6624
rect 11520 6604 11572 6624
rect 11572 6604 11574 6624
rect 11518 6568 11574 6604
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 11426 5752 11482 5808
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 13266 8372 13268 8392
rect 13268 8372 13320 8392
rect 13320 8372 13322 8392
rect 13266 8336 13322 8372
rect 14002 7404 14058 7440
rect 14002 7384 14004 7404
rect 14004 7384 14056 7404
rect 14056 7384 14058 7404
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 11242 3848 11298 3904
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 10874 2080 10930 2136
rect 10966 1264 11022 1320
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 13910 484 13912 504
rect 13912 484 13964 504
rect 13964 484 13966 504
rect 13910 448 13966 484
<< metal3 >>
rect 10869 14514 10935 14517
rect 14200 14514 15000 14544
rect 10869 14512 15000 14514
rect 10869 14456 10874 14512
rect 10930 14456 15000 14512
rect 10869 14454 15000 14456
rect 10869 14451 10935 14454
rect 14200 14424 15000 14454
rect 14200 13698 15000 13728
rect 12758 13638 15000 13698
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 12208 13632 12528 13633
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 13567 12528 13568
rect 10501 13426 10567 13429
rect 12758 13426 12818 13638
rect 14200 13608 15000 13638
rect 10501 13424 12818 13426
rect 10501 13368 10506 13424
rect 10562 13368 12818 13424
rect 10501 13366 12818 13368
rect 10501 13363 10567 13366
rect 8208 13088 8528 13089
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 13023 8528 13024
rect 10133 12746 10199 12749
rect 14200 12746 15000 12776
rect 10133 12744 15000 12746
rect 10133 12688 10138 12744
rect 10194 12688 15000 12744
rect 10133 12686 15000 12688
rect 10133 12683 10199 12686
rect 14200 12656 15000 12686
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 12208 12544 12528 12545
rect 12208 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12528 12544
rect 12208 12479 12528 12480
rect 8208 12000 8528 12001
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 11935 8528 11936
rect 9949 11930 10015 11933
rect 14200 11930 15000 11960
rect 9949 11928 15000 11930
rect 9949 11872 9954 11928
rect 10010 11872 15000 11928
rect 9949 11870 15000 11872
rect 9949 11867 10015 11870
rect 14200 11840 15000 11870
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 12208 11456 12528 11457
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 11391 12528 11392
rect 0 11250 800 11280
rect 1485 11250 1551 11253
rect 0 11248 1551 11250
rect 0 11192 1490 11248
rect 1546 11192 1551 11248
rect 0 11190 1551 11192
rect 0 11160 800 11190
rect 1485 11187 1551 11190
rect 3601 11114 3667 11117
rect 4153 11114 4219 11117
rect 3601 11112 4219 11114
rect 3601 11056 3606 11112
rect 3662 11056 4158 11112
rect 4214 11056 4219 11112
rect 3601 11054 4219 11056
rect 3601 11051 3667 11054
rect 4153 11051 4219 11054
rect 4889 11114 4955 11117
rect 6269 11114 6335 11117
rect 7373 11114 7439 11117
rect 4889 11112 7439 11114
rect 4889 11056 4894 11112
rect 4950 11056 6274 11112
rect 6330 11056 7378 11112
rect 7434 11056 7439 11112
rect 4889 11054 7439 11056
rect 4889 11051 4955 11054
rect 6269 11051 6335 11054
rect 7373 11051 7439 11054
rect 9673 10978 9739 10981
rect 14200 10978 15000 11008
rect 9673 10976 15000 10978
rect 9673 10920 9678 10976
rect 9734 10920 15000 10976
rect 9673 10918 15000 10920
rect 9673 10915 9739 10918
rect 8208 10912 8528 10913
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 14200 10888 15000 10918
rect 8208 10847 8528 10848
rect 749 10570 815 10573
rect 6637 10570 6703 10573
rect 749 10568 6703 10570
rect 749 10512 754 10568
rect 810 10512 6642 10568
rect 6698 10512 6703 10568
rect 749 10510 6703 10512
rect 749 10507 815 10510
rect 6637 10507 6703 10510
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 12208 10368 12528 10369
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 10303 12528 10304
rect 4797 10162 4863 10165
rect 5165 10162 5231 10165
rect 5809 10162 5875 10165
rect 4797 10160 5875 10162
rect 4797 10104 4802 10160
rect 4858 10104 5170 10160
rect 5226 10104 5814 10160
rect 5870 10104 5875 10160
rect 4797 10102 5875 10104
rect 4797 10099 4863 10102
rect 5165 10099 5231 10102
rect 5809 10099 5875 10102
rect 10409 10162 10475 10165
rect 14200 10162 15000 10192
rect 10409 10160 15000 10162
rect 10409 10104 10414 10160
rect 10470 10104 15000 10160
rect 10409 10102 15000 10104
rect 10409 10099 10475 10102
rect 14200 10072 15000 10102
rect 5257 10026 5323 10029
rect 8017 10026 8083 10029
rect 5257 10024 8083 10026
rect 5257 9968 5262 10024
rect 5318 9968 8022 10024
rect 8078 9968 8083 10024
rect 5257 9966 8083 9968
rect 5257 9963 5323 9966
rect 8017 9963 8083 9966
rect 8208 9824 8528 9825
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 9759 8528 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 12208 9280 12528 9281
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 9215 12528 9216
rect 14200 9210 15000 9240
rect 12758 9150 15000 9210
rect 10685 9074 10751 9077
rect 12758 9074 12818 9150
rect 14200 9120 15000 9150
rect 10685 9072 12818 9074
rect 10685 9016 10690 9072
rect 10746 9016 12818 9072
rect 10685 9014 12818 9016
rect 10685 9011 10751 9014
rect 8208 8736 8528 8737
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8671 8528 8672
rect 13261 8394 13327 8397
rect 14200 8394 15000 8424
rect 13261 8392 15000 8394
rect 13261 8336 13266 8392
rect 13322 8336 15000 8392
rect 13261 8334 15000 8336
rect 13261 8331 13327 8334
rect 14200 8304 15000 8334
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 12208 8192 12528 8193
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 8127 12528 8128
rect 8208 7648 8528 7649
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 7583 8528 7584
rect 13997 7442 14063 7445
rect 14200 7442 15000 7472
rect 13997 7440 15000 7442
rect 13997 7384 14002 7440
rect 14058 7384 15000 7440
rect 13997 7382 15000 7384
rect 13997 7379 14063 7382
rect 14200 7352 15000 7382
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 12208 7104 12528 7105
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 7039 12528 7040
rect 11513 6626 11579 6629
rect 14200 6626 15000 6656
rect 11513 6624 15000 6626
rect 11513 6568 11518 6624
rect 11574 6568 15000 6624
rect 11513 6566 15000 6568
rect 11513 6563 11579 6566
rect 8208 6560 8528 6561
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 14200 6536 15000 6566
rect 8208 6495 8528 6496
rect 7005 6490 7071 6493
rect 8017 6490 8083 6493
rect 7005 6488 8083 6490
rect 7005 6432 7010 6488
rect 7066 6432 8022 6488
rect 8078 6432 8083 6488
rect 7005 6430 8083 6432
rect 7005 6427 7071 6430
rect 8017 6427 8083 6430
rect 6269 6218 6335 6221
rect 9029 6218 9095 6221
rect 6269 6216 9095 6218
rect 6269 6160 6274 6216
rect 6330 6160 9034 6216
rect 9090 6160 9095 6216
rect 6269 6158 9095 6160
rect 6269 6155 6335 6158
rect 9029 6155 9095 6158
rect 7649 6082 7715 6085
rect 9121 6084 9187 6085
rect 9070 6082 9076 6084
rect 7649 6080 9076 6082
rect 9140 6082 9187 6084
rect 9140 6080 9232 6082
rect 7649 6024 7654 6080
rect 7710 6024 9076 6080
rect 9182 6024 9232 6080
rect 7649 6022 9076 6024
rect 7649 6019 7715 6022
rect 9070 6020 9076 6022
rect 9140 6022 9232 6024
rect 9140 6020 9187 6022
rect 9121 6019 9187 6020
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 12208 6016 12528 6017
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 5951 12528 5952
rect 8569 5946 8635 5949
rect 9489 5946 9555 5949
rect 8569 5944 9555 5946
rect 8569 5888 8574 5944
rect 8630 5888 9494 5944
rect 9550 5888 9555 5944
rect 8569 5886 9555 5888
rect 8569 5883 8635 5886
rect 9489 5883 9555 5886
rect 9673 5946 9739 5949
rect 9806 5946 9812 5948
rect 9673 5944 9812 5946
rect 9673 5888 9678 5944
rect 9734 5888 9812 5944
rect 9673 5886 9812 5888
rect 9673 5883 9739 5886
rect 9806 5884 9812 5886
rect 9876 5884 9882 5948
rect 9438 5748 9444 5812
rect 9508 5810 9514 5812
rect 9581 5810 9647 5813
rect 11421 5810 11487 5813
rect 9508 5808 9647 5810
rect 9508 5752 9586 5808
rect 9642 5752 9647 5808
rect 9508 5750 9647 5752
rect 9508 5748 9514 5750
rect 9581 5747 9647 5750
rect 9768 5808 11487 5810
rect 9768 5752 11426 5808
rect 11482 5752 11487 5808
rect 9768 5750 11487 5752
rect 7189 5674 7255 5677
rect 9213 5676 9279 5677
rect 9213 5674 9260 5676
rect 7189 5672 9260 5674
rect 7189 5616 7194 5672
rect 7250 5616 9218 5672
rect 7189 5614 9260 5616
rect 7189 5611 7255 5614
rect 9213 5612 9260 5614
rect 9324 5612 9330 5676
rect 9397 5674 9463 5677
rect 9768 5674 9828 5750
rect 11421 5747 11487 5750
rect 9397 5672 9828 5674
rect 9397 5616 9402 5672
rect 9458 5616 9828 5672
rect 9397 5614 9828 5616
rect 10961 5674 11027 5677
rect 14200 5674 15000 5704
rect 10961 5672 15000 5674
rect 10961 5616 10966 5672
rect 11022 5616 15000 5672
rect 10961 5614 15000 5616
rect 9213 5611 9279 5612
rect 9397 5611 9463 5614
rect 10961 5611 11027 5614
rect 14200 5584 15000 5614
rect 8753 5538 8819 5541
rect 9489 5538 9555 5541
rect 10961 5538 11027 5541
rect 8753 5536 9555 5538
rect 8753 5480 8758 5536
rect 8814 5480 9494 5536
rect 9550 5480 9555 5536
rect 8753 5478 9555 5480
rect 8753 5475 8819 5478
rect 9489 5475 9555 5478
rect 9630 5536 11027 5538
rect 9630 5480 10966 5536
rect 11022 5480 11027 5536
rect 9630 5478 11027 5480
rect 8208 5472 8528 5473
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 5407 8528 5408
rect 9630 5303 9690 5478
rect 10961 5475 11027 5478
rect 9630 5298 9739 5303
rect 9630 5242 9678 5298
rect 9734 5242 9739 5298
rect 9630 5240 9739 5242
rect 9673 5237 9739 5240
rect 7557 5130 7623 5133
rect 9305 5130 9371 5133
rect 9581 5130 9647 5133
rect 7557 5128 9371 5130
rect 7557 5072 7562 5128
rect 7618 5072 9310 5128
rect 9366 5072 9371 5128
rect 7557 5070 9371 5072
rect 7557 5067 7623 5070
rect 9305 5067 9371 5070
rect 9446 5128 9647 5130
rect 9446 5072 9586 5128
rect 9642 5072 9647 5128
rect 9446 5070 9647 5072
rect 6085 4994 6151 4997
rect 9446 4994 9506 5070
rect 9581 5067 9647 5070
rect 10869 5130 10935 5133
rect 10869 5128 12818 5130
rect 10869 5072 10874 5128
rect 10930 5072 12818 5128
rect 10869 5070 12818 5072
rect 10869 5067 10935 5070
rect 6085 4992 9506 4994
rect 6085 4936 6090 4992
rect 6146 4936 9506 4992
rect 6085 4934 9506 4936
rect 9581 4994 9647 4997
rect 9765 4994 9831 4997
rect 10041 4994 10107 4997
rect 9581 4992 9690 4994
rect 9581 4936 9586 4992
rect 9642 4936 9690 4992
rect 6085 4931 6151 4934
rect 9581 4931 9690 4936
rect 9765 4992 10107 4994
rect 9765 4936 9770 4992
rect 9826 4936 10046 4992
rect 10102 4936 10107 4992
rect 9765 4934 10107 4936
rect 9765 4931 9831 4934
rect 10041 4931 10107 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 8937 4858 9003 4861
rect 9630 4858 9690 4931
rect 12208 4928 12528 4929
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4863 12528 4864
rect 8937 4856 9690 4858
rect 8937 4800 8942 4856
rect 8998 4800 9690 4856
rect 8937 4798 9690 4800
rect 9949 4858 10015 4861
rect 11053 4858 11119 4861
rect 9949 4856 11119 4858
rect 9949 4800 9954 4856
rect 10010 4800 11058 4856
rect 11114 4800 11119 4856
rect 9949 4798 11119 4800
rect 12758 4858 12818 5070
rect 14200 4858 15000 4888
rect 12758 4798 15000 4858
rect 8937 4795 9003 4798
rect 9949 4795 10015 4798
rect 11053 4795 11119 4798
rect 14200 4768 15000 4798
rect 9765 4724 9831 4725
rect 9765 4720 9812 4724
rect 9876 4722 9882 4724
rect 9765 4664 9770 4720
rect 9765 4660 9812 4664
rect 9876 4662 9922 4722
rect 9876 4660 9882 4662
rect 9765 4659 9831 4660
rect 9070 4388 9076 4452
rect 9140 4450 9146 4452
rect 9213 4450 9279 4453
rect 9140 4448 9279 4450
rect 9140 4392 9218 4448
rect 9274 4392 9279 4448
rect 9140 4390 9279 4392
rect 9140 4388 9146 4390
rect 9213 4387 9279 4390
rect 9438 4388 9444 4452
rect 9508 4450 9514 4452
rect 9581 4450 9647 4453
rect 9508 4448 9647 4450
rect 9508 4392 9586 4448
rect 9642 4392 9647 4448
rect 9508 4390 9647 4392
rect 9508 4388 9514 4390
rect 9581 4387 9647 4390
rect 8208 4384 8528 4385
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 4319 8528 4320
rect 9254 4252 9260 4316
rect 9324 4314 9330 4316
rect 9397 4314 9463 4317
rect 9324 4312 9463 4314
rect 9324 4256 9402 4312
rect 9458 4256 9463 4312
rect 9324 4254 9463 4256
rect 9324 4252 9330 4254
rect 9397 4251 9463 4254
rect 3417 4178 3483 4181
rect 5349 4178 5415 4181
rect 5625 4178 5691 4181
rect 6637 4178 6703 4181
rect 3417 4176 6703 4178
rect 3417 4120 3422 4176
rect 3478 4120 5354 4176
rect 5410 4120 5630 4176
rect 5686 4120 6642 4176
rect 6698 4120 6703 4176
rect 3417 4118 6703 4120
rect 3417 4115 3483 4118
rect 5349 4115 5415 4118
rect 5625 4115 5691 4118
rect 6637 4115 6703 4118
rect 9857 4178 9923 4181
rect 10317 4178 10383 4181
rect 9857 4176 10383 4178
rect 9857 4120 9862 4176
rect 9918 4120 10322 4176
rect 10378 4120 10383 4176
rect 9857 4118 10383 4120
rect 9857 4115 9923 4118
rect 10317 4115 10383 4118
rect 5901 4042 5967 4045
rect 8293 4042 8359 4045
rect 5901 4040 8359 4042
rect 5901 3984 5906 4040
rect 5962 3984 8298 4040
rect 8354 3984 8359 4040
rect 5901 3982 8359 3984
rect 5901 3979 5967 3982
rect 8293 3979 8359 3982
rect 8845 4042 8911 4045
rect 8845 4040 12818 4042
rect 8845 3984 8850 4040
rect 8906 3984 12818 4040
rect 8845 3982 12818 3984
rect 8845 3979 8911 3982
rect 9673 3906 9739 3909
rect 11237 3906 11303 3909
rect 9673 3904 11303 3906
rect 9673 3848 9678 3904
rect 9734 3848 11242 3904
rect 11298 3848 11303 3904
rect 9673 3846 11303 3848
rect 12758 3906 12818 3982
rect 14200 3906 15000 3936
rect 12758 3846 15000 3906
rect 9673 3843 9739 3846
rect 11237 3843 11303 3846
rect 4208 3840 4528 3841
rect 0 3770 800 3800
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 12208 3840 12528 3841
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 14200 3816 15000 3846
rect 12208 3775 12528 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 6269 3634 6335 3637
rect 8661 3634 8727 3637
rect 6269 3632 8727 3634
rect 6269 3576 6274 3632
rect 6330 3576 8666 3632
rect 8722 3576 8727 3632
rect 6269 3574 8727 3576
rect 6269 3571 6335 3574
rect 8661 3571 8727 3574
rect 8293 3498 8359 3501
rect 9581 3498 9647 3501
rect 8293 3496 9647 3498
rect 8293 3440 8298 3496
rect 8354 3440 9586 3496
rect 9642 3440 9647 3496
rect 8293 3438 9647 3440
rect 8293 3435 8359 3438
rect 9581 3435 9647 3438
rect 8208 3296 8528 3297
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 3231 8528 3232
rect 3877 3090 3943 3093
rect 6085 3090 6151 3093
rect 3877 3088 6151 3090
rect 3877 3032 3882 3088
rect 3938 3032 6090 3088
rect 6146 3032 6151 3088
rect 3877 3030 6151 3032
rect 3877 3027 3943 3030
rect 6085 3027 6151 3030
rect 9857 3090 9923 3093
rect 14200 3090 15000 3120
rect 9857 3088 15000 3090
rect 9857 3032 9862 3088
rect 9918 3032 15000 3088
rect 9857 3030 15000 3032
rect 9857 3027 9923 3030
rect 14200 3000 15000 3030
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 12208 2752 12528 2753
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 2687 12528 2688
rect 8208 2208 8528 2209
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 2143 8528 2144
rect 10869 2138 10935 2141
rect 14200 2138 15000 2168
rect 10869 2136 15000 2138
rect 10869 2080 10874 2136
rect 10930 2080 15000 2136
rect 10869 2078 15000 2080
rect 10869 2075 10935 2078
rect 14200 2048 15000 2078
rect 4208 1664 4528 1665
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1599 4528 1600
rect 12208 1664 12528 1665
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1599 12528 1600
rect 10961 1322 11027 1325
rect 14200 1322 15000 1352
rect 10961 1320 15000 1322
rect 10961 1264 10966 1320
rect 11022 1264 15000 1320
rect 10961 1262 15000 1264
rect 10961 1259 11027 1262
rect 14200 1232 15000 1262
rect 8208 1120 8528 1121
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1055 8528 1056
rect 13905 506 13971 509
rect 14200 506 15000 536
rect 13905 504 15000 506
rect 13905 448 13910 504
rect 13966 448 15000 504
rect 13905 446 15000 448
rect 13905 443 13971 446
rect 14200 416 15000 446
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 9076 6080 9140 6084
rect 9076 6024 9126 6080
rect 9126 6024 9140 6080
rect 9076 6020 9140 6024
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 9812 5884 9876 5948
rect 9444 5748 9508 5812
rect 9260 5672 9324 5676
rect 9260 5616 9274 5672
rect 9274 5616 9324 5672
rect 9260 5612 9324 5616
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 9812 4720 9876 4724
rect 9812 4664 9826 4720
rect 9826 4664 9876 4720
rect 9812 4660 9876 4664
rect 9076 4388 9140 4452
rect 9444 4388 9508 4452
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 9260 4252 9324 4316
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 9075 6084 9141 6085
rect 9075 6020 9076 6084
rect 9140 6020 9141 6084
rect 9075 6019 9141 6020
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 9078 4453 9138 6019
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 9811 5948 9877 5949
rect 9811 5884 9812 5948
rect 9876 5884 9877 5948
rect 9811 5883 9877 5884
rect 9443 5812 9509 5813
rect 9443 5748 9444 5812
rect 9508 5748 9509 5812
rect 9443 5747 9509 5748
rect 9259 5676 9325 5677
rect 9259 5612 9260 5676
rect 9324 5612 9325 5676
rect 9259 5611 9325 5612
rect 9075 4452 9141 4453
rect 9075 4388 9076 4452
rect 9140 4388 9141 4452
rect 9075 4387 9141 4388
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 9262 4317 9322 5611
rect 9446 4453 9506 5747
rect 9814 4725 9874 5883
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 9811 4724 9877 4725
rect 9811 4660 9812 4724
rect 9876 4660 9877 4724
rect 9811 4659 9877 4660
rect 12208 4488 12528 4864
rect 9443 4452 9509 4453
rect 9443 4388 9444 4452
rect 9508 4388 9509 4452
rect 9443 4387 9509 4388
rect 9259 4316 9325 4317
rect 9259 4252 9260 4316
rect 9324 4252 9325 4316
rect 9259 4251 9325 4252
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 4250 4252 4486 4488
rect 8250 8252 8486 8488
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 12250 4252 12486 4488
<< metal5 >>
rect 1104 12488 13892 12530
rect 1104 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 13892 12488
rect 1104 12210 13892 12252
rect 1104 8488 13892 8530
rect 1104 8252 8250 8488
rect 8486 8252 13892 8488
rect 1104 8210 13892 8252
rect 1104 4488 13892 4530
rect 1104 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 13892 4488
rect 1104 4210 13892 4252
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 2300 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 2484 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1380 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1932 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635271187
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _333_
timestamp 1635271187
transform 1 0 2024 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _364_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1380 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1635271187
transform 1 0 3128 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__D
timestamp 1635271187
transform -1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _365_
timestamp 1635271187
transform 1 0 3312 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _366_
timestamp 1635271187
transform -1 0 5704 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1635271187
transform 1 0 5704 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1635271187
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1635271187
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6992 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6348 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5244 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6348 0 -1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1635271187
transform 1 0 8464 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__B
timestamp 1635271187
transform -1 0 8832 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1635271187
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7268 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 7912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8188 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8188 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1635271187
transform 1 0 8924 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7912 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A1
timestamp 1635271187
transform -1 0 11132 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__S
timestamp 1635271187
transform -1 0 11316 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 11408 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1635271187
transform 1 0 9844 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1635271187
transform 1 0 10672 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1635271187
transform 1 0 9568 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1635271187
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1635271187
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1635271187
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1635271187
transform 1 0 13156 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1635271187
transform 1 0 11500 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1635271187
transform 1 0 11500 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1635271187
transform 1 0 12420 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1635271187
transform -1 0 12420 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__S
timestamp 1635271187
transform 1 0 13432 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1635271187
transform 1 0 13432 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635271187
transform -1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635271187
transform -1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1635271187
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635271187
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _321_
timestamp 1635271187
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A
timestamp 1635271187
transform 1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A
timestamp 1635271187
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1635271187
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_24
timestamp 1635271187
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1635271187
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 4692 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _319_
timestamp 1635271187
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _331_
timestamp 1635271187
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_44
timestamp 1635271187
transform 1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0
timestamp 1635271187
transform 1 0 5704 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1635271187
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__S
timestamp 1635271187
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1635271187
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1635271187
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7360 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1635271187
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7820 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A1
timestamp 1635271187
transform -1 0 10948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__S
timestamp 1635271187
transform 1 0 10948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1635271187
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_109
timestamp 1635271187
transform 1 0 11132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _334_
timestamp 1635271187
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1635271187
transform 1 0 9752 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A1
timestamp 1635271187
transform -1 0 11776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__S
timestamp 1635271187
transform 1 0 11408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__S
timestamp 1635271187
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1635271187
transform -1 0 12604 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1635271187
transform 1 0 12604 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635271187
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1635271187
transform -1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1635271187
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_8
timestamp 1635271187
transform 1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635271187
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _376_
timestamp 1635271187
transform 1 0 2024 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _378_
timestamp 1635271187
transform 1 0 3956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1635271187
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1635271187
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp 1635271187
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1635271187
transform 1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A1
timestamp 1635271187
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__S
timestamp 1635271187
transform 1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A1
timestamp 1635271187
transform -1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1635271187
transform 1 0 8464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_85
timestamp 1635271187
transform 1 0 8924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1635271187
transform 1 0 7636 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1635271187
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _236_
timestamp 1635271187
transform 1 0 9936 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1635271187
transform -1 0 11224 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A1
timestamp 1635271187
transform -1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__S
timestamp 1635271187
transform 1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A1
timestamp 1635271187
transform -1 0 11408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1635271187
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1635271187
transform 1 0 12144 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1635271187
transform 1 0 11500 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A1
timestamp 1635271187
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_135
timestamp 1635271187
transform 1 0 13524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635271187
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1635271187
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635271187
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _374_
timestamp 1635271187
transform 1 0 1472 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1635271187
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1635271187
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1635271187
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4324 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1635271187
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp 1635271187
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _255_
timestamp 1635271187
transform -1 0 5796 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _375_
timestamp 1635271187
transform 1 0 6256 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1635271187
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8188 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1635271187
transform -1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _286_
timestamp 1635271187
transform -1 0 10948 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _290_
timestamp 1635271187
transform 1 0 9752 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1635271187
transform 1 0 10948 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1635271187
transform 1 0 11960 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635271187
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A
timestamp 1635271187
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_11
timestamp 1635271187
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635271187
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 2668 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp 1635271187
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_26
timestamp 1635271187
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1635271187
transform 1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4232 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _264_
timestamp 1635271187
transform -1 0 4232 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1635271187
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _247_
timestamp 1635271187
transform -1 0 6992 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1635271187
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _266_
timestamp 1635271187
transform 1 0 5152 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _268_
timestamp 1635271187
transform -1 0 7636 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1635271187
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A1
timestamp 1635271187
transform -1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1635271187
transform 1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _322_
timestamp 1635271187
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1635271187
transform -1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_105
timestamp 1635271187
transform 1 0 10764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_109
timestamp 1635271187
transform 1 0 11132 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_89
timestamp 1635271187
transform 1 0 9292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_99
timestamp 1635271187
transform 1 0 10212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1635271187
transform -1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _296_
timestamp 1635271187
transform 1 0 10304 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 9660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__S
timestamp 1635271187
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__S
timestamp 1635271187
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1635271187
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1635271187
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1635271187
transform -1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1635271187
transform -1 0 12144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1635271187
transform 1 0 12144 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1635271187
transform 1 0 12788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1635271187
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635271187
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 1635271187
transform -1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1635271187
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635271187
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635271187
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1635271187
transform -1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _269_
timestamp 1635271187
transform -1 0 3680 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _273_
timestamp 1635271187
transform 1 0 2392 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _325_
timestamp 1635271187
transform 1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _372_
timestamp 1635271187
transform -1 0 3312 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1635271187
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_28
timestamp 1635271187
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_32
timestamp 1635271187
transform 1 0 4048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1635271187
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1635271187
transform 1 0 3772 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _250_
timestamp 1635271187
transform -1 0 5244 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_2  _253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4600 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _259_
timestamp 1635271187
transform 1 0 4140 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_2  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5428 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _246_
timestamp 1635271187
transform -1 0 6256 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1635271187
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_50
timestamp 1635271187
transform 1 0 5704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1635271187
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__o32a_2  _249_
timestamp 1635271187
transform 1 0 6348 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _228_
timestamp 1635271187
transform 1 0 6624 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1635271187
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 1635271187
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_59
timestamp 1635271187
transform 1 0 6532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A1
timestamp 1635271187
transform -1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1635271187
transform 1 0 7452 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_2  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8556 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _234_
timestamp 1635271187
transform 1 0 7176 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1635271187
transform -1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_2  _304_
timestamp 1635271187
transform 1 0 8556 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_2  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 9108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1635271187
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1635271187
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1635271187
transform 1 0 8280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1635271187
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A1
timestamp 1635271187
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A1
timestamp 1635271187
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_105
timestamp 1635271187
transform 1 0 10764 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_91
timestamp 1635271187
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_2  _301_
timestamp 1635271187
transform 1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _312_
timestamp 1635271187
transform 1 0 9936 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1635271187
transform -1 0 11408 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1635271187
transform 1 0 10856 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_6_124
timestamp 1635271187
transform 1 0 12512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1635271187
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _238_
timestamp 1635271187
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1635271187
transform 1 0 12604 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1635271187
transform 1 0 11960 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1635271187
transform 1 0 11500 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_6_135
timestamp 1635271187
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635271187
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635271187
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1635271187
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1635271187
transform 1 0 2392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_16
timestamp 1635271187
transform 1 0 2576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1635271187
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635271187
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _271_
timestamp 1635271187
transform 1 0 2668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _324_
timestamp 1635271187
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_24
timestamp 1635271187
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1635271187
transform 1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1635271187
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1635271187
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4416 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _244_
timestamp 1635271187
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_8_58
timestamp 1635271187
transform 1 0 6440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1635271187
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _230_
timestamp 1635271187
transform -1 0 7360 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _251_
timestamp 1635271187
transform -1 0 5796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _260_
timestamp 1635271187
transform -1 0 6440 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__S
timestamp 1635271187
transform 1 0 8556 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp 1635271187
transform 1 0 7636 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1635271187
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1635271187
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1635271187
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _306_
timestamp 1635271187
transform 1 0 7728 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1635271187
transform -1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _302_
timestamp 1635271187
transform -1 0 10120 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1635271187
transform 1 0 10396 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_122
timestamp 1635271187
transform 1 0 12328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _309_
timestamp 1635271187
transform 1 0 11224 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1635271187
transform 1 0 12420 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1635271187
transform 1 0 11684 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1635271187
transform 1 0 12696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1635271187
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A1
timestamp 1635271187
transform -1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__S
timestamp 1635271187
transform 1 0 13248 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635271187
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635271187
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _373_
timestamp 1635271187
transform 1 0 1380 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_9_42
timestamp 1635271187
transform 1 0 4968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 4968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _262_
timestamp 1635271187
transform 1 0 5060 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_2  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_9_52
timestamp 1635271187
transform 1 0 5888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1635271187
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1635271187
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1635271187
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__S
timestamp 1635271187
transform 1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1635271187
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_80
timestamp 1635271187
transform 1 0 8464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1635271187
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _288_
timestamp 1635271187
transform 1 0 7268 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_2  _295_
timestamp 1635271187
transform -1 0 9660 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1635271187
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__S
timestamp 1635271187
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A1
timestamp 1635271187
transform -1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp 1635271187
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _239_
timestamp 1635271187
transform -1 0 10396 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _300_
timestamp 1635271187
transform 1 0 10396 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A1
timestamp 1635271187
transform -1 0 11408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1635271187
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1635271187
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1635271187
transform 1 0 12604 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1635271187
transform 1 0 11592 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635271187
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1635271187
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1635271187
transform 1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp 1635271187
transform 1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1635271187
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1635271187
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635271187
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _197_
timestamp 1635271187
transform -1 0 2760 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _318_
timestamp 1635271187
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1635271187
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and4_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _240_
timestamp 1635271187
transform -1 0 3680 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _242_
timestamp 1635271187
transform 1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1635271187
transform 1 0 5244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _377_
timestamp 1635271187
transform 1 0 5428 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_10_75
timestamp 1635271187
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1635271187
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1635271187
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_2  _291_
timestamp 1635271187
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1635271187
transform 1 0 7360 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _289_
timestamp 1635271187
transform -1 0 10212 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1635271187
transform -1 0 11040 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1635271187
transform 1 0 11040 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_117
timestamp 1635271187
transform 1 0 11868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1635271187
transform 1 0 11960 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635271187
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635271187
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _379_
timestamp 1635271187
transform 1 0 1380 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1635271187
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1635271187
transform 1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4416 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1635271187
transform 1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_45
timestamp 1635271187
transform 1 0 5244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1635271187
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1635271187
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1635271187
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _263_
timestamp 1635271187
transform 1 0 5336 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _320_
timestamp 1635271187
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1635271187
transform 1 0 8464 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1635271187
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_2  _294_
timestamp 1635271187
transform -1 0 9568 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1635271187
transform 1 0 7176 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1635271187
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 9568 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1635271187
transform -1 0 11408 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A1
timestamp 1635271187
transform -1 0 11960 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__S
timestamp 1635271187
transform 1 0 11592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1635271187
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1635271187
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1635271187
transform 1 0 11960 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1635271187
transform 1 0 12788 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635271187
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635271187
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _380_
timestamp 1635271187
transform -1 0 3312 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_12_24
timestamp 1635271187
transform 1 0 3312 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1635271187
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _316_
timestamp 1635271187
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _381_
timestamp 1635271187
transform -1 0 5704 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A1
timestamp 1635271187
transform 1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1635271187
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_59
timestamp 1635271187
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _226_
timestamp 1635271187
transform 1 0 5704 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1635271187
transform 1 0 7084 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1635271187
transform -1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__S
timestamp 1635271187
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1635271187
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_2  _293_
timestamp 1635271187
transform -1 0 9844 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_2  _297_
timestamp 1635271187
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1635271187
transform 1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_2  _298_
timestamp 1635271187
transform -1 0 10488 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 11224 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1
timestamp 1635271187
transform -1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__S
timestamp 1635271187
transform 1 0 12420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A1
timestamp 1635271187
transform -1 0 11776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__S
timestamp 1635271187
transform 1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1635271187
transform 1 0 11224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1635271187
transform 1 0 12788 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1635271187
transform 1 0 11776 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635271187
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _335_
timestamp 1635271187
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _317_
timestamp 1635271187
transform 1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635271187
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635271187
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1635271187
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1635271187
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1635271187
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 1635271187
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _196_
timestamp 1635271187
transform 1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_15
timestamp 1635271187
transform 1 0 2484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1635271187
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _367_
timestamp 1635271187
transform 1 0 2852 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1635271187
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_40
timestamp 1635271187
transform 1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1635271187
transform 1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_34
timestamp 1635271187
transform 1 0 4232 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_40
timestamp 1635271187
transform 1 0 4784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1635271187
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1635271187
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _330_
timestamp 1635271187
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _382_
timestamp 1635271187
transform 1 0 4876 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp 1635271187
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1635271187
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1635271187
transform 1 0 5520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1635271187
transform 1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1635271187
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1635271187
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1635271187
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_59
timestamp 1635271187
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635271187
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 1635271187
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1635271187
transform 1 0 6992 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1635271187
transform -1 0 8832 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A1
timestamp 1635271187
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__S
timestamp 1635271187
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_76
timestamp 1635271187
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1635271187
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1635271187
transform -1 0 9752 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1635271187
transform 1 0 7452 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1635271187
transform 1 0 8648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_109
timestamp 1635271187
transform 1 0 11132 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_105
timestamp 1635271187
transform 1 0 10764 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_94
timestamp 1635271187
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1635271187
transform 1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1635271187
transform 1 0 9844 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1635271187
transform 1 0 9200 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1635271187
transform 1 0 9844 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1635271187
transform 1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1635271187
transform 1 0 10856 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A1
timestamp 1635271187
transform -1 0 11408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_122
timestamp 1635271187
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1635271187
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1635271187
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1635271187
transform 1 0 12788 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1635271187
transform 1 0 11500 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1635271187
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1635271187
transform 1 0 12420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A1
timestamp 1635271187
transform -1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635271187
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635271187
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635271187
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _386_
timestamp 1635271187
transform 1 0 1380 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_2  _188_
timestamp 1635271187
transform -1 0 4048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _194_
timestamp 1635271187
transform 1 0 4692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _282_
timestamp 1635271187
transform -1 0 4692 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 1635271187
transform 1 0 5796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1635271187
transform 1 0 5428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1635271187
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _314_
timestamp 1635271187
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _383_
timestamp 1635271187
transform 1 0 6348 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_15_86
timestamp 1635271187
transform 1 0 9016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1635271187
transform 1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _223_
timestamp 1635271187
transform 1 0 8280 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1635271187
transform 1 0 9108 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1635271187
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1635271187
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__S
timestamp 1635271187
transform 1 0 12512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1635271187
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1635271187
transform -1 0 13064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1635271187
transform 1 0 13064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1635271187
transform 1 0 11500 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__S
timestamp 1635271187
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1635271187
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635271187
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A
timestamp 1635271187
transform 1 0 2392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_16
timestamp 1635271187
transform 1 0 2576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1635271187
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1635271187
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635271187
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1635271187
transform -1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _329_
timestamp 1635271187
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1635271187
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1635271187
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1635271187
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _219_
timestamp 1635271187
transform 1 0 3956 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__B1
timestamp 1635271187
transform 1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1635271187
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1635271187
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _193_
timestamp 1635271187
transform 1 0 5796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _215_
timestamp 1635271187
transform 1 0 7084 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1635271187
transform 1 0 8188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1635271187
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _201_
timestamp 1635271187
transform 1 0 7728 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _214_
timestamp 1635271187
transform -1 0 8832 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_2  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1635271187
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__S
timestamp 1635271187
transform 1 0 10488 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1635271187
transform -1 0 10304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1635271187
transform 1 0 10672 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_16_122
timestamp 1635271187
transform 1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1635271187
transform -1 0 12328 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1635271187
transform 1 0 12604 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1635271187
transform 1 0 13524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635271187
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1635271187
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635271187
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _368_
timestamp 1635271187
transform 1 0 1380 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_17_36
timestamp 1635271187
transform 1 0 4416 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1635271187
transform 1 0 4140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_2  _283_
timestamp 1635271187
transform 1 0 3312 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1635271187
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_64
timestamp 1635271187
transform 1 0 6992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1635271187
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1635271187
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _213_
timestamp 1635271187
transform -1 0 7912 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _221_
timestamp 1635271187
transform 1 0 5244 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _279_
timestamp 1635271187
transform -1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _217_
timestamp 1635271187
transform 1 0 8556 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7912 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A1
timestamp 1635271187
transform 1 0 9476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__B1
timestamp 1635271187
transform 1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_104
timestamp 1635271187
transform 1 0 10672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_90
timestamp 1635271187
transform 1 0 9384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1635271187
transform -1 0 10488 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1635271187
transform 1 0 10764 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A1
timestamp 1635271187
transform -1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1635271187
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1635271187
transform -1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1635271187
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1635271187
transform 1 0 12512 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1635271187
transform -1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1635271187
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635271187
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_15
timestamp 1635271187
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1635271187
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635271187
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _281_
timestamp 1635271187
transform 1 0 2760 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1635271187
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1635271187
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _277_
timestamp 1635271187
transform 1 0 4508 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1635271187
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_62
timestamp 1635271187
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _203_
timestamp 1635271187
transform -1 0 7636 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _274_
timestamp 1635271187
transform -1 0 6808 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _280_
timestamp 1635271187
transform 1 0 5336 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 1635271187
transform -1 0 8740 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_78
timestamp 1635271187
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1635271187
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1635271187
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _202_
timestamp 1635271187
transform -1 0 8280 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _224_
timestamp 1635271187
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _287_
timestamp 1635271187
transform 1 0 9752 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1635271187
transform 1 0 10212 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1635271187
transform 1 0 11868 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_18_135
timestamp 1635271187
transform 1 0 13524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635271187
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1635271187
transform 1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_21
timestamp 1635271187
transform 1 0 3036 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635271187
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635271187
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _326_
timestamp 1635271187
transform -1 0 2852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _371_
timestamp 1635271187
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1635271187
transform -1 0 2576 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_20_24
timestamp 1635271187
transform 1 0 3312 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1635271187
transform 1 0 4416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1635271187
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _191_
timestamp 1635271187
transform -1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _220_
timestamp 1635271187
transform 1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _276_
timestamp 1635271187
transform -1 0 4416 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _327_
timestamp 1635271187
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _370_
timestamp 1635271187
transform 1 0 3128 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1635271187
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1635271187
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1635271187
transform 1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1635271187
transform -1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _198_
timestamp 1635271187
transform -1 0 6256 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _199_
timestamp 1635271187
transform 1 0 5244 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _204_
timestamp 1635271187
transform 1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_2  _205_
timestamp 1635271187
transform -1 0 6716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _211_
timestamp 1635271187
transform -1 0 8832 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _207_
timestamp 1635271187
transform 1 0 7636 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _206_
timestamp 1635271187
transform 1 0 7452 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_19_70
timestamp 1635271187
transform 1 0 7544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1635271187
transform 1 0 7176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1635271187
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _209_
timestamp 1635271187
transform -1 0 9384 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8924 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1635271187
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_84
timestamp 1635271187
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_78
timestamp 1635271187
transform 1 0 8280 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1635271187
transform -1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A1
timestamp 1635271187
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__B1
timestamp 1635271187
transform 1 0 9844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_93
timestamp 1635271187
transform 1 0 9660 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_99
timestamp 1635271187
transform 1 0 10212 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1635271187
transform 1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1635271187
transform -1 0 10580 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1635271187
transform 1 0 10580 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1635271187
transform 1 0 10304 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1635271187
transform -1 0 12328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1635271187
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1635271187
transform 1 0 11316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1635271187
transform -1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1635271187
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_116
timestamp 1635271187
transform 1 0 11776 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1635271187
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__S
timestamp 1635271187
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A1
timestamp 1635271187
transform -1 0 11408 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1635271187
transform 1 0 12328 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1635271187
transform 1 0 12972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1635271187
transform 1 0 12236 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_19_133
timestamp 1635271187
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1635271187
transform 1 0 13524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635271187
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635271187
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1635271187
transform 1 0 13248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1635271187
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1635271187
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635271187
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _369_
timestamp 1635271187
transform 1 0 2300 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _385_
timestamp 1635271187
transform 1 0 4232 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1635271187
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1635271187
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _384_
timestamp 1635271187
transform 1 0 6348 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_21_81
timestamp 1635271187
transform 1 0 8556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp 1635271187
transform -1 0 8556 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1635271187
transform -1 0 9476 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A1
timestamp 1635271187
transform -1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_93
timestamp 1635271187
transform 1 0 9660 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1635271187
transform 1 0 9752 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1635271187
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1635271187
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1635271187
transform 1 0 11684 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635271187
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1635271187
transform 1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1635271187
transform 1 0 2484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_21
timestamp 1635271187
transform 1 0 3036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1635271187
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635271187
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1635271187
transform -1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1635271187
transform -1 0 3588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1635271187
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_31
timestamp 1635271187
transform 1 0 3956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_43
timestamp 1635271187
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1635271187
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _328_
timestamp 1635271187
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__RESET_B
timestamp 1635271187
transform -1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_48
timestamp 1635271187
transform 1 0 5520 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1635271187
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1635271187
transform 1 0 5244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _192_
timestamp 1635271187
transform 1 0 6348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _200_
timestamp 1635271187
transform 1 0 7084 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1635271187
transform -1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A1
timestamp 1635271187
transform 1 0 8464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A1
timestamp 1635271187
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_73
timestamp 1635271187
transform 1 0 7820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1635271187
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1635271187
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1635271187
transform -1 0 7820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1635271187
transform -1 0 9752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__S
timestamp 1635271187
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__S
timestamp 1635271187
transform 1 0 9936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1635271187
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_98
timestamp 1635271187
transform 1 0 10120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1635271187
transform 1 0 10212 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1635271187
transform -1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_113
timestamp 1635271187
transform 1 0 11500 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1635271187
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1635271187
transform 1 0 12052 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1635271187
transform 1 0 12696 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_22_133
timestamp 1635271187
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635271187
transform -1 0 13892 0 1 13056
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 8210 13892 8530 6 VGND
port 0 nsew ground input
rlabel metal4 s 8208 1040 8528 13648 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 4210 13892 4530 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 12210 13892 12530 6 VPWR
port 1 nsew power input
rlabel metal4 s 4208 1040 4528 13648 6 VPWR
port 1 nsew power input
rlabel metal4 s 12208 1040 12528 13648 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 3680 800 3800 6 clockp[0]
port 2 nsew signal tristate
rlabel metal3 s 0 11160 800 11280 6 clockp[1]
port 3 nsew signal tristate
rlabel metal3 s 14200 14424 15000 14544 6 dco
port 4 nsew signal input
rlabel metal3 s 14200 10072 15000 10192 6 div[0]
port 5 nsew signal input
rlabel metal3 s 14200 10888 15000 11008 6 div[1]
port 6 nsew signal input
rlabel metal3 s 14200 11840 15000 11960 6 div[2]
port 7 nsew signal input
rlabel metal3 s 14200 12656 15000 12776 6 div[3]
port 8 nsew signal input
rlabel metal3 s 14200 13608 15000 13728 6 div[4]
port 9 nsew signal input
rlabel metal3 s 14200 9120 15000 9240 6 enable
port 10 nsew signal input
rlabel metal2 s 754 14200 810 15000 6 ext_trim[0]
port 11 nsew signal input
rlabel metal3 s 14200 416 15000 536 6 ext_trim[10]
port 12 nsew signal input
rlabel metal3 s 14200 1232 15000 1352 6 ext_trim[11]
port 13 nsew signal input
rlabel metal3 s 14200 2048 15000 2168 6 ext_trim[12]
port 14 nsew signal input
rlabel metal3 s 14200 3000 15000 3120 6 ext_trim[13]
port 15 nsew signal input
rlabel metal3 s 14200 3816 15000 3936 6 ext_trim[14]
port 16 nsew signal input
rlabel metal3 s 14200 4768 15000 4888 6 ext_trim[15]
port 17 nsew signal input
rlabel metal3 s 14200 5584 15000 5704 6 ext_trim[16]
port 18 nsew signal input
rlabel metal3 s 14200 6536 15000 6656 6 ext_trim[17]
port 19 nsew signal input
rlabel metal3 s 14200 7352 15000 7472 6 ext_trim[18]
port 20 nsew signal input
rlabel metal3 s 14200 8304 15000 8424 6 ext_trim[19]
port 21 nsew signal input
rlabel metal2 s 2226 14200 2282 15000 6 ext_trim[1]
port 22 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 ext_trim[20]
port 23 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 ext_trim[21]
port 24 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 ext_trim[22]
port 25 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 ext_trim[23]
port 26 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 ext_trim[24]
port 27 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 ext_trim[25]
port 28 nsew signal input
rlabel metal2 s 3698 14200 3754 15000 6 ext_trim[2]
port 29 nsew signal input
rlabel metal2 s 5170 14200 5226 15000 6 ext_trim[3]
port 30 nsew signal input
rlabel metal2 s 6734 14200 6790 15000 6 ext_trim[4]
port 31 nsew signal input
rlabel metal2 s 8206 14200 8262 15000 6 ext_trim[5]
port 32 nsew signal input
rlabel metal2 s 9678 14200 9734 15000 6 ext_trim[6]
port 33 nsew signal input
rlabel metal2 s 11242 14200 11298 15000 6 ext_trim[7]
port 34 nsew signal input
rlabel metal2 s 12714 14200 12770 15000 6 ext_trim[8]
port 35 nsew signal input
rlabel metal2 s 14186 14200 14242 15000 6 ext_trim[9]
port 36 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 osc
port 37 nsew signal input
rlabel metal2 s 938 0 994 800 6 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
