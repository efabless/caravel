magic
tech sky130A
magscale 1 2
timestamp 1665777668
<< error_s >>
rect 147395 223457 147404 223466
rect 147743 223457 147752 223466
rect 147386 223448 147395 223457
rect 147752 223448 147761 223457
rect 147386 223397 147395 223406
rect 147752 223397 147761 223406
rect 147395 223388 147404 223397
rect 147743 223388 147752 223397
<< locali >>
rect 676932 708260 676938 708478
rect 40621 604574 40627 604792
rect 40621 603378 40627 603596
rect 40621 602182 40627 602400
rect 40621 600986 40627 601204
rect 40621 599790 40627 600008
rect 40621 598594 40627 598812
rect 676932 447436 676938 447654
rect 676932 446240 676938 446458
rect 676932 445044 676938 445262
rect 676932 443848 676938 444066
rect 676932 442652 676938 442870
rect 676932 441456 676938 441674
rect 676932 440260 676938 440478
rect 40643 346393 40649 346611
rect 40643 345197 40649 345415
rect 40643 344001 40649 344219
rect 40643 342805 40649 343023
rect 40643 341609 40649 341827
rect 40643 340413 40649 340631
rect 40643 339217 40649 339435
rect 40643 338021 40649 338239
rect 40643 336825 40649 337043
rect 40643 335629 40649 335847
rect 134848 223204 135066 223210
rect 136044 223204 136262 223210
rect 137240 223204 137458 223210
rect 138436 223204 138654 223210
rect 139632 223204 139850 223210
rect 140828 223204 141046 223210
rect 142024 223204 142242 223210
rect 143220 223204 143438 223210
rect 144416 223204 144634 223210
rect 145612 223204 145830 223210
rect 148004 223204 148222 223210
rect 149200 223204 149418 223210
rect 150396 223204 150614 223210
rect 151592 223204 151810 223210
rect 152788 223204 153006 223210
rect 153984 223204 154202 223210
rect 394848 223204 395066 223210
rect 396044 223204 396262 223210
rect 397240 223204 397458 223210
rect 398436 223204 398654 223210
rect 399632 223204 399850 223210
rect 400828 223204 401046 223210
rect 402024 223204 402242 223210
rect 403220 223204 403438 223210
rect 404416 223204 404634 223210
rect 405612 223204 405830 223210
rect 408004 223204 408222 223210
rect 409200 223204 409418 223210
rect 410396 223204 410614 223210
rect 411592 223204 411810 223210
rect 412788 223204 413006 223210
rect 413984 223204 414202 223210
<< viali >>
rect 676938 708260 676972 708478
rect 677482 708162 677652 708196
rect 676870 707516 677040 707550
rect 677550 707334 677584 707552
rect 40587 604574 40621 604792
rect 39907 604476 40077 604510
rect 39975 603648 40009 603866
rect 40519 603830 40689 603864
rect 40587 603378 40621 603596
rect 39907 603280 40077 603314
rect 39975 602452 40009 602670
rect 40519 602634 40689 602668
rect 40587 602182 40621 602400
rect 39907 602084 40077 602118
rect 39975 601256 40009 601474
rect 40519 601438 40689 601472
rect 40587 600986 40621 601204
rect 39907 600888 40077 600922
rect 39975 600060 40009 600278
rect 40519 600242 40689 600276
rect 40587 599790 40621 600008
rect 39907 599692 40077 599726
rect 39975 598864 40009 599082
rect 40519 599046 40689 599080
rect 40587 598594 40621 598812
rect 39907 598496 40077 598530
rect 39975 597668 40009 597886
rect 40519 597850 40689 597884
rect 676938 447436 676972 447654
rect 677482 447338 677652 447372
rect 676870 446692 677040 446726
rect 677550 446510 677584 446728
rect 676938 446240 676972 446458
rect 677482 446142 677652 446176
rect 676870 445496 677040 445530
rect 677550 445314 677584 445532
rect 676938 445044 676972 445262
rect 677482 444946 677652 444980
rect 676870 444300 677040 444334
rect 677550 444118 677584 444336
rect 676938 443848 676972 444066
rect 677482 443750 677652 443784
rect 676870 443104 677040 443138
rect 677550 442922 677584 443140
rect 676938 442652 676972 442870
rect 677482 442554 677652 442588
rect 676870 441908 677040 441942
rect 677550 441726 677584 441944
rect 676938 441456 676972 441674
rect 677482 441358 677652 441392
rect 676870 440712 677040 440746
rect 677550 440530 677584 440748
rect 676938 440260 676972 440478
rect 677482 440162 677652 440196
rect 676870 439516 677040 439550
rect 677550 439334 677584 439552
rect 40609 346393 40643 346611
rect 39929 346295 40099 346329
rect 39997 345467 40031 345685
rect 40541 345649 40711 345683
rect 40609 345197 40643 345415
rect 39929 345099 40099 345133
rect 39997 344271 40031 344489
rect 40541 344453 40711 344487
rect 40609 344001 40643 344219
rect 39929 343903 40099 343937
rect 39997 343075 40031 343293
rect 40541 343257 40711 343291
rect 40609 342805 40643 343023
rect 39929 342707 40099 342741
rect 39997 341879 40031 342097
rect 40541 342061 40711 342095
rect 40609 341609 40643 341827
rect 39929 341511 40099 341545
rect 39997 340683 40031 340901
rect 40541 340865 40711 340899
rect 40609 340413 40643 340631
rect 39929 340315 40099 340349
rect 39997 339487 40031 339705
rect 40541 339669 40711 339703
rect 40609 339217 40643 339435
rect 39929 339119 40099 339153
rect 39997 338291 40031 338509
rect 40541 338473 40711 338507
rect 40609 338021 40643 338239
rect 39929 337923 40099 337957
rect 39997 337095 40031 337313
rect 40541 337277 40711 337311
rect 40609 336825 40643 337043
rect 39929 336727 40099 336761
rect 39997 335899 40031 336117
rect 40541 336081 40711 336115
rect 40609 335629 40643 335847
rect 39929 335531 40099 335565
rect 39997 334703 40031 334921
rect 40541 334885 40711 334919
rect 134104 223102 134138 223272
rect 134848 223170 135066 223204
rect 135300 223102 135334 223272
rect 136044 223170 136262 223204
rect 136496 223102 136530 223272
rect 137240 223170 137458 223204
rect 137692 223102 137726 223272
rect 138436 223170 138654 223204
rect 138888 223102 138922 223272
rect 139632 223170 139850 223204
rect 140084 223102 140118 223272
rect 140828 223170 141046 223204
rect 141280 223102 141314 223272
rect 142024 223170 142242 223204
rect 142476 223102 142510 223272
rect 143220 223170 143438 223204
rect 143672 223102 143706 223272
rect 144416 223170 144634 223204
rect 144868 223102 144902 223272
rect 145612 223170 145830 223204
rect 147260 223102 147294 223272
rect 148004 223170 148222 223204
rect 148456 223102 148490 223272
rect 149200 223170 149418 223204
rect 149652 223102 149686 223272
rect 150396 223170 150614 223204
rect 150848 223102 150882 223272
rect 151592 223170 151810 223204
rect 152044 223102 152078 223272
rect 152788 223170 153006 223204
rect 153240 223102 153274 223272
rect 153984 223170 154202 223204
rect 394104 223102 394138 223272
rect 394848 223170 395066 223204
rect 395300 223102 395334 223272
rect 396044 223170 396262 223204
rect 396496 223102 396530 223272
rect 397240 223170 397458 223204
rect 397692 223102 397726 223272
rect 398436 223170 398654 223204
rect 398888 223102 398922 223272
rect 399632 223170 399850 223204
rect 400084 223102 400118 223272
rect 400828 223170 401046 223204
rect 401280 223102 401314 223272
rect 402024 223170 402242 223204
rect 402476 223102 402510 223272
rect 403220 223170 403438 223204
rect 403672 223102 403706 223272
rect 404416 223170 404634 223204
rect 404868 223102 404902 223272
rect 405612 223170 405830 223204
rect 407260 223102 407294 223272
rect 408004 223170 408222 223204
rect 408456 223102 408490 223272
rect 409200 223170 409418 223204
rect 409652 223102 409686 223272
rect 410396 223170 410614 223204
rect 410848 223102 410882 223272
rect 411592 223170 411810 223204
rect 412044 223102 412078 223272
rect 412788 223170 413006 223204
rect 413240 223102 413274 223272
rect 413984 223170 414202 223204
rect 135118 222558 135336 222592
rect 135946 222490 135980 222660
rect 136314 222558 136532 222592
rect 137142 222490 137176 222660
rect 137510 222558 137728 222592
rect 138338 222490 138372 222660
rect 138706 222558 138924 222592
rect 139534 222490 139568 222660
rect 139902 222558 140120 222592
rect 140730 222490 140764 222660
rect 141098 222558 141316 222592
rect 141926 222490 141960 222660
rect 142294 222558 142512 222592
rect 143122 222490 143156 222660
rect 143490 222558 143708 222592
rect 144318 222490 144352 222660
rect 144686 222558 144904 222592
rect 145514 222490 145548 222660
rect 145882 222558 146100 222592
rect 146710 222490 146744 222660
rect 148274 222558 148492 222592
rect 149102 222490 149136 222660
rect 149470 222558 149688 222592
rect 150298 222490 150332 222660
rect 150666 222558 150884 222592
rect 151494 222490 151528 222660
rect 151862 222558 152080 222592
rect 152690 222490 152724 222660
rect 153240 222490 153274 222660
rect 153884 222558 154102 222592
rect 395118 222558 395336 222592
rect 395946 222490 395980 222660
rect 396314 222558 396532 222592
rect 397142 222490 397176 222660
rect 397510 222558 397728 222592
rect 398338 222490 398372 222660
rect 398706 222558 398924 222592
rect 399534 222490 399568 222660
rect 399902 222558 400120 222592
rect 400730 222490 400764 222660
rect 401098 222558 401316 222592
rect 401926 222490 401960 222660
rect 402294 222558 402512 222592
rect 403122 222490 403156 222660
rect 403490 222558 403708 222592
rect 404318 222490 404352 222660
rect 404686 222558 404904 222592
rect 405514 222490 405548 222660
rect 405882 222558 406100 222592
rect 406710 222490 406744 222660
rect 408274 222558 408492 222592
rect 409102 222490 409136 222660
rect 409470 222558 409688 222592
rect 410298 222490 410332 222660
rect 410666 222558 410884 222592
rect 411494 222490 411528 222660
rect 411862 222558 412080 222592
rect 412690 222490 412724 222660
rect 413240 222490 413274 222660
rect 413884 222558 414102 222592
<< metal1 >>
rect 676296 708223 676324 714921
rect 676352 708417 676380 715121
rect 676928 708478 676980 708490
rect 676352 708411 676404 708417
rect 676352 708353 676404 708359
rect 676928 708248 676980 708260
rect 676296 708217 676348 708223
rect 676296 708159 676348 708165
rect 677470 708152 677482 708204
rect 677652 708152 677664 708204
rect 676356 707568 676408 707574
rect 676356 707510 676408 707516
rect 676324 707450 676352 707455
rect 676300 707444 676352 707450
rect 676300 707386 676352 707392
rect 40579 604792 40631 604804
rect 41203 604731 41231 613556
rect 41179 604725 41231 604731
rect 41179 604667 41231 604673
rect 40579 604562 40631 604574
rect 41259 604537 41287 613356
rect 41235 604531 41287 604537
rect 39895 604466 39907 604518
rect 40077 604466 40089 604518
rect 41235 604473 41287 604479
rect 41175 603882 41227 603888
rect 39967 603866 40019 603878
rect 40507 603820 40519 603872
rect 40689 603820 40701 603872
rect 41175 603824 41227 603830
rect 39967 603636 40019 603648
rect 40579 603596 40631 603608
rect 40579 603366 40631 603378
rect 39895 603270 39907 603322
rect 40077 603270 40089 603322
rect 39967 602670 40019 602682
rect 40507 602624 40519 602676
rect 40689 602624 40701 602676
rect 39967 602440 40019 602452
rect 40579 602400 40631 602412
rect 40579 602170 40631 602182
rect 39895 602074 39907 602126
rect 40077 602074 40089 602126
rect 39967 601474 40019 601486
rect 40507 601428 40519 601480
rect 40689 601428 40701 601480
rect 39967 601244 40019 601256
rect 40579 601204 40631 601216
rect 40579 600974 40631 600986
rect 39895 600878 39907 600930
rect 40077 600878 40089 600930
rect 39967 600278 40019 600290
rect 40507 600232 40519 600284
rect 40689 600232 40701 600284
rect 39967 600048 40019 600060
rect 40579 600008 40631 600020
rect 40579 599778 40631 599790
rect 39895 599682 39907 599734
rect 40077 599682 40089 599734
rect 39967 599082 40019 599094
rect 40507 599036 40519 599088
rect 40689 599036 40701 599088
rect 39967 598852 40019 598864
rect 40579 598812 40631 598824
rect 40579 598582 40631 598594
rect 39895 598486 39907 598538
rect 40077 598486 40089 598538
rect 39967 597886 40019 597898
rect 40507 597840 40519 597892
rect 40689 597840 40701 597892
rect 39967 597656 40019 597668
rect 40601 346611 40653 346623
rect 41175 346550 41203 603824
rect 41151 346544 41203 346550
rect 41151 346486 41203 346492
rect 41231 603758 41283 603764
rect 41231 603700 41283 603706
rect 40601 346381 40653 346393
rect 41231 346356 41259 603700
rect 41315 603535 41343 613156
rect 41291 603529 41343 603535
rect 41291 603471 41343 603477
rect 41371 603341 41399 612956
rect 41347 603335 41399 603341
rect 41347 603277 41399 603283
rect 41207 346350 41259 346356
rect 39917 346285 39929 346337
rect 40099 346285 40111 346337
rect 41207 346292 41259 346298
rect 41287 602686 41339 602692
rect 41287 602628 41339 602634
rect 41147 345701 41199 345707
rect 39989 345685 40041 345697
rect 40529 345639 40541 345691
rect 40711 345639 40723 345691
rect 41147 345643 41199 345649
rect 39989 345455 40041 345467
rect 40601 345415 40653 345427
rect 40601 345185 40653 345197
rect 39917 345089 39929 345141
rect 40099 345089 40111 345141
rect 39989 344489 40041 344501
rect 40529 344443 40541 344495
rect 40711 344443 40723 344495
rect 39989 344259 40041 344271
rect 40601 344219 40653 344231
rect 40601 343989 40653 344001
rect 39917 343893 39929 343945
rect 40099 343893 40111 343945
rect 39989 343293 40041 343305
rect 40529 343247 40541 343299
rect 40711 343247 40723 343299
rect 39989 343063 40041 343075
rect 40601 343023 40653 343035
rect 40601 342793 40653 342805
rect 39917 342697 39929 342749
rect 40099 342697 40111 342749
rect 39989 342097 40041 342109
rect 40529 342051 40541 342103
rect 40711 342051 40723 342103
rect 39989 341867 40041 341879
rect 40601 341827 40653 341839
rect 40601 341597 40653 341609
rect 39917 341501 39929 341553
rect 40099 341501 40111 341553
rect 39989 340901 40041 340913
rect 40529 340855 40541 340907
rect 40711 340855 40723 340907
rect 39989 340671 40041 340683
rect 40601 340631 40653 340643
rect 40601 340401 40653 340413
rect 39917 340305 39929 340357
rect 40099 340305 40111 340357
rect 39989 339705 40041 339717
rect 40529 339659 40541 339711
rect 40711 339659 40723 339711
rect 39989 339475 40041 339487
rect 40601 339435 40653 339447
rect 40601 339205 40653 339217
rect 39917 339109 39929 339161
rect 40099 339109 40111 339161
rect 39989 338509 40041 338521
rect 40529 338463 40541 338515
rect 40711 338463 40723 338515
rect 39989 338279 40041 338291
rect 40601 338239 40653 338251
rect 40601 338009 40653 338021
rect 39917 337913 39929 337965
rect 40099 337913 40111 337965
rect 39989 337313 40041 337325
rect 40529 337267 40541 337319
rect 40711 337267 40723 337319
rect 39989 337083 40041 337095
rect 40601 337043 40653 337055
rect 40601 336813 40653 336825
rect 39917 336717 39929 336769
rect 40099 336717 40111 336769
rect 39989 336117 40041 336129
rect 40529 336071 40541 336123
rect 40711 336071 40723 336123
rect 39989 335887 40041 335899
rect 40601 335847 40653 335859
rect 40601 335617 40653 335629
rect 39917 335521 39929 335573
rect 40099 335521 40111 335573
rect 39989 334921 40041 334933
rect 40529 334875 40541 334927
rect 40711 334875 40723 334927
rect 39989 334691 40041 334703
rect 41147 224252 41175 345643
rect 41203 345577 41255 345583
rect 41203 345519 41255 345525
rect 41203 224308 41231 345519
rect 41287 345354 41315 602628
rect 41263 345348 41315 345354
rect 41263 345290 41315 345296
rect 41343 602562 41395 602568
rect 41343 602504 41395 602510
rect 41343 345160 41371 602504
rect 41427 602339 41455 612756
rect 41403 602333 41455 602339
rect 41403 602275 41455 602281
rect 41483 602145 41511 612556
rect 41459 602139 41511 602145
rect 41459 602081 41511 602087
rect 41319 345154 41371 345160
rect 41319 345096 41371 345102
rect 41399 601490 41451 601496
rect 41399 601432 41451 601438
rect 41259 344505 41311 344511
rect 41259 344447 41311 344453
rect 41259 224364 41287 344447
rect 41315 344381 41367 344387
rect 41315 344323 41367 344329
rect 41315 224420 41343 344323
rect 41399 344158 41427 601432
rect 41375 344152 41427 344158
rect 41375 344094 41427 344100
rect 41455 601366 41507 601372
rect 41455 601308 41507 601314
rect 41455 343964 41483 601308
rect 41539 601143 41567 612356
rect 41515 601137 41567 601143
rect 41515 601079 41567 601085
rect 41595 600949 41623 612156
rect 41571 600943 41623 600949
rect 41571 600885 41623 600891
rect 41431 343958 41483 343964
rect 41431 343900 41483 343906
rect 41511 600294 41563 600300
rect 41511 600236 41563 600242
rect 41371 343309 41423 343315
rect 41371 343251 41423 343257
rect 41371 224476 41399 343251
rect 41427 343185 41479 343191
rect 41427 343127 41479 343133
rect 41427 224532 41455 343127
rect 41511 342962 41539 600236
rect 41487 342956 41539 342962
rect 41487 342898 41539 342904
rect 41567 600170 41619 600176
rect 41567 600112 41619 600118
rect 41567 342768 41595 600112
rect 41651 599947 41679 611956
rect 41627 599941 41679 599947
rect 41627 599883 41679 599889
rect 41707 599753 41735 611756
rect 41683 599747 41735 599753
rect 41683 599689 41735 599695
rect 41543 342762 41595 342768
rect 41543 342704 41595 342710
rect 41623 599098 41675 599104
rect 41623 599040 41675 599046
rect 41483 342113 41535 342119
rect 41483 342055 41535 342061
rect 41483 224588 41511 342055
rect 41539 341989 41591 341995
rect 41539 341931 41591 341937
rect 41539 224644 41567 341931
rect 41623 341766 41651 599040
rect 41599 341760 41651 341766
rect 41599 341702 41651 341708
rect 41679 598974 41731 598980
rect 41679 598916 41731 598922
rect 41679 341572 41707 598916
rect 41763 598751 41791 611556
rect 41739 598745 41791 598751
rect 41739 598687 41791 598693
rect 41819 598557 41847 611356
rect 41795 598551 41847 598557
rect 41795 598493 41847 598499
rect 41655 341566 41707 341572
rect 41655 341508 41707 341514
rect 41735 597902 41787 597908
rect 41735 597844 41787 597850
rect 41595 340917 41647 340923
rect 41595 340859 41647 340865
rect 41595 224700 41623 340859
rect 41651 340793 41703 340799
rect 41651 340735 41703 340741
rect 41651 224756 41679 340735
rect 41735 340570 41763 597844
rect 41711 340564 41763 340570
rect 41711 340506 41763 340512
rect 41791 597778 41843 597784
rect 41791 597720 41843 597726
rect 41791 340376 41819 597720
rect 675624 440223 675652 454055
rect 675680 440417 675708 454255
rect 675736 441419 675764 454455
rect 675792 441613 675820 454655
rect 675848 442615 675876 454855
rect 675904 442809 675932 455055
rect 675960 443811 675988 455255
rect 676016 444005 676044 455455
rect 676072 445007 676100 455655
rect 676128 445201 676156 455855
rect 676184 446203 676212 456055
rect 676240 446397 676268 456255
rect 676324 455108 676352 707386
rect 676296 455079 676352 455108
rect 676296 447399 676324 455079
rect 676380 455050 676408 707510
rect 676858 707506 676870 707558
rect 677040 707506 677052 707558
rect 677540 707552 677592 707564
rect 677540 707322 677592 707334
rect 677213 706869 677309 707220
rect 677213 706512 677234 706869
rect 677294 706512 677309 706869
rect 677213 706498 677309 706512
rect 676352 455020 676408 455050
rect 676352 447593 676380 455020
rect 676928 447654 676980 447666
rect 676352 447587 676404 447593
rect 676352 447529 676404 447535
rect 676928 447424 676980 447436
rect 676296 447393 676348 447399
rect 676296 447335 676348 447341
rect 677470 447328 677482 447380
rect 677652 447328 677664 447380
rect 676356 446744 676408 446750
rect 676356 446686 676408 446692
rect 676300 446620 676352 446626
rect 676300 446562 676352 446568
rect 676240 446391 676292 446397
rect 676240 446333 676292 446339
rect 676184 446197 676236 446203
rect 676184 446139 676236 446145
rect 676244 445548 676296 445554
rect 676244 445490 676296 445496
rect 676188 445424 676240 445430
rect 676188 445366 676240 445372
rect 676128 445195 676180 445201
rect 676128 445137 676180 445143
rect 676072 445001 676124 445007
rect 676072 444943 676124 444949
rect 676132 444352 676184 444358
rect 676132 444294 676184 444300
rect 676076 444228 676128 444234
rect 676076 444170 676128 444176
rect 676016 443999 676068 444005
rect 676016 443941 676068 443947
rect 675960 443805 676012 443811
rect 675960 443747 676012 443753
rect 676020 443156 676072 443162
rect 676020 443098 676072 443104
rect 675964 443032 676016 443038
rect 675964 442974 676016 442980
rect 675904 442803 675956 442809
rect 675904 442745 675956 442751
rect 675848 442609 675900 442615
rect 675848 442551 675900 442557
rect 675908 441960 675960 441966
rect 675908 441902 675960 441908
rect 675852 441836 675904 441842
rect 675852 441778 675904 441784
rect 675792 441607 675844 441613
rect 675792 441549 675844 441555
rect 675736 441413 675788 441419
rect 675736 441355 675788 441361
rect 675796 440764 675848 440770
rect 675796 440706 675848 440712
rect 675740 440640 675792 440646
rect 675740 440582 675792 440588
rect 675680 440411 675732 440417
rect 675680 440353 675732 440359
rect 675624 440217 675676 440223
rect 675624 440159 675676 440165
rect 675684 439568 675736 439574
rect 675684 439510 675736 439516
rect 675628 439444 675680 439450
rect 675628 439386 675680 439392
rect 41767 340370 41819 340376
rect 41767 340312 41819 340318
rect 41707 339721 41759 339727
rect 41707 339663 41759 339669
rect 41707 224812 41735 339663
rect 41763 339597 41815 339603
rect 41763 339539 41815 339545
rect 41763 224868 41791 339539
rect 41847 339374 41875 354730
rect 41823 339368 41875 339374
rect 41823 339310 41875 339316
rect 41903 339180 41931 354530
rect 41879 339174 41931 339180
rect 41879 339116 41931 339122
rect 41819 338525 41871 338531
rect 41819 338467 41871 338473
rect 41819 224924 41847 338467
rect 41875 338401 41927 338407
rect 41875 338343 41927 338349
rect 41875 224980 41903 338343
rect 41959 338178 41987 354330
rect 41935 338172 41987 338178
rect 41935 338114 41987 338120
rect 42015 337984 42043 354130
rect 41991 337978 42043 337984
rect 41991 337920 42043 337926
rect 41931 337329 41983 337335
rect 41931 337271 41983 337277
rect 41931 225036 41959 337271
rect 41987 337205 42039 337211
rect 41987 337147 42039 337153
rect 41987 225092 42015 337147
rect 42071 336958 42099 353930
rect 42047 336952 42099 336958
rect 42047 336894 42099 336900
rect 42127 336788 42155 353730
rect 42103 336782 42155 336788
rect 42103 336724 42155 336730
rect 42043 336133 42095 336139
rect 42043 336075 42095 336081
rect 42043 225148 42071 336075
rect 42099 336009 42151 336015
rect 42099 335951 42151 335957
rect 42099 225204 42127 335951
rect 42183 335786 42211 353530
rect 42159 335780 42211 335786
rect 42159 335722 42211 335728
rect 42239 335592 42267 353330
rect 42215 335586 42267 335592
rect 42215 335528 42267 335534
rect 42155 334937 42207 334943
rect 42155 334879 42207 334885
rect 42155 225260 42183 334879
rect 42211 334813 42263 334819
rect 42211 334755 42263 334761
rect 42211 225316 42239 334755
rect 394098 225344 394104 225368
rect 134098 225316 134104 225340
rect 42211 225288 134104 225316
rect 134156 225288 134162 225340
rect 134941 225292 134947 225344
rect 134999 225316 394104 225344
rect 394156 225316 394162 225368
rect 394941 225320 394947 225372
rect 394999 225344 675568 225372
rect 394999 225320 395005 225344
rect 134999 225292 135005 225316
rect 395170 225288 395176 225312
rect 135170 225260 135176 225284
rect 42155 225232 135176 225260
rect 135228 225232 135234 225284
rect 135943 225236 135949 225288
rect 136001 225260 395176 225288
rect 395228 225260 395234 225312
rect 395943 225264 395949 225316
rect 396001 225288 675512 225316
rect 396001 225264 396007 225288
rect 136001 225236 136007 225260
rect 395294 225232 395300 225256
rect 135294 225204 135300 225228
rect 42099 225176 135300 225204
rect 135352 225176 135358 225228
rect 136137 225180 136143 225232
rect 136195 225204 395300 225232
rect 395352 225204 395358 225256
rect 396137 225208 396143 225260
rect 396195 225232 675456 225260
rect 396195 225208 396201 225232
rect 136195 225180 136201 225204
rect 396366 225176 396372 225200
rect 136366 225148 136372 225172
rect 42043 225120 136372 225148
rect 136424 225120 136430 225172
rect 137139 225124 137145 225176
rect 137197 225148 396372 225176
rect 396424 225148 396430 225200
rect 397139 225152 397145 225204
rect 397197 225176 675400 225204
rect 397197 225152 397203 225176
rect 137197 225124 137203 225148
rect 396490 225120 396496 225144
rect 136490 225092 136496 225116
rect 41987 225064 136496 225092
rect 136548 225064 136554 225116
rect 137333 225068 137339 225120
rect 137391 225092 396496 225120
rect 396548 225092 396554 225144
rect 397333 225096 397339 225148
rect 397391 225120 675344 225148
rect 397391 225096 397397 225120
rect 137391 225068 137397 225092
rect 397562 225064 397568 225088
rect 137562 225036 137568 225060
rect 41931 225008 137568 225036
rect 137620 225008 137626 225060
rect 138335 225012 138341 225064
rect 138393 225036 397568 225064
rect 397620 225036 397626 225088
rect 398335 225040 398341 225092
rect 398393 225064 675288 225092
rect 398393 225040 398399 225064
rect 138393 225012 138399 225036
rect 397686 225008 397692 225032
rect 137686 224980 137692 225004
rect 41875 224952 137692 224980
rect 137744 224952 137750 225004
rect 138529 224956 138535 225008
rect 138587 224980 397692 225008
rect 397744 224980 397750 225032
rect 398529 224984 398535 225036
rect 398587 225008 675232 225036
rect 398587 224984 398593 225008
rect 138587 224956 138593 224980
rect 398758 224952 398764 224976
rect 138758 224924 138764 224948
rect 41819 224896 138764 224924
rect 138816 224896 138822 224948
rect 139531 224900 139537 224952
rect 139589 224924 398764 224952
rect 398816 224924 398822 224976
rect 399531 224928 399537 224980
rect 399589 224952 675176 224980
rect 399589 224928 399595 224952
rect 139589 224900 139595 224924
rect 398882 224896 398888 224920
rect 138882 224868 138888 224892
rect 41763 224840 138888 224868
rect 138940 224840 138946 224892
rect 139725 224844 139731 224896
rect 139783 224868 398888 224896
rect 398940 224868 398946 224920
rect 399725 224872 399731 224924
rect 399783 224896 675120 224924
rect 399783 224872 399789 224896
rect 139783 224844 139789 224868
rect 399954 224840 399960 224864
rect 139954 224812 139960 224836
rect 41707 224784 139960 224812
rect 140012 224784 140018 224836
rect 140727 224788 140733 224840
rect 140785 224812 399960 224840
rect 400012 224812 400018 224864
rect 400727 224816 400733 224868
rect 400785 224840 675064 224868
rect 400785 224816 400791 224840
rect 140785 224788 140791 224812
rect 400078 224784 400084 224808
rect 140078 224756 140084 224780
rect 41651 224728 140084 224756
rect 140136 224728 140142 224780
rect 140897 224732 140903 224784
rect 140955 224756 400084 224784
rect 400136 224756 400142 224808
rect 400897 224760 400903 224812
rect 400955 224784 675008 224812
rect 400955 224760 400961 224784
rect 140955 224732 140961 224756
rect 401150 224728 401156 224752
rect 141150 224700 141156 224724
rect 41595 224672 141156 224700
rect 141208 224672 141214 224724
rect 141923 224676 141929 224728
rect 141981 224700 401156 224728
rect 401208 224700 401214 224752
rect 401923 224704 401929 224756
rect 401981 224728 674952 224756
rect 401981 224704 401987 224728
rect 141981 224676 141987 224700
rect 401274 224672 401280 224696
rect 141274 224644 141280 224668
rect 41539 224616 141280 224644
rect 141332 224616 141338 224668
rect 142117 224620 142123 224672
rect 142175 224644 401280 224672
rect 401332 224644 401338 224696
rect 402117 224648 402123 224700
rect 402175 224672 674896 224700
rect 402175 224648 402181 224672
rect 142175 224620 142181 224644
rect 402346 224616 402352 224640
rect 142346 224588 142352 224612
rect 41483 224560 142352 224588
rect 142404 224560 142410 224612
rect 143119 224564 143125 224616
rect 143177 224588 402352 224616
rect 402404 224588 402410 224640
rect 403119 224592 403125 224644
rect 403177 224616 674840 224644
rect 403177 224592 403183 224616
rect 143177 224564 143183 224588
rect 402470 224560 402476 224584
rect 142470 224532 142476 224556
rect 41427 224504 142476 224532
rect 142528 224504 142534 224556
rect 143289 224508 143295 224560
rect 143347 224532 402476 224560
rect 402528 224532 402534 224584
rect 403289 224536 403295 224588
rect 403347 224560 674784 224588
rect 403347 224536 403353 224560
rect 143347 224508 143353 224532
rect 403542 224504 403548 224528
rect 143542 224476 143548 224500
rect 41371 224448 143548 224476
rect 143600 224448 143606 224500
rect 144315 224452 144321 224504
rect 144373 224476 403548 224504
rect 403600 224476 403606 224528
rect 404315 224480 404321 224532
rect 404373 224504 674728 224532
rect 404373 224480 404379 224504
rect 144373 224452 144379 224476
rect 403666 224448 403672 224472
rect 143666 224420 143672 224444
rect 41315 224392 143672 224420
rect 143724 224392 143730 224444
rect 144509 224396 144515 224448
rect 144567 224420 403672 224448
rect 403724 224420 403730 224472
rect 404509 224424 404515 224476
rect 404567 224448 674672 224476
rect 404567 224424 404573 224448
rect 144567 224396 144573 224420
rect 404738 224392 404744 224416
rect 144738 224364 144744 224388
rect 41259 224336 144744 224364
rect 144796 224336 144802 224388
rect 145511 224340 145517 224392
rect 145569 224364 404744 224392
rect 404796 224364 404802 224416
rect 405511 224368 405517 224420
rect 405569 224392 674616 224420
rect 405569 224368 405575 224392
rect 145569 224340 145575 224364
rect 404862 224336 404868 224360
rect 144862 224308 144868 224332
rect 41203 224280 144868 224308
rect 144920 224280 144926 224332
rect 145705 224284 145711 224336
rect 145763 224308 404868 224336
rect 404920 224308 404926 224360
rect 405705 224312 405711 224364
rect 405763 224336 674560 224364
rect 405763 224312 405769 224336
rect 145763 224284 145769 224308
rect 405934 224280 405940 224304
rect 145934 224252 145940 224276
rect 41147 224224 145940 224252
rect 145992 224224 145998 224276
rect 146600 224252 146713 224280
rect 146707 224228 146713 224252
rect 146765 224252 405940 224280
rect 405992 224252 405998 224304
rect 406707 224256 406713 224308
rect 406765 224280 674504 224308
rect 406765 224256 406771 224280
rect 146765 224228 146771 224252
rect 407254 224224 407260 224248
rect 147254 224196 147260 224220
rect 131123 224168 147260 224196
rect 147312 224168 147318 224220
rect 148097 224172 148103 224224
rect 148155 224196 407260 224224
rect 407312 224196 407318 224248
rect 408097 224200 408103 224252
rect 408155 224224 674448 224252
rect 408155 224200 408161 224224
rect 148155 224172 148161 224196
rect 408326 224168 408332 224192
rect 148326 224140 148332 224164
rect 131323 224112 148332 224140
rect 148384 224112 148390 224164
rect 149099 224116 149105 224168
rect 149157 224140 408332 224168
rect 408384 224140 408390 224192
rect 409099 224144 409105 224196
rect 409157 224168 674392 224196
rect 409157 224144 409163 224168
rect 149157 224116 149163 224140
rect 408450 224112 408456 224136
rect 148450 224084 148456 224108
rect 131523 224056 148456 224084
rect 148508 224056 148514 224108
rect 149293 224060 149299 224112
rect 149351 224084 408456 224112
rect 408508 224084 408514 224136
rect 409293 224088 409299 224140
rect 409351 224112 674336 224140
rect 409351 224088 409357 224112
rect 149351 224060 149357 224084
rect 409522 224056 409528 224080
rect 149522 224028 149528 224052
rect 131723 224000 149528 224028
rect 149580 224000 149586 224052
rect 150295 224004 150301 224056
rect 150353 224028 409528 224056
rect 409580 224028 409586 224080
rect 410295 224032 410301 224084
rect 410353 224056 674280 224084
rect 410353 224032 410359 224056
rect 150353 224004 150359 224028
rect 409646 224000 409652 224024
rect 149646 223972 149652 223996
rect 131923 223944 149652 223972
rect 149704 223944 149710 223996
rect 150465 223948 150471 224000
rect 150523 223972 409652 224000
rect 409704 223972 409710 224024
rect 410465 223976 410471 224028
rect 410523 224000 674224 224028
rect 410523 223976 410529 224000
rect 150523 223948 150529 223972
rect 410718 223944 410724 223968
rect 150718 223916 150724 223940
rect 132123 223888 150724 223916
rect 150776 223888 150782 223940
rect 151491 223892 151497 223944
rect 151549 223916 410724 223944
rect 410776 223916 410782 223968
rect 411491 223920 411497 223972
rect 411549 223944 674168 223972
rect 411549 223920 411555 223944
rect 151549 223892 151555 223916
rect 410842 223888 410848 223912
rect 150842 223860 150848 223884
rect 132323 223832 150848 223860
rect 150900 223832 150906 223884
rect 151685 223836 151691 223888
rect 151743 223860 410848 223888
rect 410900 223860 410906 223912
rect 411685 223864 411691 223916
rect 411743 223888 674112 223916
rect 411743 223864 411749 223888
rect 151743 223836 151749 223860
rect 411914 223832 411920 223856
rect 151914 223804 151920 223828
rect 132523 223776 151920 223804
rect 151972 223776 151978 223828
rect 152687 223780 152693 223832
rect 152745 223804 411920 223832
rect 411972 223804 411978 223856
rect 412687 223808 412693 223860
rect 412745 223832 674056 223860
rect 412745 223808 412751 223832
rect 152745 223780 152751 223804
rect 412038 223776 412044 223800
rect 152038 223748 152044 223772
rect 132723 223720 152044 223748
rect 152096 223720 152102 223772
rect 152857 223724 152863 223776
rect 152915 223748 412044 223776
rect 412096 223748 412102 223800
rect 412857 223752 412863 223804
rect 412915 223776 674000 223804
rect 412915 223752 412921 223776
rect 152915 223724 152921 223748
rect 413110 223720 413116 223744
rect 153110 223692 153116 223716
rect 132923 223664 153116 223692
rect 153168 223664 153174 223716
rect 153883 223668 153889 223720
rect 153941 223692 413116 223720
rect 413168 223692 413174 223744
rect 413883 223696 413889 223748
rect 413941 223720 673944 223748
rect 413941 223696 413947 223720
rect 153941 223668 153947 223692
rect 413234 223664 413240 223688
rect 153234 223636 153240 223660
rect 133123 223608 153240 223636
rect 153292 223608 153298 223660
rect 154077 223612 154083 223664
rect 154135 223636 413240 223664
rect 413292 223636 413298 223688
rect 414077 223640 414083 223692
rect 414135 223664 673888 223692
rect 414135 223640 414141 223664
rect 154135 223612 154141 223636
rect 134094 223272 134146 223284
rect 135290 223272 135342 223284
rect 134836 223162 134848 223214
rect 135066 223162 135078 223214
rect 134094 223090 134146 223102
rect 136486 223272 136538 223284
rect 136032 223162 136044 223214
rect 136262 223162 136274 223214
rect 135290 223090 135342 223102
rect 137682 223272 137734 223284
rect 137228 223162 137240 223214
rect 137458 223162 137470 223214
rect 136486 223090 136538 223102
rect 138878 223272 138930 223284
rect 138424 223162 138436 223214
rect 138654 223162 138666 223214
rect 137682 223090 137734 223102
rect 140074 223272 140126 223284
rect 139620 223162 139632 223214
rect 139850 223162 139862 223214
rect 138878 223090 138930 223102
rect 141270 223272 141322 223284
rect 140816 223162 140828 223214
rect 141046 223162 141058 223214
rect 140074 223090 140126 223102
rect 142466 223272 142518 223284
rect 142012 223162 142024 223214
rect 142242 223162 142254 223214
rect 141270 223090 141322 223102
rect 143662 223272 143714 223284
rect 143208 223162 143220 223214
rect 143438 223162 143450 223214
rect 142466 223090 142518 223102
rect 144858 223272 144910 223284
rect 144404 223162 144416 223214
rect 144634 223162 144646 223214
rect 143662 223090 143714 223102
rect 147250 223272 147302 223284
rect 145600 223162 145612 223214
rect 145830 223162 145842 223214
rect 144858 223090 144910 223102
rect 148446 223272 148498 223284
rect 147992 223162 148004 223214
rect 148222 223162 148234 223214
rect 147250 223090 147302 223102
rect 149642 223272 149694 223284
rect 149188 223162 149200 223214
rect 149418 223162 149430 223214
rect 148446 223090 148498 223102
rect 150838 223272 150890 223284
rect 150384 223162 150396 223214
rect 150614 223162 150626 223214
rect 149642 223090 149694 223102
rect 152034 223272 152086 223284
rect 151580 223162 151592 223214
rect 151810 223162 151822 223214
rect 150838 223090 150890 223102
rect 153230 223272 153282 223284
rect 152776 223162 152788 223214
rect 153006 223162 153018 223214
rect 152034 223090 152086 223102
rect 394094 223272 394146 223284
rect 153972 223162 153984 223214
rect 154202 223162 154214 223214
rect 153230 223090 153282 223102
rect 395290 223272 395342 223284
rect 394836 223162 394848 223214
rect 395066 223162 395078 223214
rect 394094 223090 394146 223102
rect 396486 223272 396538 223284
rect 396032 223162 396044 223214
rect 396262 223162 396274 223214
rect 395290 223090 395342 223102
rect 397682 223272 397734 223284
rect 397228 223162 397240 223214
rect 397458 223162 397470 223214
rect 396486 223090 396538 223102
rect 398878 223272 398930 223284
rect 398424 223162 398436 223214
rect 398654 223162 398666 223214
rect 397682 223090 397734 223102
rect 400074 223272 400126 223284
rect 399620 223162 399632 223214
rect 399850 223162 399862 223214
rect 398878 223090 398930 223102
rect 401270 223272 401322 223284
rect 400816 223162 400828 223214
rect 401046 223162 401058 223214
rect 400074 223090 400126 223102
rect 402466 223272 402518 223284
rect 402012 223162 402024 223214
rect 402242 223162 402254 223214
rect 401270 223090 401322 223102
rect 403662 223272 403714 223284
rect 403208 223162 403220 223214
rect 403438 223162 403450 223214
rect 402466 223090 402518 223102
rect 404858 223272 404910 223284
rect 404404 223162 404416 223214
rect 404634 223162 404646 223214
rect 403662 223090 403714 223102
rect 407250 223272 407302 223284
rect 405600 223162 405612 223214
rect 405830 223162 405842 223214
rect 404858 223090 404910 223102
rect 408446 223272 408498 223284
rect 407992 223162 408004 223214
rect 408222 223162 408234 223214
rect 407250 223090 407302 223102
rect 409642 223272 409694 223284
rect 409188 223162 409200 223214
rect 409418 223162 409430 223214
rect 408446 223090 408498 223102
rect 410838 223272 410890 223284
rect 410384 223162 410396 223214
rect 410614 223162 410626 223214
rect 409642 223090 409694 223102
rect 412034 223272 412086 223284
rect 411580 223162 411592 223214
rect 411810 223162 411822 223214
rect 410838 223090 410890 223102
rect 413230 223272 413282 223284
rect 412776 223162 412788 223214
rect 413006 223162 413018 223214
rect 412034 223090 412086 223102
rect 413972 223162 413984 223214
rect 414202 223162 414214 223214
rect 413230 223090 413282 223102
rect 135936 222660 135988 222672
rect 135106 222550 135118 222602
rect 135336 222550 135348 222602
rect 137132 222660 137184 222672
rect 136302 222550 136314 222602
rect 136532 222550 136544 222602
rect 135936 222478 135988 222490
rect 138328 222660 138380 222672
rect 137498 222550 137510 222602
rect 137728 222550 137740 222602
rect 137132 222478 137184 222490
rect 139524 222660 139576 222672
rect 138694 222550 138706 222602
rect 138924 222550 138936 222602
rect 138328 222478 138380 222490
rect 140720 222660 140772 222672
rect 139890 222550 139902 222602
rect 140120 222550 140132 222602
rect 139524 222478 139576 222490
rect 141916 222660 141968 222672
rect 141086 222550 141098 222602
rect 141316 222550 141328 222602
rect 140720 222478 140772 222490
rect 143112 222660 143164 222672
rect 142282 222550 142294 222602
rect 142512 222550 142524 222602
rect 141916 222478 141968 222490
rect 144308 222660 144360 222672
rect 143478 222550 143490 222602
rect 143708 222550 143720 222602
rect 143112 222478 143164 222490
rect 145504 222660 145556 222672
rect 144674 222550 144686 222602
rect 144904 222550 144916 222602
rect 144308 222478 144360 222490
rect 146700 222660 146752 222672
rect 145870 222550 145882 222602
rect 146100 222550 146112 222602
rect 145504 222478 145556 222490
rect 149092 222660 149144 222672
rect 148262 222550 148274 222602
rect 148492 222550 148504 222602
rect 146700 222478 146752 222490
rect 150288 222660 150340 222672
rect 149458 222550 149470 222602
rect 149688 222550 149700 222602
rect 149092 222478 149144 222490
rect 151484 222660 151536 222672
rect 150654 222550 150666 222602
rect 150884 222550 150896 222602
rect 150288 222478 150340 222490
rect 152680 222660 152732 222672
rect 151850 222550 151862 222602
rect 152080 222550 152092 222602
rect 151484 222478 151536 222490
rect 152680 222478 152732 222490
rect 153232 222660 153284 222672
rect 395936 222660 395988 222672
rect 153872 222550 153884 222602
rect 154102 222550 154114 222602
rect 395106 222550 395118 222602
rect 395336 222550 395348 222602
rect 153232 222478 153284 222490
rect 397132 222660 397184 222672
rect 396302 222550 396314 222602
rect 396532 222550 396544 222602
rect 395936 222478 395988 222490
rect 398328 222660 398380 222672
rect 397498 222550 397510 222602
rect 397728 222550 397740 222602
rect 397132 222478 397184 222490
rect 399524 222660 399576 222672
rect 398694 222550 398706 222602
rect 398924 222550 398936 222602
rect 398328 222478 398380 222490
rect 400720 222660 400772 222672
rect 399890 222550 399902 222602
rect 400120 222550 400132 222602
rect 399524 222478 399576 222490
rect 401916 222660 401968 222672
rect 401086 222550 401098 222602
rect 401316 222550 401328 222602
rect 400720 222478 400772 222490
rect 403112 222660 403164 222672
rect 402282 222550 402294 222602
rect 402512 222550 402524 222602
rect 401916 222478 401968 222490
rect 404308 222660 404360 222672
rect 403478 222550 403490 222602
rect 403708 222550 403720 222602
rect 403112 222478 403164 222490
rect 405504 222660 405556 222672
rect 404674 222550 404686 222602
rect 404904 222550 404916 222602
rect 404308 222478 404360 222490
rect 406700 222660 406752 222672
rect 405870 222550 405882 222602
rect 406100 222550 406112 222602
rect 405504 222478 405556 222490
rect 409092 222660 409144 222672
rect 408262 222550 408274 222602
rect 408492 222550 408504 222602
rect 406700 222478 406752 222490
rect 410288 222660 410340 222672
rect 409458 222550 409470 222602
rect 409688 222550 409700 222602
rect 409092 222478 409144 222490
rect 411484 222660 411536 222672
rect 410654 222550 410666 222602
rect 410884 222550 410896 222602
rect 410288 222478 410340 222490
rect 412680 222660 412732 222672
rect 411850 222550 411862 222602
rect 412080 222550 412092 222602
rect 411484 222478 411536 222490
rect 412680 222478 412732 222490
rect 413232 222660 413284 222672
rect 413872 222550 413884 222602
rect 414102 222550 414114 222602
rect 413232 222478 413284 222490
rect 673860 221050 673888 223664
rect 673916 220850 673944 223720
rect 673972 220650 674000 223776
rect 674028 220450 674056 223832
rect 674084 220250 674112 223888
rect 674140 220050 674168 223944
rect 674196 219850 674224 224000
rect 674252 219650 674280 224056
rect 674308 219450 674336 224112
rect 674364 219250 674392 224168
rect 674420 219050 674448 224224
rect 674476 218850 674504 224280
rect 674532 218650 674560 224336
rect 674588 218450 674616 224392
rect 674644 218250 674672 224448
rect 674700 218050 674728 224504
rect 674756 217850 674784 224560
rect 674812 217650 674840 224616
rect 674868 217450 674896 224672
rect 674924 217250 674952 224728
rect 674980 217050 675008 224784
rect 675036 216850 675064 224840
rect 675092 216650 675120 224896
rect 675148 216450 675176 224952
rect 675204 216250 675232 225008
rect 675260 216050 675288 225064
rect 675316 215850 675344 225120
rect 675372 215650 675400 225176
rect 675428 215450 675456 225232
rect 675484 215250 675512 225288
rect 675540 215050 675568 225344
rect 675652 215050 675680 439386
rect 675708 214850 675736 439510
rect 675764 214650 675792 440582
rect 675820 214450 675848 440706
rect 675876 214250 675904 441778
rect 675932 214050 675960 441902
rect 675988 213850 676016 442974
rect 676044 213650 676072 443098
rect 676100 213450 676128 444170
rect 676156 213250 676184 444294
rect 676212 213050 676240 445366
rect 676268 212850 676296 445490
rect 676324 212650 676352 446562
rect 676380 212450 676408 446686
rect 676858 446682 676870 446734
rect 677040 446682 677052 446734
rect 677540 446728 677592 446740
rect 677540 446498 677592 446510
rect 676928 446458 676980 446470
rect 676928 446228 676980 446240
rect 677470 446132 677482 446184
rect 677652 446132 677664 446184
rect 676858 445486 676870 445538
rect 677040 445486 677052 445538
rect 677540 445532 677592 445544
rect 677540 445302 677592 445314
rect 676928 445262 676980 445274
rect 676928 445032 676980 445044
rect 677470 444936 677482 444988
rect 677652 444936 677664 444988
rect 676858 444290 676870 444342
rect 677040 444290 677052 444342
rect 677540 444336 677592 444348
rect 677540 444106 677592 444118
rect 676928 444066 676980 444078
rect 676928 443836 676980 443848
rect 677470 443740 677482 443792
rect 677652 443740 677664 443792
rect 676858 443094 676870 443146
rect 677040 443094 677052 443146
rect 677540 443140 677592 443152
rect 677540 442910 677592 442922
rect 676928 442870 676980 442882
rect 676928 442640 676980 442652
rect 677470 442544 677482 442596
rect 677652 442544 677664 442596
rect 676858 441898 676870 441950
rect 677040 441898 677052 441950
rect 677540 441944 677592 441956
rect 677540 441714 677592 441726
rect 676928 441674 676980 441686
rect 676928 441444 676980 441456
rect 677470 441348 677482 441400
rect 677652 441348 677664 441400
rect 676858 440702 676870 440754
rect 677040 440702 677052 440754
rect 677540 440748 677592 440760
rect 677540 440518 677592 440530
rect 676928 440478 676980 440490
rect 676928 440248 676980 440260
rect 677470 440152 677482 440204
rect 677652 440152 677664 440204
rect 676858 439506 676870 439558
rect 677040 439506 677052 439558
rect 677540 439552 677592 439564
rect 677540 439322 677592 439334
<< via1 >>
rect 676352 708359 676404 708411
rect 676928 708260 676938 708478
rect 676938 708260 676972 708478
rect 676972 708260 676980 708478
rect 676296 708165 676348 708217
rect 677482 708196 677652 708204
rect 677482 708162 677652 708196
rect 677482 708152 677652 708162
rect 676693 707708 676753 708065
rect 677775 707708 677835 708065
rect 676356 707516 676408 707568
rect 676300 707392 676352 707444
rect 40579 604574 40587 604792
rect 40587 604574 40621 604792
rect 40621 604574 40631 604792
rect 41179 604673 41231 604725
rect 39907 604510 40077 604518
rect 39907 604476 40077 604510
rect 39907 604466 40077 604476
rect 41235 604479 41287 604531
rect 39731 604014 39791 604371
rect 40813 604014 40873 604371
rect 39967 603648 39975 603866
rect 39975 603648 40009 603866
rect 40009 603648 40019 603866
rect 40519 603864 40689 603872
rect 40519 603830 40689 603864
rect 40519 603820 40689 603830
rect 41175 603830 41227 603882
rect 40579 603378 40587 603596
rect 40587 603378 40621 603596
rect 40621 603378 40631 603596
rect 39907 603314 40077 603322
rect 39907 603280 40077 603314
rect 39907 603270 40077 603280
rect 40272 602818 40332 603175
rect 39967 602452 39975 602670
rect 39975 602452 40009 602670
rect 40009 602452 40019 602670
rect 40519 602668 40689 602676
rect 40519 602634 40689 602668
rect 40519 602624 40689 602634
rect 40579 602182 40587 602400
rect 40587 602182 40621 602400
rect 40621 602182 40631 602400
rect 39907 602118 40077 602126
rect 39907 602084 40077 602118
rect 39907 602074 40077 602084
rect 39967 601256 39975 601474
rect 39975 601256 40009 601474
rect 40009 601256 40019 601474
rect 40519 601472 40689 601480
rect 40519 601438 40689 601472
rect 40519 601428 40689 601438
rect 40579 600986 40587 601204
rect 40587 600986 40621 601204
rect 40621 600986 40631 601204
rect 39907 600922 40077 600930
rect 39907 600888 40077 600922
rect 39907 600878 40077 600888
rect 39967 600060 39975 600278
rect 39975 600060 40009 600278
rect 40009 600060 40019 600278
rect 40519 600276 40689 600284
rect 40519 600242 40689 600276
rect 40519 600232 40689 600242
rect 40579 599790 40587 600008
rect 40587 599790 40621 600008
rect 40621 599790 40631 600008
rect 39907 599726 40077 599734
rect 39907 599692 40077 599726
rect 39907 599682 40077 599692
rect 39967 598864 39975 599082
rect 39975 598864 40009 599082
rect 40009 598864 40019 599082
rect 40519 599080 40689 599088
rect 40519 599046 40689 599080
rect 40519 599036 40689 599046
rect 40579 598594 40587 598812
rect 40587 598594 40621 598812
rect 40621 598594 40631 598812
rect 39907 598530 40077 598538
rect 39907 598496 40077 598530
rect 39907 598486 40077 598496
rect 39967 597668 39975 597886
rect 39975 597668 40009 597886
rect 40009 597668 40019 597886
rect 40519 597884 40689 597892
rect 40519 597850 40689 597884
rect 40519 597840 40689 597850
rect 40601 346393 40609 346611
rect 40609 346393 40643 346611
rect 40643 346393 40653 346611
rect 41151 346492 41203 346544
rect 41231 603706 41283 603758
rect 41291 603477 41343 603529
rect 41347 603283 41399 603335
rect 39929 346329 40099 346337
rect 39929 346295 40099 346329
rect 39929 346285 40099 346295
rect 41207 346298 41259 346350
rect 41287 602634 41339 602686
rect 39989 345467 39997 345685
rect 39997 345467 40031 345685
rect 40031 345467 40041 345685
rect 40541 345683 40711 345691
rect 40541 345649 40711 345683
rect 40541 345639 40711 345649
rect 41147 345649 41199 345701
rect 40601 345197 40609 345415
rect 40609 345197 40643 345415
rect 40643 345197 40653 345415
rect 39929 345133 40099 345141
rect 39929 345099 40099 345133
rect 39929 345089 40099 345099
rect 39989 344271 39997 344489
rect 39997 344271 40031 344489
rect 40031 344271 40041 344489
rect 40541 344487 40711 344495
rect 40541 344453 40711 344487
rect 40541 344443 40711 344453
rect 40601 344001 40609 344219
rect 40609 344001 40643 344219
rect 40643 344001 40653 344219
rect 39929 343937 40099 343945
rect 39929 343903 40099 343937
rect 39929 343893 40099 343903
rect 40291 343371 40351 343728
rect 39989 343075 39997 343293
rect 39997 343075 40031 343293
rect 40031 343075 40041 343293
rect 40541 343291 40711 343299
rect 40541 343257 40711 343291
rect 40541 343247 40711 343257
rect 40601 342805 40609 343023
rect 40609 342805 40643 343023
rect 40643 342805 40653 343023
rect 39929 342741 40099 342749
rect 39929 342707 40099 342741
rect 39929 342697 40099 342707
rect 39750 342175 39810 342532
rect 40832 342175 40892 342532
rect 39989 341879 39997 342097
rect 39997 341879 40031 342097
rect 40031 341879 40041 342097
rect 40541 342095 40711 342103
rect 40541 342061 40711 342095
rect 40541 342051 40711 342061
rect 40601 341609 40609 341827
rect 40609 341609 40643 341827
rect 40643 341609 40653 341827
rect 39929 341545 40099 341553
rect 39929 341511 40099 341545
rect 39929 341501 40099 341511
rect 39989 340683 39997 340901
rect 39997 340683 40031 340901
rect 40031 340683 40041 340901
rect 40541 340899 40711 340907
rect 40541 340865 40711 340899
rect 40541 340855 40711 340865
rect 40601 340413 40609 340631
rect 40609 340413 40643 340631
rect 40643 340413 40653 340631
rect 39929 340349 40099 340357
rect 39929 340315 40099 340349
rect 39929 340305 40099 340315
rect 39989 339487 39997 339705
rect 39997 339487 40031 339705
rect 40031 339487 40041 339705
rect 40541 339703 40711 339711
rect 40541 339669 40711 339703
rect 40541 339659 40711 339669
rect 40601 339217 40609 339435
rect 40609 339217 40643 339435
rect 40643 339217 40653 339435
rect 39929 339153 40099 339161
rect 39929 339119 40099 339153
rect 39929 339109 40099 339119
rect 39989 338291 39997 338509
rect 39997 338291 40031 338509
rect 40031 338291 40041 338509
rect 40541 338507 40711 338515
rect 40541 338473 40711 338507
rect 40541 338463 40711 338473
rect 40601 338021 40609 338239
rect 40609 338021 40643 338239
rect 40643 338021 40653 338239
rect 39929 337957 40099 337965
rect 39929 337923 40099 337957
rect 39929 337913 40099 337923
rect 39989 337095 39997 337313
rect 39997 337095 40031 337313
rect 40031 337095 40041 337313
rect 40541 337311 40711 337319
rect 40541 337277 40711 337311
rect 40541 337267 40711 337277
rect 40601 336825 40609 337043
rect 40609 336825 40643 337043
rect 40643 336825 40653 337043
rect 39929 336761 40099 336769
rect 39929 336727 40099 336761
rect 39929 336717 40099 336727
rect 39989 335899 39997 336117
rect 39997 335899 40031 336117
rect 40031 335899 40041 336117
rect 40541 336115 40711 336123
rect 40541 336081 40711 336115
rect 40541 336071 40711 336081
rect 40601 335629 40609 335847
rect 40609 335629 40643 335847
rect 40643 335629 40653 335847
rect 39929 335565 40099 335573
rect 39929 335531 40099 335565
rect 39929 335521 40099 335531
rect 39989 334703 39997 334921
rect 39997 334703 40031 334921
rect 40031 334703 40041 334921
rect 40541 334919 40711 334927
rect 40541 334885 40711 334919
rect 40541 334875 40711 334885
rect 41203 345525 41255 345577
rect 41263 345296 41315 345348
rect 41343 602510 41395 602562
rect 41403 602281 41455 602333
rect 41459 602087 41511 602139
rect 41319 345102 41371 345154
rect 41399 601438 41451 601490
rect 41259 344453 41311 344505
rect 41315 344329 41367 344381
rect 41375 344100 41427 344152
rect 41455 601314 41507 601366
rect 41515 601085 41567 601137
rect 41571 600891 41623 600943
rect 41431 343906 41483 343958
rect 41511 600242 41563 600294
rect 41371 343257 41423 343309
rect 41427 343133 41479 343185
rect 41487 342904 41539 342956
rect 41567 600118 41619 600170
rect 41627 599889 41679 599941
rect 41683 599695 41735 599747
rect 41543 342710 41595 342762
rect 41623 599046 41675 599098
rect 41483 342061 41535 342113
rect 41539 341937 41591 341989
rect 41599 341708 41651 341760
rect 41679 598922 41731 598974
rect 41739 598693 41791 598745
rect 41795 598499 41847 598551
rect 41655 341514 41707 341566
rect 41735 597850 41787 597902
rect 41595 340865 41647 340917
rect 41651 340741 41703 340793
rect 41711 340512 41763 340564
rect 41791 597726 41843 597778
rect 676870 707550 677040 707558
rect 676870 707516 677040 707550
rect 676870 707506 677040 707516
rect 677540 707334 677550 707552
rect 677550 707334 677584 707552
rect 677584 707334 677592 707552
rect 677234 706512 677294 706869
rect 676352 447535 676404 447587
rect 676928 447436 676938 447654
rect 676938 447436 676972 447654
rect 676972 447436 676980 447654
rect 676296 447341 676348 447393
rect 677482 447372 677652 447380
rect 677482 447338 677652 447372
rect 677482 447328 677652 447338
rect 677226 446899 677286 447256
rect 676356 446692 676408 446744
rect 676300 446568 676352 446620
rect 676240 446339 676292 446391
rect 676184 446145 676236 446197
rect 676244 445496 676296 445548
rect 676188 445372 676240 445424
rect 676128 445143 676180 445195
rect 676072 444949 676124 445001
rect 676132 444300 676184 444352
rect 676076 444176 676128 444228
rect 676016 443947 676068 443999
rect 675960 443753 676012 443805
rect 676020 443104 676072 443156
rect 675964 442980 676016 443032
rect 675904 442751 675956 442803
rect 675848 442557 675900 442609
rect 675908 441908 675960 441960
rect 675852 441784 675904 441836
rect 675792 441555 675844 441607
rect 675736 441361 675788 441413
rect 675796 440712 675848 440764
rect 675740 440588 675792 440640
rect 675680 440359 675732 440411
rect 675624 440165 675676 440217
rect 675684 439516 675736 439568
rect 675628 439392 675680 439444
rect 41767 340318 41819 340370
rect 41707 339669 41759 339721
rect 41763 339545 41815 339597
rect 41823 339316 41875 339368
rect 41879 339122 41931 339174
rect 41819 338473 41871 338525
rect 41875 338349 41927 338401
rect 41935 338120 41987 338172
rect 41991 337926 42043 337978
rect 41931 337277 41983 337329
rect 41987 337153 42039 337205
rect 42047 336900 42099 336952
rect 42103 336730 42155 336782
rect 42043 336081 42095 336133
rect 42099 335957 42151 336009
rect 42159 335728 42211 335780
rect 42215 335534 42267 335586
rect 42155 334885 42207 334937
rect 42211 334761 42263 334813
rect 134104 225288 134156 225340
rect 134947 225292 134999 225344
rect 394104 225316 394156 225368
rect 394947 225320 394999 225372
rect 135176 225232 135228 225284
rect 135949 225236 136001 225288
rect 395176 225260 395228 225312
rect 395949 225264 396001 225316
rect 135300 225176 135352 225228
rect 136143 225180 136195 225232
rect 395300 225204 395352 225256
rect 396143 225208 396195 225260
rect 136372 225120 136424 225172
rect 137145 225124 137197 225176
rect 396372 225148 396424 225200
rect 397145 225152 397197 225204
rect 136496 225064 136548 225116
rect 137339 225068 137391 225120
rect 396496 225092 396548 225144
rect 397339 225096 397391 225148
rect 137568 225008 137620 225060
rect 138341 225012 138393 225064
rect 397568 225036 397620 225088
rect 398341 225040 398393 225092
rect 137692 224952 137744 225004
rect 138535 224956 138587 225008
rect 397692 224980 397744 225032
rect 398535 224984 398587 225036
rect 138764 224896 138816 224948
rect 139537 224900 139589 224952
rect 398764 224924 398816 224976
rect 399537 224928 399589 224980
rect 138888 224840 138940 224892
rect 139731 224844 139783 224896
rect 398888 224868 398940 224920
rect 399731 224872 399783 224924
rect 139960 224784 140012 224836
rect 140733 224788 140785 224840
rect 399960 224812 400012 224864
rect 400733 224816 400785 224868
rect 140084 224728 140136 224780
rect 140903 224732 140955 224784
rect 400084 224756 400136 224808
rect 400903 224760 400955 224812
rect 141156 224672 141208 224724
rect 141929 224676 141981 224728
rect 401156 224700 401208 224752
rect 401929 224704 401981 224756
rect 141280 224616 141332 224668
rect 142123 224620 142175 224672
rect 401280 224644 401332 224696
rect 402123 224648 402175 224700
rect 142352 224560 142404 224612
rect 143125 224564 143177 224616
rect 402352 224588 402404 224640
rect 403125 224592 403177 224644
rect 142476 224504 142528 224556
rect 143295 224508 143347 224560
rect 402476 224532 402528 224584
rect 403295 224536 403347 224588
rect 143548 224448 143600 224500
rect 144321 224452 144373 224504
rect 403548 224476 403600 224528
rect 404321 224480 404373 224532
rect 143672 224392 143724 224444
rect 144515 224396 144567 224448
rect 403672 224420 403724 224472
rect 404515 224424 404567 224476
rect 144744 224336 144796 224388
rect 145517 224340 145569 224392
rect 404744 224364 404796 224416
rect 405517 224368 405569 224420
rect 144868 224280 144920 224332
rect 145711 224284 145763 224336
rect 404868 224308 404920 224360
rect 405711 224312 405763 224364
rect 145940 224224 145992 224276
rect 146713 224228 146765 224280
rect 405940 224252 405992 224304
rect 406713 224256 406765 224308
rect 147260 224168 147312 224220
rect 148103 224172 148155 224224
rect 407260 224196 407312 224248
rect 408103 224200 408155 224252
rect 148332 224112 148384 224164
rect 149105 224116 149157 224168
rect 408332 224140 408384 224192
rect 409105 224144 409157 224196
rect 148456 224056 148508 224108
rect 149299 224060 149351 224112
rect 408456 224084 408508 224136
rect 409299 224088 409351 224140
rect 149528 224000 149580 224052
rect 150301 224004 150353 224056
rect 409528 224028 409580 224080
rect 410301 224032 410353 224084
rect 149652 223944 149704 223996
rect 150471 223948 150523 224000
rect 409652 223972 409704 224024
rect 410471 223976 410523 224028
rect 150724 223888 150776 223940
rect 151497 223892 151549 223944
rect 410724 223916 410776 223968
rect 411497 223920 411549 223972
rect 150848 223832 150900 223884
rect 151691 223836 151743 223888
rect 410848 223860 410900 223912
rect 411691 223864 411743 223916
rect 151920 223776 151972 223828
rect 152693 223780 152745 223832
rect 411920 223804 411972 223856
rect 412693 223808 412745 223860
rect 152044 223720 152096 223772
rect 152863 223724 152915 223776
rect 412044 223748 412096 223800
rect 412863 223752 412915 223804
rect 153116 223664 153168 223716
rect 153889 223668 153941 223720
rect 413116 223692 413168 223744
rect 413889 223696 413941 223748
rect 153240 223608 153292 223660
rect 154083 223612 154135 223664
rect 413240 223636 413292 223688
rect 414083 223640 414135 223692
rect 147395 223397 147752 223457
rect 406226 223390 406583 223450
rect 134094 223102 134104 223272
rect 134104 223102 134138 223272
rect 134138 223102 134146 223272
rect 134848 223204 135066 223214
rect 134848 223170 135066 223204
rect 134848 223162 135066 223170
rect 135290 223102 135300 223272
rect 135300 223102 135334 223272
rect 135334 223102 135342 223272
rect 136044 223204 136262 223214
rect 136044 223170 136262 223204
rect 136044 223162 136262 223170
rect 136486 223102 136496 223272
rect 136496 223102 136530 223272
rect 136530 223102 136538 223272
rect 137240 223204 137458 223214
rect 137240 223170 137458 223204
rect 137240 223162 137458 223170
rect 137682 223102 137692 223272
rect 137692 223102 137726 223272
rect 137726 223102 137734 223272
rect 138436 223204 138654 223214
rect 138436 223170 138654 223204
rect 138436 223162 138654 223170
rect 138878 223102 138888 223272
rect 138888 223102 138922 223272
rect 138922 223102 138930 223272
rect 139632 223204 139850 223214
rect 139632 223170 139850 223204
rect 139632 223162 139850 223170
rect 140074 223102 140084 223272
rect 140084 223102 140118 223272
rect 140118 223102 140126 223272
rect 140828 223204 141046 223214
rect 140828 223170 141046 223204
rect 140828 223162 141046 223170
rect 141270 223102 141280 223272
rect 141280 223102 141314 223272
rect 141314 223102 141322 223272
rect 142024 223204 142242 223214
rect 142024 223170 142242 223204
rect 142024 223162 142242 223170
rect 142466 223102 142476 223272
rect 142476 223102 142510 223272
rect 142510 223102 142518 223272
rect 143220 223204 143438 223214
rect 143220 223170 143438 223204
rect 143220 223162 143438 223170
rect 143662 223102 143672 223272
rect 143672 223102 143706 223272
rect 143706 223102 143714 223272
rect 144416 223204 144634 223214
rect 144416 223170 144634 223204
rect 144416 223162 144634 223170
rect 144858 223102 144868 223272
rect 144868 223102 144902 223272
rect 144902 223102 144910 223272
rect 145612 223204 145830 223214
rect 145612 223170 145830 223204
rect 145612 223162 145830 223170
rect 147250 223102 147260 223272
rect 147260 223102 147294 223272
rect 147294 223102 147302 223272
rect 148004 223204 148222 223214
rect 148004 223170 148222 223204
rect 148004 223162 148222 223170
rect 148446 223102 148456 223272
rect 148456 223102 148490 223272
rect 148490 223102 148498 223272
rect 149200 223204 149418 223214
rect 149200 223170 149418 223204
rect 149200 223162 149418 223170
rect 149642 223102 149652 223272
rect 149652 223102 149686 223272
rect 149686 223102 149694 223272
rect 150396 223204 150614 223214
rect 150396 223170 150614 223204
rect 150396 223162 150614 223170
rect 150838 223102 150848 223272
rect 150848 223102 150882 223272
rect 150882 223102 150890 223272
rect 151592 223204 151810 223214
rect 151592 223170 151810 223204
rect 151592 223162 151810 223170
rect 152034 223102 152044 223272
rect 152044 223102 152078 223272
rect 152078 223102 152086 223272
rect 152788 223204 153006 223214
rect 152788 223170 153006 223204
rect 152788 223162 153006 223170
rect 153230 223102 153240 223272
rect 153240 223102 153274 223272
rect 153274 223102 153282 223272
rect 153984 223204 154202 223214
rect 153984 223170 154202 223204
rect 153984 223162 154202 223170
rect 394094 223102 394104 223272
rect 394104 223102 394138 223272
rect 394138 223102 394146 223272
rect 394848 223204 395066 223214
rect 394848 223170 395066 223204
rect 394848 223162 395066 223170
rect 395290 223102 395300 223272
rect 395300 223102 395334 223272
rect 395334 223102 395342 223272
rect 396044 223204 396262 223214
rect 396044 223170 396262 223204
rect 396044 223162 396262 223170
rect 396486 223102 396496 223272
rect 396496 223102 396530 223272
rect 396530 223102 396538 223272
rect 397240 223204 397458 223214
rect 397240 223170 397458 223204
rect 397240 223162 397458 223170
rect 397682 223102 397692 223272
rect 397692 223102 397726 223272
rect 397726 223102 397734 223272
rect 398436 223204 398654 223214
rect 398436 223170 398654 223204
rect 398436 223162 398654 223170
rect 398878 223102 398888 223272
rect 398888 223102 398922 223272
rect 398922 223102 398930 223272
rect 399632 223204 399850 223214
rect 399632 223170 399850 223204
rect 399632 223162 399850 223170
rect 400074 223102 400084 223272
rect 400084 223102 400118 223272
rect 400118 223102 400126 223272
rect 400828 223204 401046 223214
rect 400828 223170 401046 223204
rect 400828 223162 401046 223170
rect 401270 223102 401280 223272
rect 401280 223102 401314 223272
rect 401314 223102 401322 223272
rect 402024 223204 402242 223214
rect 402024 223170 402242 223204
rect 402024 223162 402242 223170
rect 402466 223102 402476 223272
rect 402476 223102 402510 223272
rect 402510 223102 402518 223272
rect 403220 223204 403438 223214
rect 403220 223170 403438 223204
rect 403220 223162 403438 223170
rect 403662 223102 403672 223272
rect 403672 223102 403706 223272
rect 403706 223102 403714 223272
rect 404416 223204 404634 223214
rect 404416 223170 404634 223204
rect 404416 223162 404634 223170
rect 404858 223102 404868 223272
rect 404868 223102 404902 223272
rect 404902 223102 404910 223272
rect 405612 223204 405830 223214
rect 405612 223170 405830 223204
rect 405612 223162 405830 223170
rect 407250 223102 407260 223272
rect 407260 223102 407294 223272
rect 407294 223102 407302 223272
rect 408004 223204 408222 223214
rect 408004 223170 408222 223204
rect 408004 223162 408222 223170
rect 408446 223102 408456 223272
rect 408456 223102 408490 223272
rect 408490 223102 408498 223272
rect 409200 223204 409418 223214
rect 409200 223170 409418 223204
rect 409200 223162 409418 223170
rect 409642 223102 409652 223272
rect 409652 223102 409686 223272
rect 409686 223102 409694 223272
rect 410396 223204 410614 223214
rect 410396 223170 410614 223204
rect 410396 223162 410614 223170
rect 410838 223102 410848 223272
rect 410848 223102 410882 223272
rect 410882 223102 410890 223272
rect 411592 223204 411810 223214
rect 411592 223170 411810 223204
rect 411592 223162 411810 223170
rect 412034 223102 412044 223272
rect 412044 223102 412078 223272
rect 412078 223102 412086 223272
rect 412788 223204 413006 223214
rect 412788 223170 413006 223204
rect 412788 223162 413006 223170
rect 413230 223102 413240 223272
rect 413240 223102 413274 223272
rect 413274 223102 413282 223272
rect 413984 223204 414202 223214
rect 413984 223170 414202 223204
rect 413984 223162 414202 223170
rect 146199 222856 146556 222916
rect 405030 222849 405387 222909
rect 135118 222592 135336 222602
rect 135118 222558 135336 222592
rect 135118 222550 135336 222558
rect 135936 222490 135946 222660
rect 135946 222490 135980 222660
rect 135980 222490 135988 222660
rect 136314 222592 136532 222602
rect 136314 222558 136532 222592
rect 136314 222550 136532 222558
rect 137132 222490 137142 222660
rect 137142 222490 137176 222660
rect 137176 222490 137184 222660
rect 137510 222592 137728 222602
rect 137510 222558 137728 222592
rect 137510 222550 137728 222558
rect 138328 222490 138338 222660
rect 138338 222490 138372 222660
rect 138372 222490 138380 222660
rect 138706 222592 138924 222602
rect 138706 222558 138924 222592
rect 138706 222550 138924 222558
rect 139524 222490 139534 222660
rect 139534 222490 139568 222660
rect 139568 222490 139576 222660
rect 139902 222592 140120 222602
rect 139902 222558 140120 222592
rect 139902 222550 140120 222558
rect 140720 222490 140730 222660
rect 140730 222490 140764 222660
rect 140764 222490 140772 222660
rect 141098 222592 141316 222602
rect 141098 222558 141316 222592
rect 141098 222550 141316 222558
rect 141916 222490 141926 222660
rect 141926 222490 141960 222660
rect 141960 222490 141968 222660
rect 142294 222592 142512 222602
rect 142294 222558 142512 222592
rect 142294 222550 142512 222558
rect 143112 222490 143122 222660
rect 143122 222490 143156 222660
rect 143156 222490 143164 222660
rect 143490 222592 143708 222602
rect 143490 222558 143708 222592
rect 143490 222550 143708 222558
rect 144308 222490 144318 222660
rect 144318 222490 144352 222660
rect 144352 222490 144360 222660
rect 144686 222592 144904 222602
rect 144686 222558 144904 222592
rect 144686 222550 144904 222558
rect 145504 222490 145514 222660
rect 145514 222490 145548 222660
rect 145548 222490 145556 222660
rect 145882 222592 146100 222602
rect 145882 222558 146100 222592
rect 145882 222550 146100 222558
rect 146700 222490 146710 222660
rect 146710 222490 146744 222660
rect 146744 222490 146752 222660
rect 148274 222592 148492 222602
rect 148274 222558 148492 222592
rect 148274 222550 148492 222558
rect 149092 222490 149102 222660
rect 149102 222490 149136 222660
rect 149136 222490 149144 222660
rect 149470 222592 149688 222602
rect 149470 222558 149688 222592
rect 149470 222550 149688 222558
rect 150288 222490 150298 222660
rect 150298 222490 150332 222660
rect 150332 222490 150340 222660
rect 150666 222592 150884 222602
rect 150666 222558 150884 222592
rect 150666 222550 150884 222558
rect 151484 222490 151494 222660
rect 151494 222490 151528 222660
rect 151528 222490 151536 222660
rect 151862 222592 152080 222602
rect 151862 222558 152080 222592
rect 151862 222550 152080 222558
rect 152680 222490 152690 222660
rect 152690 222490 152724 222660
rect 152724 222490 152732 222660
rect 153232 222490 153240 222660
rect 153240 222490 153274 222660
rect 153274 222490 153284 222660
rect 153884 222592 154102 222602
rect 153884 222558 154102 222592
rect 153884 222550 154102 222558
rect 395118 222592 395336 222602
rect 395118 222558 395336 222592
rect 395118 222550 395336 222558
rect 395936 222490 395946 222660
rect 395946 222490 395980 222660
rect 395980 222490 395988 222660
rect 396314 222592 396532 222602
rect 396314 222558 396532 222592
rect 396314 222550 396532 222558
rect 397132 222490 397142 222660
rect 397142 222490 397176 222660
rect 397176 222490 397184 222660
rect 397510 222592 397728 222602
rect 397510 222558 397728 222592
rect 397510 222550 397728 222558
rect 398328 222490 398338 222660
rect 398338 222490 398372 222660
rect 398372 222490 398380 222660
rect 398706 222592 398924 222602
rect 398706 222558 398924 222592
rect 398706 222550 398924 222558
rect 399524 222490 399534 222660
rect 399534 222490 399568 222660
rect 399568 222490 399576 222660
rect 399902 222592 400120 222602
rect 399902 222558 400120 222592
rect 399902 222550 400120 222558
rect 400720 222490 400730 222660
rect 400730 222490 400764 222660
rect 400764 222490 400772 222660
rect 401098 222592 401316 222602
rect 401098 222558 401316 222592
rect 401098 222550 401316 222558
rect 401916 222490 401926 222660
rect 401926 222490 401960 222660
rect 401960 222490 401968 222660
rect 402294 222592 402512 222602
rect 402294 222558 402512 222592
rect 402294 222550 402512 222558
rect 403112 222490 403122 222660
rect 403122 222490 403156 222660
rect 403156 222490 403164 222660
rect 403490 222592 403708 222602
rect 403490 222558 403708 222592
rect 403490 222550 403708 222558
rect 404308 222490 404318 222660
rect 404318 222490 404352 222660
rect 404352 222490 404360 222660
rect 404686 222592 404904 222602
rect 404686 222558 404904 222592
rect 404686 222550 404904 222558
rect 405504 222490 405514 222660
rect 405514 222490 405548 222660
rect 405548 222490 405556 222660
rect 405882 222592 406100 222602
rect 405882 222558 406100 222592
rect 405882 222550 406100 222558
rect 406700 222490 406710 222660
rect 406710 222490 406744 222660
rect 406744 222490 406752 222660
rect 408274 222592 408492 222602
rect 408274 222558 408492 222592
rect 408274 222550 408492 222558
rect 409092 222490 409102 222660
rect 409102 222490 409136 222660
rect 409136 222490 409144 222660
rect 409470 222592 409688 222602
rect 409470 222558 409688 222592
rect 409470 222550 409688 222558
rect 410288 222490 410298 222660
rect 410298 222490 410332 222660
rect 410332 222490 410340 222660
rect 410666 222592 410884 222602
rect 410666 222558 410884 222592
rect 410666 222550 410884 222558
rect 411484 222490 411494 222660
rect 411494 222490 411528 222660
rect 411528 222490 411536 222660
rect 411862 222592 412080 222602
rect 411862 222558 412080 222592
rect 411862 222550 412080 222558
rect 412680 222490 412690 222660
rect 412690 222490 412724 222660
rect 412724 222490 412732 222660
rect 413232 222490 413240 222660
rect 413240 222490 413274 222660
rect 413274 222490 413284 222660
rect 413884 222592 414102 222602
rect 413884 222558 414102 222592
rect 413884 222550 414102 222558
rect 147395 222315 147752 222375
rect 406226 222308 406583 222368
rect 676870 446726 677040 446734
rect 676870 446692 677040 446726
rect 676870 446682 677040 446692
rect 677540 446510 677550 446728
rect 677550 446510 677584 446728
rect 677584 446510 677592 446728
rect 676928 446240 676938 446458
rect 676938 446240 676972 446458
rect 676972 446240 676980 446458
rect 677482 446176 677652 446184
rect 677482 446142 677652 446176
rect 677482 446132 677652 446142
rect 676685 445703 676745 446060
rect 677767 445703 677827 446060
rect 676870 445530 677040 445538
rect 676870 445496 677040 445530
rect 676870 445486 677040 445496
rect 677540 445314 677550 445532
rect 677550 445314 677584 445532
rect 677584 445314 677592 445532
rect 676928 445044 676938 445262
rect 676938 445044 676972 445262
rect 676972 445044 676980 445262
rect 677482 444980 677652 444988
rect 677482 444946 677652 444980
rect 677482 444936 677652 444946
rect 676870 444334 677040 444342
rect 676870 444300 677040 444334
rect 676870 444290 677040 444300
rect 677540 444118 677550 444336
rect 677550 444118 677584 444336
rect 677584 444118 677592 444336
rect 676928 443848 676938 444066
rect 676938 443848 676972 444066
rect 676972 443848 676980 444066
rect 677482 443784 677652 443792
rect 677482 443750 677652 443784
rect 677482 443740 677652 443750
rect 676870 443138 677040 443146
rect 676870 443104 677040 443138
rect 676870 443094 677040 443104
rect 677540 442922 677550 443140
rect 677550 442922 677584 443140
rect 677584 442922 677592 443140
rect 676928 442652 676938 442870
rect 676938 442652 676972 442870
rect 676972 442652 676980 442870
rect 677482 442588 677652 442596
rect 677482 442554 677652 442588
rect 677482 442544 677652 442554
rect 676870 441942 677040 441950
rect 676870 441908 677040 441942
rect 676870 441898 677040 441908
rect 677540 441726 677550 441944
rect 677550 441726 677584 441944
rect 677584 441726 677592 441944
rect 676928 441456 676938 441674
rect 676938 441456 676972 441674
rect 676972 441456 676980 441674
rect 677482 441392 677652 441400
rect 677482 441358 677652 441392
rect 677482 441348 677652 441358
rect 676870 440746 677040 440754
rect 676870 440712 677040 440746
rect 676870 440702 677040 440712
rect 677540 440530 677550 440748
rect 677550 440530 677584 440748
rect 677584 440530 677592 440748
rect 676928 440260 676938 440478
rect 676938 440260 676972 440478
rect 676972 440260 676980 440478
rect 677482 440196 677652 440204
rect 677482 440162 677652 440196
rect 677482 440152 677652 440162
rect 676870 439550 677040 439558
rect 676870 439516 677040 439550
rect 676870 439506 677040 439516
rect 677540 439334 677550 439552
rect 677550 439334 677584 439552
rect 677584 439334 677592 439552
<< metal2 >>
rect 676346 708387 676352 708411
rect 676262 708359 676352 708387
rect 676404 708387 676410 708411
rect 676922 708387 676928 708478
rect 676404 708359 676928 708387
rect 676922 708260 676928 708359
rect 676980 708260 676986 708478
rect 676290 708193 676296 708217
rect 676262 708165 676296 708193
rect 676348 708193 676354 708217
rect 677482 708204 677652 708210
rect 676348 708165 677482 708193
rect 677482 708146 677652 708152
rect 676681 708065 676767 708073
rect 676681 707708 676693 708065
rect 676753 707708 676767 708065
rect 676681 707700 676767 707708
rect 677766 708065 677852 708073
rect 677766 707708 677775 708065
rect 677835 707708 677852 708065
rect 677766 707700 677852 707708
rect 676350 707544 676356 707568
rect 676262 707516 676356 707544
rect 676408 707544 676414 707568
rect 676870 707558 677040 707564
rect 676408 707516 676870 707544
rect 676870 707500 677040 707506
rect 676294 707420 676300 707444
rect 676262 707392 676300 707420
rect 676352 707420 676358 707444
rect 677534 707420 677540 707552
rect 676352 707392 677540 707420
rect 677534 707334 677540 707392
rect 677592 707334 677598 707552
rect 677220 706869 677306 706877
rect 677220 706512 677234 706869
rect 677294 706512 677306 706869
rect 677220 706504 677306 706512
rect 40573 604574 40579 604792
rect 40631 604701 40637 604792
rect 41173 604701 41179 604725
rect 40631 604673 41179 604701
rect 41231 604701 41237 604725
rect 41231 604673 41860 604701
rect 40631 604574 40637 604673
rect 39907 604518 40077 604524
rect 41229 604507 41235 604531
rect 40077 604479 41235 604507
rect 41287 604507 41293 604531
rect 41287 604479 41860 604507
rect 39907 604460 40077 604466
rect 39714 604371 39800 604379
rect 39714 604014 39731 604371
rect 39791 604014 39800 604371
rect 39714 604006 39800 604014
rect 40799 604371 40885 604379
rect 40799 604014 40813 604371
rect 40873 604014 40885 604371
rect 40799 604006 40885 604014
rect 40519 603872 40689 603878
rect 39961 603648 39967 603866
rect 40019 603734 40025 603866
rect 41169 603858 41175 603882
rect 40689 603830 41175 603858
rect 41227 603858 41233 603882
rect 41227 603830 41860 603858
rect 40519 603814 40689 603820
rect 41225 603734 41231 603758
rect 40019 603706 41231 603734
rect 41283 603734 41289 603758
rect 41283 603706 41860 603734
rect 40019 603648 40025 603706
rect 40573 603378 40579 603596
rect 40631 603505 40637 603596
rect 41285 603505 41291 603529
rect 40631 603477 41291 603505
rect 41343 603505 41349 603529
rect 41343 603477 41860 603505
rect 40631 603378 40637 603477
rect 39907 603322 40077 603328
rect 41341 603311 41347 603335
rect 40077 603283 41347 603311
rect 41399 603311 41405 603335
rect 41399 603283 41860 603311
rect 39907 603264 40077 603270
rect 40260 603175 40346 603183
rect 40260 602818 40272 603175
rect 40332 602818 40346 603175
rect 40260 602810 40346 602818
rect 40519 602676 40689 602682
rect 39961 602452 39967 602670
rect 40019 602538 40025 602670
rect 41281 602662 41287 602686
rect 40689 602634 41287 602662
rect 41339 602662 41345 602686
rect 41339 602634 41860 602662
rect 40519 602618 40689 602624
rect 41337 602538 41343 602562
rect 40019 602510 41343 602538
rect 41395 602538 41401 602562
rect 41395 602510 41860 602538
rect 40019 602452 40025 602510
rect 40573 602182 40579 602400
rect 40631 602309 40637 602400
rect 41397 602309 41403 602333
rect 40631 602281 41403 602309
rect 41455 602309 41461 602333
rect 41455 602281 41860 602309
rect 40631 602182 40637 602281
rect 39907 602126 40077 602132
rect 41453 602115 41459 602139
rect 40077 602087 41459 602115
rect 41511 602115 41517 602139
rect 41511 602087 41860 602115
rect 39907 602068 40077 602074
rect 40519 601480 40689 601486
rect 39961 601256 39967 601474
rect 40019 601342 40025 601474
rect 41393 601466 41399 601490
rect 40689 601438 41399 601466
rect 41451 601466 41457 601490
rect 41451 601438 41860 601466
rect 40519 601422 40689 601428
rect 41449 601342 41455 601366
rect 40019 601314 41455 601342
rect 41507 601342 41513 601366
rect 41507 601314 41860 601342
rect 40019 601256 40025 601314
rect 40573 600986 40579 601204
rect 40631 601113 40637 601204
rect 41509 601113 41515 601137
rect 40631 601085 41515 601113
rect 41567 601113 41573 601137
rect 41567 601085 41860 601113
rect 40631 600986 40637 601085
rect 39907 600930 40077 600936
rect 41565 600919 41571 600943
rect 40077 600891 41571 600919
rect 41623 600919 41629 600943
rect 41623 600891 41860 600919
rect 39907 600872 40077 600878
rect 40519 600284 40689 600290
rect 39961 600060 39967 600278
rect 40019 600146 40025 600278
rect 41505 600270 41511 600294
rect 40689 600242 41511 600270
rect 41563 600270 41569 600294
rect 41563 600242 41860 600270
rect 40519 600226 40689 600232
rect 41561 600146 41567 600170
rect 40019 600118 41567 600146
rect 41619 600146 41625 600170
rect 41619 600118 41860 600146
rect 40019 600060 40025 600118
rect 40573 599790 40579 600008
rect 40631 599917 40637 600008
rect 41621 599917 41627 599941
rect 40631 599889 41627 599917
rect 41679 599917 41685 599941
rect 41679 599889 41860 599917
rect 40631 599790 40637 599889
rect 39907 599734 40077 599740
rect 41677 599723 41683 599747
rect 40077 599695 41683 599723
rect 41735 599723 41741 599747
rect 41735 599695 41860 599723
rect 39907 599676 40077 599682
rect 40519 599088 40689 599094
rect 39961 598864 39967 599082
rect 40019 598950 40025 599082
rect 41617 599074 41623 599098
rect 40689 599046 41623 599074
rect 41675 599074 41681 599098
rect 41675 599046 41860 599074
rect 40519 599030 40689 599036
rect 41673 598950 41679 598974
rect 40019 598922 41679 598950
rect 41731 598950 41737 598974
rect 41731 598922 41860 598950
rect 40019 598864 40025 598922
rect 40573 598594 40579 598812
rect 40631 598721 40637 598812
rect 41733 598721 41739 598745
rect 40631 598693 41739 598721
rect 41791 598721 41797 598745
rect 41791 598693 41860 598721
rect 40631 598594 40637 598693
rect 39907 598538 40077 598544
rect 41789 598527 41795 598551
rect 40077 598499 41795 598527
rect 41847 598527 41853 598551
rect 41847 598499 41860 598527
rect 39907 598480 40077 598486
rect 40519 597892 40689 597898
rect 39961 597668 39967 597886
rect 40019 597754 40025 597886
rect 41729 597878 41735 597902
rect 40689 597850 41735 597878
rect 41787 597878 41793 597902
rect 41787 597850 41860 597878
rect 40519 597834 40689 597840
rect 41785 597754 41791 597778
rect 40019 597726 41791 597754
rect 41843 597754 41849 597778
rect 41843 597726 41860 597754
rect 40019 597668 40025 597726
rect 676346 447563 676352 447587
rect 675590 447535 676352 447563
rect 676404 447563 676410 447587
rect 676922 447563 676928 447654
rect 676404 447535 676928 447563
rect 676922 447436 676928 447535
rect 676980 447436 676986 447654
rect 676290 447369 676296 447393
rect 675590 447341 676296 447369
rect 676348 447369 676354 447393
rect 677482 447380 677652 447386
rect 676348 447341 677482 447369
rect 677482 447322 677652 447328
rect 677212 447256 677298 447264
rect 677212 446899 677226 447256
rect 677286 446899 677298 447256
rect 677212 446891 677298 446899
rect 676350 446720 676356 446744
rect 675590 446692 676356 446720
rect 676408 446720 676414 446744
rect 676870 446734 677040 446740
rect 676408 446692 676870 446720
rect 676870 446676 677040 446682
rect 676294 446596 676300 446620
rect 675590 446568 676300 446596
rect 676352 446596 676358 446620
rect 677534 446596 677540 446728
rect 676352 446568 677540 446596
rect 677534 446510 677540 446568
rect 677592 446510 677598 446728
rect 676234 446367 676240 446391
rect 675590 446339 676240 446367
rect 676292 446367 676298 446391
rect 676922 446367 676928 446458
rect 676292 446339 676928 446367
rect 676922 446240 676928 446339
rect 676980 446240 676986 446458
rect 676178 446173 676184 446197
rect 675590 446145 676184 446173
rect 676236 446173 676242 446197
rect 677482 446184 677652 446190
rect 676236 446145 677482 446173
rect 677482 446126 677652 446132
rect 676673 446060 676759 446068
rect 676673 445703 676685 446060
rect 676745 445703 676759 446060
rect 676673 445695 676759 445703
rect 677758 446060 677844 446068
rect 677758 445703 677767 446060
rect 677827 445703 677844 446060
rect 677758 445695 677844 445703
rect 676238 445524 676244 445548
rect 675590 445496 676244 445524
rect 676296 445524 676302 445548
rect 676870 445538 677040 445544
rect 676296 445496 676870 445524
rect 676870 445480 677040 445486
rect 676182 445400 676188 445424
rect 675590 445372 676188 445400
rect 676240 445400 676246 445424
rect 677534 445400 677540 445532
rect 676240 445372 677540 445400
rect 677534 445314 677540 445372
rect 677592 445314 677598 445532
rect 676122 445171 676128 445195
rect 675590 445143 676128 445171
rect 676180 445171 676186 445195
rect 676922 445171 676928 445262
rect 676180 445143 676928 445171
rect 676922 445044 676928 445143
rect 676980 445044 676986 445262
rect 676066 444977 676072 445001
rect 675590 444949 676072 444977
rect 676124 444977 676130 445001
rect 677482 444988 677652 444994
rect 676124 444949 677482 444977
rect 677482 444930 677652 444936
rect 676126 444328 676132 444352
rect 675590 444300 676132 444328
rect 676184 444328 676190 444352
rect 676870 444342 677040 444348
rect 676184 444300 676870 444328
rect 676870 444284 677040 444290
rect 676070 444204 676076 444228
rect 675590 444176 676076 444204
rect 676128 444204 676134 444228
rect 677534 444204 677540 444336
rect 676128 444176 677540 444204
rect 677534 444118 677540 444176
rect 677592 444118 677598 444336
rect 676010 443975 676016 443999
rect 675590 443947 676016 443975
rect 676068 443975 676074 443999
rect 676922 443975 676928 444066
rect 676068 443947 676928 443975
rect 676922 443848 676928 443947
rect 676980 443848 676986 444066
rect 675954 443781 675960 443805
rect 675590 443753 675960 443781
rect 676012 443781 676018 443805
rect 677482 443792 677652 443798
rect 676012 443753 677482 443781
rect 677482 443734 677652 443740
rect 676014 443132 676020 443156
rect 675590 443104 676020 443132
rect 676072 443132 676078 443156
rect 676870 443146 677040 443152
rect 676072 443104 676870 443132
rect 676870 443088 677040 443094
rect 675958 443008 675964 443032
rect 675590 442980 675964 443008
rect 676016 443008 676022 443032
rect 677534 443008 677540 443140
rect 676016 442980 677540 443008
rect 677534 442922 677540 442980
rect 677592 442922 677598 443140
rect 675898 442779 675904 442803
rect 675590 442751 675904 442779
rect 675956 442779 675962 442803
rect 676922 442779 676928 442870
rect 675956 442751 676928 442779
rect 676922 442652 676928 442751
rect 676980 442652 676986 442870
rect 675842 442585 675848 442609
rect 675590 442557 675848 442585
rect 675900 442585 675906 442609
rect 677482 442596 677652 442602
rect 675900 442557 677482 442585
rect 677482 442538 677652 442544
rect 675902 441936 675908 441960
rect 675590 441908 675908 441936
rect 675960 441936 675966 441960
rect 676870 441950 677040 441956
rect 675960 441908 676870 441936
rect 676870 441892 677040 441898
rect 675846 441812 675852 441836
rect 675590 441784 675852 441812
rect 675904 441812 675910 441836
rect 677534 441812 677540 441944
rect 675904 441784 677540 441812
rect 677534 441726 677540 441784
rect 677592 441726 677598 441944
rect 675786 441583 675792 441607
rect 675590 441555 675792 441583
rect 675844 441583 675850 441607
rect 676922 441583 676928 441674
rect 675844 441555 676928 441583
rect 676922 441456 676928 441555
rect 676980 441456 676986 441674
rect 675730 441389 675736 441413
rect 675590 441361 675736 441389
rect 675788 441389 675794 441413
rect 677482 441400 677652 441406
rect 675788 441361 677482 441389
rect 677482 441342 677652 441348
rect 675790 440740 675796 440764
rect 675590 440712 675796 440740
rect 675848 440740 675854 440764
rect 676870 440754 677040 440760
rect 675848 440712 676870 440740
rect 676870 440696 677040 440702
rect 675734 440616 675740 440640
rect 675590 440588 675740 440616
rect 675792 440616 675798 440640
rect 677534 440616 677540 440748
rect 675792 440588 677540 440616
rect 677534 440530 677540 440588
rect 677592 440530 677598 440748
rect 675674 440387 675680 440411
rect 675590 440359 675680 440387
rect 675732 440387 675738 440411
rect 676922 440387 676928 440478
rect 675732 440359 676928 440387
rect 676922 440260 676928 440359
rect 676980 440260 676986 440478
rect 675618 440193 675624 440217
rect 675590 440165 675624 440193
rect 675676 440193 675682 440217
rect 677482 440204 677652 440210
rect 675676 440165 677482 440193
rect 677482 440146 677652 440152
rect 675678 439544 675684 439568
rect 675590 439516 675684 439544
rect 675736 439544 675742 439568
rect 676870 439558 677040 439564
rect 675736 439516 676870 439544
rect 676870 439500 677040 439506
rect 675622 439420 675628 439444
rect 675590 439392 675628 439420
rect 675680 439420 675686 439444
rect 677534 439420 677540 439552
rect 675680 439392 677540 439420
rect 677534 439334 677540 439392
rect 677592 439334 677598 439552
rect 40595 346393 40601 346611
rect 40653 346520 40659 346611
rect 41145 346520 41151 346544
rect 40653 346492 41151 346520
rect 41203 346520 41209 346544
rect 41203 346492 42288 346520
rect 40653 346393 40659 346492
rect 39929 346337 40099 346343
rect 41201 346326 41207 346350
rect 40099 346298 41207 346326
rect 41259 346326 41265 346350
rect 41259 346298 42288 346326
rect 39929 346279 40099 346285
rect 40541 345691 40711 345697
rect 39983 345467 39989 345685
rect 40041 345553 40047 345685
rect 41141 345677 41147 345701
rect 40711 345649 41147 345677
rect 41199 345677 41205 345701
rect 41199 345649 42288 345677
rect 40541 345633 40711 345639
rect 41197 345553 41203 345577
rect 40041 345525 41203 345553
rect 41255 345553 41261 345577
rect 41255 345525 42288 345553
rect 40041 345467 40047 345525
rect 40595 345197 40601 345415
rect 40653 345324 40659 345415
rect 41257 345324 41263 345348
rect 40653 345296 41263 345324
rect 41315 345324 41321 345348
rect 41315 345296 42288 345324
rect 40653 345197 40659 345296
rect 39929 345141 40099 345147
rect 41313 345130 41319 345154
rect 40099 345102 41319 345130
rect 41371 345130 41377 345154
rect 41371 345102 42288 345130
rect 39929 345083 40099 345089
rect 40541 344495 40711 344501
rect 39983 344271 39989 344489
rect 40041 344357 40047 344489
rect 41253 344481 41259 344505
rect 40711 344453 41259 344481
rect 41311 344481 41317 344505
rect 41311 344453 42288 344481
rect 40541 344437 40711 344443
rect 41309 344357 41315 344381
rect 40041 344329 41315 344357
rect 41367 344357 41373 344381
rect 41367 344329 42288 344357
rect 40041 344271 40047 344329
rect 40595 344001 40601 344219
rect 40653 344128 40659 344219
rect 41369 344128 41375 344152
rect 40653 344100 41375 344128
rect 41427 344128 41433 344152
rect 41427 344100 42288 344128
rect 40653 344001 40659 344100
rect 39929 343945 40099 343951
rect 41425 343934 41431 343958
rect 40099 343906 41431 343934
rect 41483 343934 41489 343958
rect 41483 343906 42288 343934
rect 39929 343887 40099 343893
rect 40279 343728 40365 343736
rect 40279 343371 40291 343728
rect 40351 343371 40365 343728
rect 40279 343363 40365 343371
rect 40541 343299 40711 343305
rect 39983 343075 39989 343293
rect 40041 343161 40047 343293
rect 41365 343285 41371 343309
rect 40711 343257 41371 343285
rect 41423 343285 41429 343309
rect 41423 343257 42288 343285
rect 40541 343241 40711 343247
rect 41421 343161 41427 343185
rect 40041 343133 41427 343161
rect 41479 343161 41485 343185
rect 41479 343133 42288 343161
rect 40041 343075 40047 343133
rect 40595 342805 40601 343023
rect 40653 342932 40659 343023
rect 41481 342932 41487 342956
rect 40653 342904 41487 342932
rect 41539 342932 41545 342956
rect 41539 342904 42288 342932
rect 40653 342805 40659 342904
rect 39929 342749 40099 342755
rect 41537 342738 41543 342762
rect 40099 342710 41543 342738
rect 41595 342738 41601 342762
rect 41595 342710 42288 342738
rect 39929 342691 40099 342697
rect 39733 342532 39819 342540
rect 39733 342175 39750 342532
rect 39810 342175 39819 342532
rect 39733 342167 39819 342175
rect 40818 342532 40904 342540
rect 40818 342175 40832 342532
rect 40892 342175 40904 342532
rect 40818 342167 40904 342175
rect 40541 342103 40711 342109
rect 39983 341879 39989 342097
rect 40041 341965 40047 342097
rect 41477 342089 41483 342113
rect 40711 342061 41483 342089
rect 41535 342089 41541 342113
rect 41535 342061 42288 342089
rect 40541 342045 40711 342051
rect 41533 341965 41539 341989
rect 40041 341937 41539 341965
rect 41591 341965 41597 341989
rect 41591 341937 42288 341965
rect 40041 341879 40047 341937
rect 40595 341609 40601 341827
rect 40653 341736 40659 341827
rect 41593 341736 41599 341760
rect 40653 341708 41599 341736
rect 41651 341736 41657 341760
rect 41651 341708 42288 341736
rect 40653 341609 40659 341708
rect 39929 341553 40099 341559
rect 41649 341542 41655 341566
rect 40099 341514 41655 341542
rect 41707 341542 41713 341566
rect 41707 341514 42288 341542
rect 39929 341495 40099 341501
rect 40541 340907 40711 340913
rect 39983 340683 39989 340901
rect 40041 340769 40047 340901
rect 41589 340893 41595 340917
rect 40711 340865 41595 340893
rect 41647 340893 41653 340917
rect 41647 340865 42288 340893
rect 40541 340849 40711 340855
rect 41645 340769 41651 340793
rect 40041 340741 41651 340769
rect 41703 340769 41709 340793
rect 41703 340741 42288 340769
rect 40041 340683 40047 340741
rect 40595 340413 40601 340631
rect 40653 340540 40659 340631
rect 41705 340540 41711 340564
rect 40653 340512 41711 340540
rect 41763 340540 41769 340564
rect 41763 340512 42288 340540
rect 40653 340413 40659 340512
rect 39929 340357 40099 340363
rect 41761 340346 41767 340370
rect 40099 340318 41767 340346
rect 41819 340346 41825 340370
rect 41819 340318 42288 340346
rect 39929 340299 40099 340305
rect 40541 339711 40711 339717
rect 39983 339487 39989 339705
rect 40041 339573 40047 339705
rect 41701 339697 41707 339721
rect 40711 339669 41707 339697
rect 41759 339697 41765 339721
rect 41759 339669 42288 339697
rect 40541 339653 40711 339659
rect 41757 339573 41763 339597
rect 40041 339545 41763 339573
rect 41815 339573 41821 339597
rect 41815 339545 42288 339573
rect 40041 339487 40047 339545
rect 40595 339217 40601 339435
rect 40653 339344 40659 339435
rect 41817 339344 41823 339368
rect 40653 339316 41823 339344
rect 41875 339344 41881 339368
rect 41875 339316 42288 339344
rect 40653 339217 40659 339316
rect 39929 339161 40099 339167
rect 41873 339150 41879 339174
rect 40099 339122 41879 339150
rect 41931 339150 41937 339174
rect 41931 339122 42288 339150
rect 39929 339103 40099 339109
rect 40541 338515 40711 338521
rect 39983 338291 39989 338509
rect 40041 338377 40047 338509
rect 41813 338501 41819 338525
rect 40711 338473 41819 338501
rect 41871 338501 41877 338525
rect 41871 338473 42288 338501
rect 40541 338457 40711 338463
rect 41869 338377 41875 338401
rect 40041 338349 41875 338377
rect 41927 338377 41933 338401
rect 41927 338349 42288 338377
rect 40041 338291 40047 338349
rect 40595 338021 40601 338239
rect 40653 338148 40659 338239
rect 41929 338148 41935 338172
rect 40653 338120 41935 338148
rect 41987 338148 41993 338172
rect 41987 338120 42288 338148
rect 40653 338021 40659 338120
rect 39929 337965 40099 337971
rect 41985 337954 41991 337978
rect 40099 337926 41991 337954
rect 42043 337954 42049 337978
rect 42043 337926 42288 337954
rect 39929 337907 40099 337913
rect 40541 337319 40711 337325
rect 39983 337095 39989 337313
rect 40041 337181 40047 337313
rect 41925 337305 41931 337329
rect 40711 337277 41931 337305
rect 41983 337305 41989 337329
rect 41983 337277 42288 337305
rect 40541 337261 40711 337267
rect 41981 337181 41987 337205
rect 40041 337153 41987 337181
rect 42039 337181 42045 337205
rect 42039 337153 42288 337181
rect 40041 337095 40047 337153
rect 40595 336825 40601 337043
rect 40653 336952 40659 337043
rect 40653 336924 42047 336952
rect 40653 336825 40659 336924
rect 42041 336900 42047 336924
rect 42099 336924 42288 336952
rect 42099 336900 42105 336924
rect 39929 336769 40099 336775
rect 42097 336758 42103 336782
rect 40099 336730 42103 336758
rect 42155 336758 42161 336782
rect 42155 336730 42288 336758
rect 39929 336711 40099 336717
rect 40541 336123 40711 336129
rect 39983 335899 39989 336117
rect 40041 335985 40047 336117
rect 42037 336109 42043 336133
rect 40711 336081 42043 336109
rect 42095 336109 42101 336133
rect 42095 336081 42288 336109
rect 40541 336065 40711 336071
rect 42093 335985 42099 336009
rect 40041 335957 42099 335985
rect 42151 335985 42157 336009
rect 42151 335957 42288 335985
rect 40041 335899 40047 335957
rect 40595 335629 40601 335847
rect 40653 335756 40659 335847
rect 42153 335756 42159 335780
rect 40653 335728 42159 335756
rect 42211 335756 42217 335780
rect 42211 335728 42288 335756
rect 40653 335629 40659 335728
rect 39929 335573 40099 335579
rect 42209 335562 42215 335586
rect 40099 335534 42215 335562
rect 42267 335562 42273 335586
rect 42267 335534 42288 335562
rect 39929 335515 40099 335521
rect 40541 334927 40711 334933
rect 39983 334703 39989 334921
rect 40041 334789 40047 334921
rect 42149 334913 42155 334937
rect 40711 334885 42155 334913
rect 42207 334913 42213 334937
rect 42207 334885 42288 334913
rect 40541 334869 40711 334875
rect 42205 334789 42211 334813
rect 40041 334761 42211 334789
rect 42263 334789 42269 334813
rect 42263 334761 42288 334789
rect 40041 334703 40047 334761
rect 394104 225374 394132 225393
rect 394947 225378 394975 225393
rect 394104 225368 394156 225374
rect 134104 225346 134132 225365
rect 134947 225350 134975 225365
rect 134104 225340 134156 225346
rect 134104 225282 134156 225288
rect 134947 225344 134999 225350
rect 134947 225286 134999 225292
rect 135176 225290 135204 225365
rect 134104 223272 134132 225282
rect 134088 223102 134094 223272
rect 134146 223102 134152 223272
rect 134947 223220 134975 225286
rect 135176 225284 135228 225290
rect 135176 225226 135228 225232
rect 135300 225234 135328 225365
rect 135949 225294 135977 225365
rect 135949 225288 136001 225294
rect 135300 225228 135352 225234
rect 134848 223214 135066 223220
rect 134848 223156 135066 223162
rect 135176 222608 135204 225226
rect 135300 225170 135352 225176
rect 135949 225230 136001 225236
rect 136143 225238 136171 225365
rect 136143 225232 136195 225238
rect 135300 223272 135328 225170
rect 135284 223102 135290 223272
rect 135342 223102 135348 223272
rect 135949 222660 135977 225230
rect 136143 225174 136195 225180
rect 136372 225178 136400 225365
rect 136143 223220 136171 225174
rect 136372 225172 136424 225178
rect 136372 225114 136424 225120
rect 136496 225122 136524 225365
rect 137145 225182 137173 225365
rect 137145 225176 137197 225182
rect 136496 225116 136548 225122
rect 136044 223214 136262 223220
rect 136044 223156 136262 223162
rect 135118 222602 135336 222608
rect 135118 222544 135336 222550
rect 135930 222490 135936 222660
rect 135988 222490 135994 222660
rect 136372 222608 136400 225114
rect 136496 225058 136548 225064
rect 137145 225118 137197 225124
rect 137339 225126 137367 225365
rect 137339 225120 137391 225126
rect 136496 223272 136524 225058
rect 136480 223102 136486 223272
rect 136538 223102 136544 223272
rect 137145 222660 137173 225118
rect 137339 225062 137391 225068
rect 137568 225066 137596 225365
rect 137339 223220 137367 225062
rect 137568 225060 137620 225066
rect 137568 225002 137620 225008
rect 137692 225010 137720 225365
rect 138341 225070 138369 225365
rect 138341 225064 138393 225070
rect 137692 225004 137744 225010
rect 137240 223214 137458 223220
rect 137240 223156 137458 223162
rect 136314 222602 136532 222608
rect 136314 222544 136532 222550
rect 137126 222490 137132 222660
rect 137184 222490 137190 222660
rect 137568 222608 137596 225002
rect 137692 224946 137744 224952
rect 138341 225006 138393 225012
rect 138535 225014 138563 225365
rect 138535 225008 138587 225014
rect 137692 223272 137720 224946
rect 137676 223102 137682 223272
rect 137734 223102 137740 223272
rect 138341 222660 138369 225006
rect 138535 224950 138587 224956
rect 138764 224954 138792 225365
rect 138535 223220 138563 224950
rect 138764 224948 138816 224954
rect 138764 224890 138816 224896
rect 138888 224898 138916 225365
rect 139537 224958 139565 225365
rect 139537 224952 139589 224958
rect 138888 224892 138940 224898
rect 138436 223214 138654 223220
rect 138436 223156 138654 223162
rect 137510 222602 137728 222608
rect 137510 222544 137728 222550
rect 138322 222490 138328 222660
rect 138380 222490 138386 222660
rect 138764 222608 138792 224890
rect 138888 224834 138940 224840
rect 139537 224894 139589 224900
rect 139731 224902 139759 225365
rect 139731 224896 139783 224902
rect 138888 223272 138916 224834
rect 138872 223102 138878 223272
rect 138930 223102 138936 223272
rect 139537 222660 139565 224894
rect 139731 224838 139783 224844
rect 139960 224842 139988 225365
rect 139731 223220 139759 224838
rect 139960 224836 140012 224842
rect 139960 224778 140012 224784
rect 140084 224786 140112 225365
rect 140733 224846 140761 225365
rect 140733 224840 140785 224846
rect 140927 224790 140955 225365
rect 140084 224780 140136 224786
rect 139632 223214 139850 223220
rect 139632 223156 139850 223162
rect 138706 222602 138924 222608
rect 138706 222544 138924 222550
rect 139518 222490 139524 222660
rect 139576 222490 139582 222660
rect 139960 222608 139988 224778
rect 140084 224722 140136 224728
rect 140733 224782 140785 224788
rect 140903 224784 140955 224790
rect 140084 223272 140112 224722
rect 140068 223102 140074 223272
rect 140126 223102 140132 223272
rect 140733 222660 140761 224782
rect 140903 224726 140955 224732
rect 140927 223220 140955 224726
rect 141156 224730 141184 225365
rect 141156 224724 141208 224730
rect 141156 224666 141208 224672
rect 141280 224674 141308 225365
rect 141929 224734 141957 225365
rect 141929 224728 141981 224734
rect 141280 224668 141332 224674
rect 140828 223214 141046 223220
rect 140828 223156 141046 223162
rect 139902 222602 140120 222608
rect 139902 222544 140120 222550
rect 140714 222490 140720 222660
rect 140772 222490 140778 222660
rect 141156 222608 141184 224666
rect 141280 224610 141332 224616
rect 141929 224670 141981 224676
rect 142123 224678 142151 225365
rect 142123 224672 142175 224678
rect 141280 223272 141308 224610
rect 141264 223102 141270 223272
rect 141322 223102 141328 223272
rect 141929 222660 141957 224670
rect 142123 224614 142175 224620
rect 142352 224618 142380 225365
rect 142123 223220 142151 224614
rect 142352 224612 142404 224618
rect 142352 224554 142404 224560
rect 142476 224562 142504 225365
rect 143125 224622 143153 225365
rect 143125 224616 143177 224622
rect 143319 224566 143347 225365
rect 142476 224556 142528 224562
rect 142024 223214 142242 223220
rect 142024 223156 142242 223162
rect 141098 222602 141316 222608
rect 141098 222544 141316 222550
rect 141910 222490 141916 222660
rect 141968 222490 141974 222660
rect 142352 222608 142380 224554
rect 142476 224498 142528 224504
rect 143125 224558 143177 224564
rect 143295 224560 143347 224566
rect 142476 223272 142504 224498
rect 142460 223102 142466 223272
rect 142518 223102 142524 223272
rect 143125 222660 143153 224558
rect 143295 224502 143347 224508
rect 143319 223220 143347 224502
rect 143548 224506 143576 225365
rect 143548 224500 143600 224506
rect 143548 224442 143600 224448
rect 143672 224450 143700 225365
rect 144321 224510 144349 225365
rect 144321 224504 144373 224510
rect 143672 224444 143724 224450
rect 143220 223214 143438 223220
rect 143220 223156 143438 223162
rect 142294 222602 142512 222608
rect 142294 222544 142512 222550
rect 143106 222490 143112 222660
rect 143164 222490 143170 222660
rect 143548 222608 143576 224442
rect 143672 224386 143724 224392
rect 144321 224446 144373 224452
rect 144515 224454 144543 225365
rect 144515 224448 144567 224454
rect 143672 223272 143700 224386
rect 143656 223102 143662 223272
rect 143714 223102 143720 223272
rect 144321 222660 144349 224446
rect 144515 224390 144567 224396
rect 144744 224394 144772 225365
rect 144515 223220 144543 224390
rect 144744 224388 144796 224394
rect 144744 224330 144796 224336
rect 144868 224338 144896 225365
rect 145517 224398 145545 225365
rect 145517 224392 145569 224398
rect 144868 224332 144920 224338
rect 144416 223214 144634 223220
rect 144416 223156 144634 223162
rect 143490 222602 143708 222608
rect 143490 222544 143708 222550
rect 144302 222490 144308 222660
rect 144360 222490 144366 222660
rect 144744 222608 144772 224330
rect 144868 224274 144920 224280
rect 145517 224334 145569 224340
rect 145711 224342 145739 225365
rect 145711 224336 145763 224342
rect 144868 223272 144896 224274
rect 144852 223102 144858 223272
rect 144910 223102 144916 223272
rect 145517 222660 145545 224334
rect 145711 224278 145763 224284
rect 145940 224282 145968 225365
rect 146713 224286 146741 225365
rect 145711 223220 145739 224278
rect 145940 224276 145992 224282
rect 145940 224218 145992 224224
rect 146713 224280 146765 224286
rect 146713 224222 146765 224228
rect 147260 224226 147288 225365
rect 148103 224230 148131 225365
rect 145612 223214 145830 223220
rect 145612 223156 145830 223162
rect 144686 222602 144904 222608
rect 144686 222544 144904 222550
rect 145498 222490 145504 222660
rect 145556 222490 145562 222660
rect 145940 222608 145968 224218
rect 146191 222916 146564 222930
rect 146191 222856 146199 222916
rect 146556 222856 146564 222916
rect 146191 222844 146564 222856
rect 146713 222660 146741 224222
rect 147260 224220 147312 224226
rect 147260 224162 147312 224168
rect 148103 224224 148155 224230
rect 148103 224166 148155 224172
rect 148332 224170 148360 225365
rect 147260 223272 147288 224162
rect 147244 223102 147250 223272
rect 147302 223102 147308 223272
rect 148103 223220 148131 224166
rect 148332 224164 148384 224170
rect 148332 224106 148384 224112
rect 148456 224114 148484 225365
rect 149105 224174 149133 225365
rect 149105 224168 149157 224174
rect 148456 224108 148508 224114
rect 148004 223214 148222 223220
rect 148004 223156 148222 223162
rect 145882 222602 146100 222608
rect 145882 222544 146100 222550
rect 146694 222490 146700 222660
rect 146752 222490 146758 222660
rect 148332 222608 148360 224106
rect 148456 224050 148508 224056
rect 149105 224110 149157 224116
rect 149299 224118 149327 225365
rect 149299 224112 149351 224118
rect 148456 223272 148484 224050
rect 148440 223102 148446 223272
rect 148498 223102 148504 223272
rect 149105 222660 149133 224110
rect 149299 224054 149351 224060
rect 149528 224058 149556 225365
rect 149299 223220 149327 224054
rect 149528 224052 149580 224058
rect 149528 223994 149580 224000
rect 149652 224002 149680 225365
rect 150301 224062 150329 225365
rect 150301 224056 150353 224062
rect 150495 224006 150523 225365
rect 149652 223996 149704 224002
rect 149200 223214 149418 223220
rect 149200 223156 149418 223162
rect 148274 222602 148492 222608
rect 148274 222544 148492 222550
rect 149086 222490 149092 222660
rect 149144 222490 149150 222660
rect 149528 222608 149556 223994
rect 149652 223938 149704 223944
rect 150301 223998 150353 224004
rect 150471 224000 150523 224006
rect 149652 223272 149680 223938
rect 149636 223102 149642 223272
rect 149694 223102 149700 223272
rect 150301 222660 150329 223998
rect 150471 223942 150523 223948
rect 150495 223220 150523 223942
rect 150724 223946 150752 225365
rect 150724 223940 150776 223946
rect 150724 223882 150776 223888
rect 150848 223890 150876 225365
rect 151497 223950 151525 225365
rect 151497 223944 151549 223950
rect 150848 223884 150900 223890
rect 150396 223214 150614 223220
rect 150396 223156 150614 223162
rect 149470 222602 149688 222608
rect 149470 222544 149688 222550
rect 150282 222490 150288 222660
rect 150340 222490 150346 222660
rect 150724 222608 150752 223882
rect 150848 223826 150900 223832
rect 151497 223886 151549 223892
rect 151691 223894 151719 225365
rect 151691 223888 151743 223894
rect 150848 223272 150876 223826
rect 150832 223102 150838 223272
rect 150890 223102 150896 223272
rect 151497 222660 151525 223886
rect 151691 223830 151743 223836
rect 151920 223834 151948 225365
rect 151691 223220 151719 223830
rect 151920 223828 151972 223834
rect 151920 223770 151972 223776
rect 152044 223778 152072 225365
rect 152693 223838 152721 225365
rect 152693 223832 152745 223838
rect 152887 223782 152915 225365
rect 152044 223772 152096 223778
rect 151592 223214 151810 223220
rect 151592 223156 151810 223162
rect 150666 222602 150884 222608
rect 150666 222544 150884 222550
rect 151478 222490 151484 222660
rect 151536 222490 151542 222660
rect 151920 222608 151948 223770
rect 152044 223714 152096 223720
rect 152693 223774 152745 223780
rect 152863 223776 152915 223782
rect 152044 223272 152072 223714
rect 152028 223102 152034 223272
rect 152086 223102 152092 223272
rect 152693 222660 152721 223774
rect 152863 223718 152915 223724
rect 152887 223220 152915 223718
rect 153116 223722 153144 225365
rect 153116 223716 153168 223722
rect 153116 223658 153168 223664
rect 153240 223666 153268 225365
rect 153889 223726 153917 225365
rect 153889 223720 153941 223726
rect 153240 223660 153292 223666
rect 152788 223214 153006 223220
rect 152788 223156 153006 223162
rect 153116 222848 153144 223658
rect 153240 223602 153292 223608
rect 153889 223662 153941 223668
rect 154083 223670 154111 225365
rect 394104 225310 394156 225316
rect 394947 225372 394999 225378
rect 394947 225314 394999 225320
rect 395176 225318 395204 225393
rect 154083 223664 154135 223670
rect 153240 223272 153268 223602
rect 153224 223102 153230 223272
rect 153282 223102 153288 223272
rect 153889 222848 153917 223662
rect 154083 223606 154135 223612
rect 154083 223220 154111 223606
rect 394104 223272 394132 225310
rect 153984 223214 154202 223220
rect 153984 223156 154202 223162
rect 394088 223102 394094 223272
rect 394146 223102 394152 223272
rect 394947 223220 394975 225314
rect 395176 225312 395228 225318
rect 395176 225254 395228 225260
rect 395300 225262 395328 225393
rect 395949 225322 395977 225393
rect 395949 225316 396001 225322
rect 395300 225256 395352 225262
rect 394848 223214 395066 223220
rect 394848 223156 395066 223162
rect 153116 222820 153271 222848
rect 153889 222820 154044 222848
rect 153243 222660 153271 222820
rect 151862 222602 152080 222608
rect 151862 222544 152080 222550
rect 152674 222490 152680 222660
rect 152732 222490 152738 222660
rect 153226 222490 153232 222660
rect 153284 222490 153290 222660
rect 154016 222608 154044 222820
rect 395176 222608 395204 225254
rect 395300 225198 395352 225204
rect 395949 225258 396001 225264
rect 396143 225266 396171 225393
rect 396143 225260 396195 225266
rect 395300 223272 395328 225198
rect 395284 223102 395290 223272
rect 395342 223102 395348 223272
rect 395949 222660 395977 225258
rect 396143 225202 396195 225208
rect 396372 225206 396400 225393
rect 396143 223220 396171 225202
rect 396372 225200 396424 225206
rect 396372 225142 396424 225148
rect 396496 225150 396524 225393
rect 397145 225210 397173 225393
rect 397145 225204 397197 225210
rect 396496 225144 396548 225150
rect 396044 223214 396262 223220
rect 396044 223156 396262 223162
rect 153884 222602 154102 222608
rect 153884 222544 154102 222550
rect 395118 222602 395336 222608
rect 395118 222544 395336 222550
rect 395930 222490 395936 222660
rect 395988 222490 395994 222660
rect 396372 222608 396400 225142
rect 396496 225086 396548 225092
rect 397145 225146 397197 225152
rect 397339 225154 397367 225393
rect 397339 225148 397391 225154
rect 396496 223272 396524 225086
rect 396480 223102 396486 223272
rect 396538 223102 396544 223272
rect 397145 222660 397173 225146
rect 397339 225090 397391 225096
rect 397568 225094 397596 225393
rect 397339 223220 397367 225090
rect 397568 225088 397620 225094
rect 397568 225030 397620 225036
rect 397692 225038 397720 225393
rect 398341 225098 398369 225393
rect 398341 225092 398393 225098
rect 397692 225032 397744 225038
rect 397240 223214 397458 223220
rect 397240 223156 397458 223162
rect 396314 222602 396532 222608
rect 396314 222544 396532 222550
rect 397126 222490 397132 222660
rect 397184 222490 397190 222660
rect 397568 222608 397596 225030
rect 397692 224974 397744 224980
rect 398341 225034 398393 225040
rect 398535 225042 398563 225393
rect 398535 225036 398587 225042
rect 397692 223272 397720 224974
rect 397676 223102 397682 223272
rect 397734 223102 397740 223272
rect 398341 222660 398369 225034
rect 398535 224978 398587 224984
rect 398764 224982 398792 225393
rect 398535 223220 398563 224978
rect 398764 224976 398816 224982
rect 398764 224918 398816 224924
rect 398888 224926 398916 225393
rect 399537 224986 399565 225393
rect 399537 224980 399589 224986
rect 398888 224920 398940 224926
rect 398436 223214 398654 223220
rect 398436 223156 398654 223162
rect 397510 222602 397728 222608
rect 397510 222544 397728 222550
rect 398322 222490 398328 222660
rect 398380 222490 398386 222660
rect 398764 222608 398792 224918
rect 398888 224862 398940 224868
rect 399537 224922 399589 224928
rect 399731 224930 399759 225393
rect 399731 224924 399783 224930
rect 398888 223272 398916 224862
rect 398872 223102 398878 223272
rect 398930 223102 398936 223272
rect 399537 222660 399565 224922
rect 399731 224866 399783 224872
rect 399960 224870 399988 225393
rect 399731 223220 399759 224866
rect 399960 224864 400012 224870
rect 399960 224806 400012 224812
rect 400084 224814 400112 225393
rect 400733 224874 400761 225393
rect 400733 224868 400785 224874
rect 400927 224818 400955 225393
rect 400084 224808 400136 224814
rect 399632 223214 399850 223220
rect 399632 223156 399850 223162
rect 398706 222602 398924 222608
rect 398706 222544 398924 222550
rect 399518 222490 399524 222660
rect 399576 222490 399582 222660
rect 399960 222608 399988 224806
rect 400084 224750 400136 224756
rect 400733 224810 400785 224816
rect 400903 224812 400955 224818
rect 400084 223272 400112 224750
rect 400068 223102 400074 223272
rect 400126 223102 400132 223272
rect 400733 222660 400761 224810
rect 400903 224754 400955 224760
rect 400927 223220 400955 224754
rect 401156 224758 401184 225393
rect 401156 224752 401208 224758
rect 401156 224694 401208 224700
rect 401280 224702 401308 225393
rect 401929 224762 401957 225393
rect 401929 224756 401981 224762
rect 401280 224696 401332 224702
rect 400828 223214 401046 223220
rect 400828 223156 401046 223162
rect 399902 222602 400120 222608
rect 399902 222544 400120 222550
rect 400714 222490 400720 222660
rect 400772 222490 400778 222660
rect 401156 222608 401184 224694
rect 401280 224638 401332 224644
rect 401929 224698 401981 224704
rect 402123 224706 402151 225393
rect 402123 224700 402175 224706
rect 401280 223272 401308 224638
rect 401264 223102 401270 223272
rect 401322 223102 401328 223272
rect 401929 222660 401957 224698
rect 402123 224642 402175 224648
rect 402352 224646 402380 225393
rect 402123 223220 402151 224642
rect 402352 224640 402404 224646
rect 402352 224582 402404 224588
rect 402476 224590 402504 225393
rect 403125 224650 403153 225393
rect 403125 224644 403177 224650
rect 403319 224594 403347 225393
rect 402476 224584 402528 224590
rect 402024 223214 402242 223220
rect 402024 223156 402242 223162
rect 401098 222602 401316 222608
rect 401098 222544 401316 222550
rect 401910 222490 401916 222660
rect 401968 222490 401974 222660
rect 402352 222608 402380 224582
rect 402476 224526 402528 224532
rect 403125 224586 403177 224592
rect 403295 224588 403347 224594
rect 402476 223272 402504 224526
rect 402460 223102 402466 223272
rect 402518 223102 402524 223272
rect 403125 222660 403153 224586
rect 403295 224530 403347 224536
rect 403319 223220 403347 224530
rect 403548 224534 403576 225393
rect 403548 224528 403600 224534
rect 403548 224470 403600 224476
rect 403672 224478 403700 225393
rect 404321 224538 404349 225393
rect 404321 224532 404373 224538
rect 403672 224472 403724 224478
rect 403220 223214 403438 223220
rect 403220 223156 403438 223162
rect 402294 222602 402512 222608
rect 402294 222544 402512 222550
rect 403106 222490 403112 222660
rect 403164 222490 403170 222660
rect 403548 222608 403576 224470
rect 403672 224414 403724 224420
rect 404321 224474 404373 224480
rect 404515 224482 404543 225393
rect 404515 224476 404567 224482
rect 403672 223272 403700 224414
rect 403656 223102 403662 223272
rect 403714 223102 403720 223272
rect 404321 222660 404349 224474
rect 404515 224418 404567 224424
rect 404744 224422 404772 225393
rect 404515 223220 404543 224418
rect 404744 224416 404796 224422
rect 404744 224358 404796 224364
rect 404868 224366 404896 225393
rect 405517 224426 405545 225393
rect 405517 224420 405569 224426
rect 404868 224360 404920 224366
rect 404416 223214 404634 223220
rect 404416 223156 404634 223162
rect 403490 222602 403708 222608
rect 403490 222544 403708 222550
rect 404302 222490 404308 222660
rect 404360 222490 404366 222660
rect 404744 222608 404772 224358
rect 404868 224302 404920 224308
rect 405517 224362 405569 224368
rect 405711 224370 405739 225393
rect 405711 224364 405763 224370
rect 404868 223272 404896 224302
rect 404852 223102 404858 223272
rect 404910 223102 404916 223272
rect 405022 222909 405395 222923
rect 405022 222849 405030 222909
rect 405387 222849 405395 222909
rect 405022 222837 405395 222849
rect 405517 222660 405545 224362
rect 405711 224306 405763 224312
rect 405940 224310 405968 225393
rect 406713 224314 406741 225393
rect 405711 223220 405739 224306
rect 405940 224304 405992 224310
rect 405940 224246 405992 224252
rect 406713 224308 406765 224314
rect 406713 224250 406765 224256
rect 407260 224254 407288 225393
rect 408103 224258 408131 225393
rect 405612 223214 405830 223220
rect 405612 223156 405830 223162
rect 404686 222602 404904 222608
rect 404686 222544 404904 222550
rect 405498 222490 405504 222660
rect 405556 222490 405562 222660
rect 405940 222608 405968 224246
rect 406218 223450 406591 223462
rect 406218 223390 406226 223450
rect 406583 223390 406591 223450
rect 406218 223376 406591 223390
rect 406713 222660 406741 224250
rect 407260 224248 407312 224254
rect 407260 224190 407312 224196
rect 408103 224252 408155 224258
rect 408103 224194 408155 224200
rect 408332 224198 408360 225393
rect 407260 223272 407288 224190
rect 407244 223102 407250 223272
rect 407302 223102 407308 223272
rect 408103 223220 408131 224194
rect 408332 224192 408384 224198
rect 408332 224134 408384 224140
rect 408456 224142 408484 225393
rect 409105 224202 409133 225393
rect 409105 224196 409157 224202
rect 408456 224136 408508 224142
rect 408004 223214 408222 223220
rect 408004 223156 408222 223162
rect 405882 222602 406100 222608
rect 405882 222544 406100 222550
rect 406694 222490 406700 222660
rect 406752 222490 406758 222660
rect 408332 222608 408360 224134
rect 408456 224078 408508 224084
rect 409105 224138 409157 224144
rect 409299 224146 409327 225393
rect 409299 224140 409351 224146
rect 408456 223272 408484 224078
rect 408440 223102 408446 223272
rect 408498 223102 408504 223272
rect 409105 222660 409133 224138
rect 409299 224082 409351 224088
rect 409528 224086 409556 225393
rect 409299 223220 409327 224082
rect 409528 224080 409580 224086
rect 409528 224022 409580 224028
rect 409652 224030 409680 225393
rect 410301 224090 410329 225393
rect 410301 224084 410353 224090
rect 410495 224034 410523 225393
rect 409652 224024 409704 224030
rect 409200 223214 409418 223220
rect 409200 223156 409418 223162
rect 408274 222602 408492 222608
rect 408274 222544 408492 222550
rect 409086 222490 409092 222660
rect 409144 222490 409150 222660
rect 409528 222608 409556 224022
rect 409652 223966 409704 223972
rect 410301 224026 410353 224032
rect 410471 224028 410523 224034
rect 409652 223272 409680 223966
rect 409636 223102 409642 223272
rect 409694 223102 409700 223272
rect 410301 222660 410329 224026
rect 410471 223970 410523 223976
rect 410495 223220 410523 223970
rect 410724 223974 410752 225393
rect 410724 223968 410776 223974
rect 410724 223910 410776 223916
rect 410848 223918 410876 225393
rect 411497 223978 411525 225393
rect 411497 223972 411549 223978
rect 410848 223912 410900 223918
rect 410396 223214 410614 223220
rect 410396 223156 410614 223162
rect 409470 222602 409688 222608
rect 409470 222544 409688 222550
rect 410282 222490 410288 222660
rect 410340 222490 410346 222660
rect 410724 222608 410752 223910
rect 410848 223854 410900 223860
rect 411497 223914 411549 223920
rect 411691 223922 411719 225393
rect 411691 223916 411743 223922
rect 410848 223272 410876 223854
rect 410832 223102 410838 223272
rect 410890 223102 410896 223272
rect 411497 222660 411525 223914
rect 411691 223858 411743 223864
rect 411920 223862 411948 225393
rect 411691 223220 411719 223858
rect 411920 223856 411972 223862
rect 411920 223798 411972 223804
rect 412044 223806 412072 225393
rect 412693 223866 412721 225393
rect 412693 223860 412745 223866
rect 412887 223810 412915 225393
rect 412044 223800 412096 223806
rect 411592 223214 411810 223220
rect 411592 223156 411810 223162
rect 410666 222602 410884 222608
rect 410666 222544 410884 222550
rect 411478 222490 411484 222660
rect 411536 222490 411542 222660
rect 411920 222608 411948 223798
rect 412044 223742 412096 223748
rect 412693 223802 412745 223808
rect 412863 223804 412915 223810
rect 412044 223272 412072 223742
rect 412028 223102 412034 223272
rect 412086 223102 412092 223272
rect 412693 222660 412721 223802
rect 412863 223746 412915 223752
rect 412887 223220 412915 223746
rect 413116 223750 413144 225393
rect 413116 223744 413168 223750
rect 413116 223686 413168 223692
rect 413240 223694 413268 225393
rect 413889 223754 413917 225393
rect 413889 223748 413941 223754
rect 413240 223688 413292 223694
rect 412788 223214 413006 223220
rect 412788 223156 413006 223162
rect 413116 222834 413144 223686
rect 413240 223630 413292 223636
rect 413889 223690 413941 223696
rect 414083 223698 414111 225393
rect 414083 223692 414135 223698
rect 413240 223272 413268 223630
rect 413224 223102 413230 223272
rect 413282 223102 413288 223272
rect 413889 222834 413917 223690
rect 414083 223634 414135 223640
rect 414083 223220 414111 223634
rect 413984 223214 414202 223220
rect 413984 223156 414202 223162
rect 413116 222806 413271 222834
rect 413889 222806 414044 222834
rect 413243 222660 413271 222806
rect 411862 222602 412080 222608
rect 411862 222544 412080 222550
rect 412674 222490 412680 222660
rect 412732 222490 412738 222660
rect 413226 222490 413232 222660
rect 413284 222490 413290 222660
rect 414016 222608 414044 222806
rect 413884 222602 414102 222608
rect 413884 222544 414102 222550
rect 147387 222375 147760 222384
rect 147387 222315 147395 222375
rect 147752 222315 147760 222375
rect 147387 222298 147760 222315
rect 406218 222368 406591 222377
rect 406218 222308 406226 222368
rect 406583 222308 406591 222368
rect 406218 222291 406591 222308
<< via2 >>
rect 676693 707708 676753 708065
rect 677775 707708 677835 708065
rect 677234 706512 677294 706869
rect 39731 604014 39791 604371
rect 40813 604014 40873 604371
rect 40272 602818 40332 603175
rect 677226 446899 677286 447256
rect 676685 445703 676745 446060
rect 677767 445703 677827 446060
rect 40291 343371 40351 343728
rect 39750 342175 39810 342532
rect 40832 342175 40892 342532
rect 146199 222856 146556 222916
rect 147395 223397 147752 223457
rect 405030 222849 405387 222909
rect 406226 223390 406583 223450
rect 147395 222315 147752 222375
rect 406226 222308 406583 222368
<< metal3 >>
rect 676678 708065 678183 708074
rect 676678 707708 676693 708065
rect 676753 707708 677775 708065
rect 677835 707708 678183 708065
rect 676678 707701 678183 707708
rect 677220 706869 678183 706876
rect 677220 706512 677234 706869
rect 677294 706512 678183 706869
rect 677220 706506 678183 706512
rect 39383 604371 40888 604378
rect 39383 604014 39731 604371
rect 39791 604014 40813 604371
rect 40873 604014 40888 604371
rect 39383 604005 40888 604014
rect 39383 603175 40346 603181
rect 39383 602818 40272 603175
rect 40332 602818 40346 603175
rect 39383 602811 40346 602818
rect 677212 447256 678175 447263
rect 677212 446899 677226 447256
rect 677286 446899 678175 447256
rect 677212 446893 678175 446899
rect 676670 446060 678175 446069
rect 676670 445703 676685 446060
rect 676745 445703 677767 446060
rect 677827 445703 678175 446060
rect 676670 445696 678175 445703
rect 39402 343728 40365 343734
rect 39402 343371 40291 343728
rect 40351 343371 40365 343728
rect 39402 343364 40365 343371
rect 39402 342532 40907 342539
rect 39402 342175 39750 342532
rect 39810 342175 40832 342532
rect 40892 342175 40907 342532
rect 39402 342166 40907 342175
rect 147388 223457 147761 223472
rect 147388 223397 147395 223457
rect 147752 223397 147761 223457
rect 146193 222916 146563 222930
rect 146193 222856 146199 222916
rect 146556 222856 146563 222916
rect 146193 221967 146563 222856
rect 147388 222375 147761 223397
rect 406219 223450 406592 223465
rect 406219 223390 406226 223450
rect 406583 223390 406592 223450
rect 147388 222315 147395 222375
rect 147752 222315 147761 222375
rect 147388 221967 147761 222315
rect 405024 222909 405394 222923
rect 405024 222849 405030 222909
rect 405387 222849 405394 222909
rect 405024 221960 405394 222849
rect 406219 222368 406592 223390
rect 406219 222308 406226 222368
rect 406583 222308 406592 222368
rect 406219 221960 406592 222308
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 134996 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_2
timestamp 1663859327
transform 1 0 148244 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_3
timestamp 1663859327
transform -1 0 149348 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_4
timestamp 1663859327
transform 1 0 150636 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_5
timestamp 1663859327
transform -1 0 151740 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_6
timestamp 1663859327
transform 1 0 151832 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_7
timestamp 1663859327
transform -1 0 152936 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_8
timestamp 1663859327
transform -1 0 154132 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_9
timestamp 1663859327
transform -1 0 154132 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_12
timestamp 1663859327
transform 0 -1 677805 1 0 439304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_13
timestamp 1663859327
transform 0 1 676717 -1 0 440408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_24
timestamp 1663859327
transform 0 -1 677805 1 0 707304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_25
timestamp 1663859327
transform 0 1 676717 -1 0 708408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_34
timestamp 1663859327
transform 0 1 676717 -1 0 446388
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_35
timestamp 1663859327
transform 0 -1 677805 1 0 445284
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_36
timestamp 1663859327
transform 0 1 676717 -1 0 447584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_37
timestamp 1663859327
transform 0 -1 677805 1 0 446480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_46
timestamp 1663859327
transform 0 1 676717 -1 0 441604
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_47
timestamp 1663859327
transform 0 -1 677805 1 0 440500
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_48
timestamp 1663859327
transform 0 -1 677805 1 0 441696
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_49
timestamp 1663859327
transform 0 1 676717 -1 0 442800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_50
timestamp 1663859327
transform 0 -1 677805 1 0 442892
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_51
timestamp 1663859327
transform 0 1 676717 -1 0 443996
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_52
timestamp 1663859327
transform 0 -1 677805 1 0 444088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_53
timestamp 1663859327
transform 0 1 676717 -1 0 445192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_54
timestamp 1663859327
transform 1 0 147048 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_55
timestamp 1663859327
transform -1 0 148152 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_64
timestamp 1663859327
transform 1 0 145852 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_65
timestamp 1663859327
transform -1 0 146956 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_66
timestamp 1663859327
transform -1 0 145760 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_67
timestamp 1663859327
transform 1 0 144656 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_68
timestamp 1663859327
transform 1 0 143460 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_69
timestamp 1663859327
transform -1 0 144564 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_70
timestamp 1663859327
transform 1 0 142264 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_71
timestamp 1663859327
transform -1 0 143368 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_72
timestamp 1663859327
transform 1 0 141068 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_73
timestamp 1663859327
transform -1 0 142172 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_74
timestamp 1663859327
transform 1 0 139872 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_75
timestamp 1663859327
transform -1 0 140976 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_76
timestamp 1663859327
transform 1 0 138676 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_77
timestamp 1663859327
transform -1 0 139780 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_78
timestamp 1663859327
transform -1 0 138584 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_79
timestamp 1663859327
transform 1 0 137480 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_80
timestamp 1663859327
transform 1 0 136284 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_81
timestamp 1663859327
transform -1 0 137388 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_82
timestamp 1663859327
transform 1 0 135088 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_83
timestamp 1663859327
transform -1 0 136192 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_84
timestamp 1663859327
transform -1 0 150544 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_85
timestamp 1663859327
transform 1 0 149440 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_86
timestamp 1663859327
transform -1 0 394996 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_88
timestamp 1663859327
transform -1 0 396192 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_89
timestamp 1663859327
transform 1 0 395088 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_90
timestamp 1663859327
transform 1 0 396284 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_91
timestamp 1663859327
transform -1 0 397388 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_92
timestamp 1663859327
transform -1 0 398584 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_93
timestamp 1663859327
transform 1 0 397480 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_94
timestamp 1663859327
transform -1 0 399780 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_95
timestamp 1663859327
transform 1 0 398676 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_96
timestamp 1663859327
transform 1 0 399872 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_97
timestamp 1663859327
transform 1 0 401068 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_98
timestamp 1663859327
transform -1 0 400976 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_99
timestamp 1663859327
transform -1 0 402172 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_100
timestamp 1663859327
transform 1 0 402264 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_101
timestamp 1663859327
transform 1 0 403460 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_102
timestamp 1663859327
transform 1 0 404656 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_103
timestamp 1663859327
transform -1 0 403368 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_104
timestamp 1663859327
transform -1 0 404564 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_105
timestamp 1663859327
transform -1 0 405760 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_106
timestamp 1663859327
transform -1 0 406956 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_107
timestamp 1663859327
transform 1 0 405852 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_116
timestamp 1663859327
transform 1 0 407048 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_117
timestamp 1663859327
transform -1 0 408152 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_118
timestamp 1663859327
transform -1 0 409348 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_119
timestamp 1663859327
transform 1 0 408244 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_120
timestamp 1663859327
transform -1 0 410544 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_121
timestamp 1663859327
transform 1 0 409440 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_122
timestamp 1663859327
transform 1 0 410636 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_123
timestamp 1663859327
transform -1 0 411740 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_124
timestamp 1663859327
transform 1 0 411832 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_125
timestamp 1663859327
transform -1 0 414132 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_126
timestamp 1663859327
transform -1 0 412936 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_127
timestamp 1663859327
transform -1 0 414132 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_128
timestamp 1663859327
transform 0 -1 40864 -1 0 335777
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_129
timestamp 1663859327
transform 0 1 39776 1 0 334673
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_130
timestamp 1663859327
transform 0 -1 40864 -1 0 336973
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_131
timestamp 1663859327
transform 0 1 39776 1 0 335869
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_132
timestamp 1663859327
transform 0 -1 40864 -1 0 338169
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_133
timestamp 1663859327
transform 0 1 39776 1 0 337065
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_134
timestamp 1663859327
transform 0 -1 40864 -1 0 341757
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_135
timestamp 1663859327
transform 0 1 39776 1 0 340653
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_136
timestamp 1663859327
transform 0 -1 40864 -1 0 340561
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_137
timestamp 1663859327
transform 0 1 39776 1 0 339457
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_138
timestamp 1663859327
transform 0 1 39776 1 0 338261
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_139
timestamp 1663859327
transform 0 -1 40864 -1 0 339365
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_140
timestamp 1663859327
transform 0 1 39776 1 0 343045
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_141
timestamp 1663859327
transform 0 -1 40864 -1 0 344149
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_142
timestamp 1663859327
transform 0 1 39776 1 0 341849
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_143
timestamp 1663859327
transform 0 -1 40864 -1 0 342953
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_146
timestamp 1663859327
transform 0 1 39776 1 0 345437
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_147
timestamp 1663859327
transform 0 -1 40864 -1 0 346541
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_148
timestamp 1663859327
transform 0 1 39776 1 0 344241
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_149
timestamp 1663859327
transform 0 -1 40864 -1 0 345345
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_168
timestamp 1663859327
transform 0 1 39754 1 0 603618
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_169
timestamp 1663859327
transform 0 -1 40842 -1 0 604722
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_170
timestamp 1663859327
transform 0 1 39754 1 0 602422
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_171
timestamp 1663859327
transform 0 -1 40842 -1 0 603526
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_172
timestamp 1663859327
transform 0 -1 40842 -1 0 602330
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_173
timestamp 1663859327
transform 0 1 39754 1 0 601226
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_174
timestamp 1663859327
transform 0 1 39754 1 0 600030
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_175
timestamp 1663859327
transform 0 -1 40842 -1 0 601134
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_176
timestamp 1663859327
transform 0 1 39754 1 0 598834
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_177
timestamp 1663859327
transform 0 -1 40842 -1 0 599938
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_178
timestamp 1663859327
transform 0 1 39754 1 0 597638
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_179
timestamp 1663859327
transform 0 -1 40842 -1 0 598742
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 0 -1 677805 -1 0 707304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1663859327
transform 0 -1 677805 -1 0 708500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1663859327
transform -1 0 133892 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1663859327
transform -1 0 150636 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1663859327
transform -1 0 150636 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1663859327
transform -1 0 148244 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1663859327
transform -1 0 148244 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1663859327
transform -1 0 151832 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1663859327
transform -1 0 151832 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1663859327
transform -1 0 153028 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1663859327
transform -1 0 153028 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1663859327
transform -1 0 154224 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1663859327
transform -1 0 154224 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1663859327
transform 0 1 676717 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1663859327
transform 0 -1 677805 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1663859327
transform 0 1 676717 -1 0 707304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1663859327
transform 0 1 676717 -1 0 708500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1663859327
transform 0 1 676717 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1663859327
transform 0 -1 677805 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1663859327
transform 0 -1 677805 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1663859327
transform 0 1 676717 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1663859327
transform 0 -1 677805 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1663859327
transform 0 1 676717 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1663859327
transform 0 -1 677805 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1663859327
transform 0 1 676717 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1663859327
transform 0 -1 677805 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1663859327
transform 0 1 676717 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1663859327
transform 0 -1 677805 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1663859327
transform 0 1 676717 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1663859327
transform 0 -1 677805 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1663859327
transform 0 1 676717 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1663859327
transform -1 0 147048 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1663859327
transform -1 0 147048 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1663859327
transform -1 0 145852 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1663859327
transform -1 0 145852 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1663859327
transform -1 0 144656 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1663859327
transform -1 0 144656 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1663859327
transform -1 0 143460 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1663859327
transform -1 0 143460 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1663859327
transform -1 0 142264 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1663859327
transform -1 0 142264 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1663859327
transform -1 0 141068 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1663859327
transform -1 0 141068 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1663859327
transform -1 0 139872 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1663859327
transform -1 0 139872 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1663859327
transform -1 0 138676 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1663859327
transform -1 0 138676 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1663859327
transform -1 0 137480 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1663859327
transform -1 0 137480 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1663859327
transform -1 0 136284 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1663859327
transform -1 0 136284 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1663859327
transform -1 0 135088 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1663859327
transform -1 0 135088 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1663859327
transform -1 0 149440 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1663859327
transform -1 0 149440 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1663859327
transform -1 0 393892 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1663859327
transform -1 0 395088 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1663859327
transform -1 0 395088 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1663859327
transform -1 0 396284 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1663859327
transform -1 0 396284 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1663859327
transform -1 0 398676 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1663859327
transform -1 0 398676 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1663859327
transform -1 0 397480 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1663859327
transform -1 0 397480 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1663859327
transform -1 0 399872 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1663859327
transform -1 0 401068 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1663859327
transform -1 0 402264 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1663859327
transform -1 0 399872 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1663859327
transform -1 0 401068 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1663859327
transform -1 0 402264 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1663859327
transform -1 0 403460 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1663859327
transform -1 0 404656 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1663859327
transform -1 0 403460 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1663859327
transform -1 0 404656 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1663859327
transform -1 0 405852 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1663859327
transform -1 0 405852 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1663859327
transform -1 0 407048 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1663859327
transform -1 0 407048 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1663859327
transform -1 0 408244 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1663859327
transform -1 0 408244 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1663859327
transform -1 0 409440 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1663859327
transform -1 0 409440 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1663859327
transform -1 0 410636 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1663859327
transform -1 0 410636 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1663859327
transform -1 0 411832 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1663859327
transform -1 0 413028 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1663859327
transform -1 0 414224 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1663859327
transform -1 0 411832 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1663859327
transform -1 0 413028 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1663859327
transform -1 0 414224 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1663859327
transform 0 -1 40864 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1663859327
transform 0 1 39776 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1663859327
transform 0 -1 40864 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1663859327
transform 0 1 39776 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1663859327
transform 0 -1 40864 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1663859327
transform 0 1 39776 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1663859327
transform 0 1 39776 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1663859327
transform 0 -1 40864 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1663859327
transform 0 1 39776 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1663859327
transform 0 -1 40864 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1663859327
transform 0 1 39776 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1663859327
transform 0 -1 40864 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1663859327
transform 0 -1 40864 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1663859327
transform 0 1 39776 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1663859327
transform 0 -1 40864 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1663859327
transform 0 1 39776 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1663859327
transform 0 -1 40864 -1 0 346633
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1663859327
transform 0 1 39776 -1 0 346633
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1663859327
transform 0 -1 40864 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1663859327
transform 0 1 39776 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1663859327
transform 0 -1 40864 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1663859327
transform 0 1 39776 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_182
timestamp 1663859327
transform 0 1 39754 -1 0 604814
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_183
timestamp 1663859327
transform 0 -1 40842 -1 0 604814
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1663859327
transform 0 1 39754 -1 0 603618
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1663859327
transform 0 -1 40842 -1 0 603618
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1663859327
transform 0 -1 40842 -1 0 602422
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1663859327
transform 0 1 39754 -1 0 602422
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1663859327
transform 0 1 39754 -1 0 601226
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1663859327
transform 0 -1 40842 -1 0 601226
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1663859327
transform 0 1 39754 -1 0 598834
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1663859327
transform 0 1 39754 -1 0 600030
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1663859327
transform 0 -1 40842 -1 0 598834
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1663859327
transform 0 -1 40842 -1 0 600030
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1663859327
transform 0 1 39754 -1 0 597638
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1663859327
transform 0 -1 40842 -1 0 597638
box -38 -48 130 592
<< labels >>
flabel metal1 133123 223608 133374 223636 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[37]
port 93 nsew signal output
flabel metal3 146226 221997 146532 222091 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 147432 221997 147738 222091 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 405051 221984 405357 222078 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 406244 221978 406550 222072 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 39436 343400 39526 343697 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 39434 342201 39524 342498 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 39413 604045 39503 604342 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 678062 446931 678152 447228 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal1 132923 223664 133174 223692 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[36]
port 92 nsew signal output
flabel metal1 132723 223720 132974 223748 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[35]
port 91 nsew signal output
flabel metal1 132523 223776 132774 223804 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[37]
port 87 nsew signal input
flabel metal1 132323 223832 132574 223860 0 FreeSans 288 0 0 0 mgmt_io_out_buf[37]
port 86 nsew signal output
flabel metal1 132123 223888 132374 223916 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[36]
port 88 nsew signal input
flabel metal1 131923 223944 132174 223972 0 FreeSans 288 0 0 0 mgmt_io_out_buf[36]
port 85 nsew signal output
flabel metal1 131723 224000 131974 224028 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[35]
port 89 nsew signal input
flabel metal1 131523 224056 131774 224084 0 FreeSans 288 0 0 0 mgmt_io_out_buf[35]
port 84 nsew signal output
flabel metal1 131323 224112 131574 224140 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[34]
port 90 nsew signal input
flabel metal1 131123 224168 131374 224196 0 FreeSans 288 0 0 0 mgmt_io_out_buf[34]
port 83 nsew signal output
flabel metal3 39413 602844 39503 603141 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 678064 445738 678154 446035 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 678061 706542 678151 706839 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 678070 707739 678160 708036 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal1 41819 611095 41847 611356 0 FreeSans 288 90 0 0 mgmt_io_out_buf[29]
port 67 nsew signal output
flabel metal1 42183 353236 42211 353530 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[33]
port 78 nsew signal input
flabel metal1 42127 353436 42155 353730 0 FreeSans 288 90 0 0 mgmt_io_out_buf[32]
port 76 nsew signal output
flabel metal1 42071 353636 42099 353930 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[32]
port 79 nsew signal input
flabel metal1 42015 353836 42043 354130 0 FreeSans 288 90 0 0 mgmt_io_out_buf[31]
port 75 nsew signal output
flabel metal1 41959 354036 41987 354330 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[31]
port 80 nsew signal input
flabel metal1 41903 354236 41931 354530 0 FreeSans 288 90 0 0 mgmt_io_out_buf[30]
port 74 nsew signal output
flabel metal1 41847 354436 41875 354730 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[30]
port 81 nsew signal input
flabel metal1 41763 611295 41791 611556 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[29]
port 68 nsew signal input
flabel metal1 41707 611495 41735 611756 0 FreeSans 288 90 0 0 mgmt_io_out_buf[28]
port 66 nsew signal output
flabel metal1 41651 611695 41679 611956 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[28]
port 69 nsew signal input
flabel metal1 41595 611895 41623 612156 0 FreeSans 288 90 0 0 mgmt_io_out_buf[27]
port 65 nsew signal output
flabel metal1 41539 612095 41567 612356 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[27]
port 70 nsew signal input
flabel metal1 41483 612295 41511 612556 0 FreeSans 288 90 0 0 mgmt_io_out_buf[26]
port 64 nsew signal output
flabel metal1 41427 612495 41455 612756 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[26]
port 71 nsew signal input
flabel metal1 41371 612695 41399 612956 0 FreeSans 288 90 0 0 mgmt_io_out_buf[25]
port 63 nsew signal output
flabel metal1 41315 612895 41343 613156 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[25]
port 72 nsew signal input
flabel metal1 41259 613095 41287 613356 0 FreeSans 288 90 0 0 mgmt_io_out_buf[24]
port 62 nsew signal output
flabel metal1 41203 613295 41231 613556 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[24]
port 73 nsew signal input
flabel metal1 42239 353036 42267 353330 0 FreeSans 288 90 0 0 mgmt_io_out_buf[33]
port 77 nsew signal output
flabel metal1 676296 714634 676324 714921 0 FreeSans 288 90 0 0 mgmt_io_out_buf[13]
port 12 nsew signal output
flabel metal1 675624 453768 675652 454055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[7]
port 19 nsew signal output
flabel metal1 675652 215050 675680 215337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[7]
port 25 nsew signal input
flabel metal1 675540 215050 675568 215333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[33]
port 105 nsew signal input
flabel metal1 675708 214850 675736 215137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[7]
port 48 nsew signal output
flabel metal1 675764 214650 675792 214937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[8]
port 26 nsew signal input
flabel metal1 675820 214450 675848 214737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[8]
port 47 nsew signal output
flabel metal1 675876 214250 675904 214537 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[9]
port 27 nsew signal input
flabel metal1 675932 214050 675960 214337 0 FreeSans 288 90 0 0 mgmt_io_in_buf[9]
port 46 nsew signal output
flabel metal1 675988 213850 676016 214137 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[10]
port 28 nsew signal input
flabel metal1 676044 213650 676072 213937 0 FreeSans 288 90 0 0 mgmt_io_in_buf[10]
port 45 nsew signal output
flabel metal1 676100 213450 676128 213737 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[11]
port 29 nsew signal input
flabel metal1 676156 213250 676184 213537 0 FreeSans 288 90 0 0 mgmt_io_in_buf[11]
port 44 nsew signal output
flabel metal1 676212 213050 676240 213337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[12]
port 30 nsew signal input
flabel metal1 676268 212850 676296 213137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[12]
port 43 nsew signal output
flabel metal1 676324 212650 676352 212937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[13]
port 31 nsew signal input
flabel metal1 676380 212450 676408 212737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[13]
port 42 nsew signal output
flabel metal1 675484 215250 675512 215533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[33]
port 134 nsew signal output
flabel metal1 675428 215450 675456 215733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[32]
port 106 nsew signal input
flabel metal1 675372 215650 675400 215933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[32]
port 133 nsew signal output
flabel metal1 675316 215850 675344 216133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[31]
port 107 nsew signal input
flabel metal1 675260 216050 675288 216333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[31]
port 132 nsew signal output
flabel metal1 675204 216250 675232 216533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[30]
port 108 nsew signal input
flabel metal1 675148 216450 675176 216733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[30]
port 131 nsew signal output
flabel metal1 675092 216650 675120 216933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[29]
port 109 nsew signal input
flabel metal1 675036 216850 675064 217133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[29]
port 130 nsew signal output
flabel metal1 674980 217050 675008 217333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[28]
port 110 nsew signal input
flabel metal1 674924 217250 674952 217533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[28]
port 129 nsew signal output
flabel metal1 674868 217450 674896 217733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[27]
port 111 nsew signal input
flabel metal1 674812 217650 674840 217933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[27]
port 128 nsew signal output
flabel metal1 674756 217850 674784 218133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[26]
port 112 nsew signal input
flabel metal1 674700 218050 674728 218333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[26]
port 127 nsew signal output
flabel metal1 674644 218250 674672 218533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[25]
port 113 nsew signal input
flabel metal1 674588 218450 674616 218733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[25]
port 126 nsew signal output
flabel metal1 674532 218650 674560 218933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[24]
port 114 nsew signal input
flabel metal1 674476 218850 674504 219133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[24]
port 125 nsew signal output
flabel metal1 676352 714834 676380 715121 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[13]
port 10 nsew signal input
flabel metal1 675680 453968 675708 454255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[7]
port 18 nsew signal input
flabel metal1 675736 454168 675764 454455 0 FreeSans 288 90 0 0 mgmt_io_out_buf[8]
port 20 nsew signal output
flabel metal1 675792 454368 675820 454655 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[8]
port 17 nsew signal input
flabel metal1 675848 454568 675876 454855 0 FreeSans 288 90 0 0 mgmt_io_out_buf[9]
port 21 nsew signal output
flabel metal1 675904 454768 675932 455055 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[9]
port 16 nsew signal input
flabel metal1 675960 454968 675988 455255 0 FreeSans 288 90 0 0 mgmt_io_out_buf[10]
port 22 nsew signal output
flabel metal1 676016 455168 676044 455455 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[10]
port 15 nsew signal input
flabel metal1 676072 455368 676100 455655 0 FreeSans 288 90 0 0 mgmt_io_out_buf[11]
port 23 nsew signal output
flabel metal1 676128 455568 676156 455855 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[11]
port 14 nsew signal input
flabel metal1 676184 455768 676212 456055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[12]
port 24 nsew signal output
flabel metal1 676240 455968 676268 456255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[12]
port 13 nsew signal input
flabel metal1 673860 221050 673888 221287 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[37]
port 94 nsew signal input
flabel metal1 674420 219050 674448 219287 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[34]
port 101 nsew signal input
flabel metal1 674364 219250 674392 219487 0 FreeSans 288 90 0 0 mgmt_io_in_buf[34]
port 100 nsew signal output
flabel metal1 674308 219450 674336 219687 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[35]
port 102 nsew signal input
flabel metal1 674252 219650 674280 219887 0 FreeSans 288 90 0 0 mgmt_io_in_buf[35]
port 99 nsew signal output
flabel metal1 674196 219850 674224 220087 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[36]
port 103 nsew signal input
flabel metal1 674140 220050 674168 220287 0 FreeSans 288 90 0 0 mgmt_io_in_buf[36]
port 98 nsew signal output
flabel metal1 674084 220250 674112 220487 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[37]
port 104 nsew signal input
flabel metal1 674028 220450 674056 220687 0 FreeSans 288 90 0 0 mgmt_io_in_buf[37]
port 97 nsew signal output
flabel metal1 673972 220650 674000 220887 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[35]
port 96 nsew signal input
flabel metal1 673916 220850 673944 221087 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[36]
port 95 nsew signal input
<< end >>
