magic
tech sky130A
magscale 1 2
timestamp 1637551221
<< isosubstrate >>
rect 1110 1538 2650 4514
<< locali >>
rect 5089 9435 5123 9537
rect 3709 8823 3743 8925
rect 9505 3519 9539 3689
<< viali >>
rect 1317 11305 1351 11339
rect 1777 11305 1811 11339
rect 5273 11305 5307 11339
rect 5549 11305 5583 11339
rect 5917 11305 5951 11339
rect 6285 11305 6319 11339
rect 6653 11305 6687 11339
rect 7021 11305 7055 11339
rect 7757 11305 7791 11339
rect 8125 11305 8159 11339
rect 2053 11237 2087 11271
rect 3433 11237 3467 11271
rect 4169 11237 4203 11271
rect 7481 11237 7515 11271
rect 8769 11237 8803 11271
rect 9229 11237 9263 11271
rect 1501 11101 1535 11135
rect 1593 11101 1627 11135
rect 1869 11101 1903 11135
rect 2145 11101 2179 11135
rect 2605 11101 2639 11135
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 3249 11101 3283 11135
rect 4353 11101 4387 11135
rect 4629 11101 4663 11135
rect 4997 11101 5031 11135
rect 5089 11101 5123 11135
rect 5365 11101 5399 11135
rect 5733 11101 5767 11135
rect 6193 11101 6227 11135
rect 6837 11101 6871 11135
rect 7297 11101 7331 11135
rect 7665 11101 7699 11135
rect 8309 11101 8343 11135
rect 8953 11101 8987 11135
rect 9045 11101 9079 11135
rect 3617 11033 3651 11067
rect 3801 11033 3835 11067
rect 3985 11033 4019 11067
rect 2329 10965 2363 10999
rect 2421 10965 2455 10999
rect 2697 10965 2731 10999
rect 3157 10965 3191 10999
rect 4445 10965 4479 10999
rect 4813 10965 4847 10999
rect 8493 10965 8527 10999
rect 1317 10761 1351 10795
rect 8953 10761 8987 10795
rect 4721 10693 4755 10727
rect 1501 10625 1535 10659
rect 1777 10625 1811 10659
rect 2053 10625 2087 10659
rect 2145 10625 2179 10659
rect 2421 10625 2455 10659
rect 3157 10625 3191 10659
rect 3801 10625 3835 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 4973 10625 5007 10659
rect 5273 10625 5307 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 6193 10625 6227 10659
rect 8033 10625 8067 10659
rect 8585 10625 8619 10659
rect 8769 10625 8803 10659
rect 9229 10625 9263 10659
rect 6561 10557 6595 10591
rect 9045 10557 9079 10591
rect 3617 10489 3651 10523
rect 4261 10489 4295 10523
rect 6009 10489 6043 10523
rect 8493 10489 8527 10523
rect 1593 10421 1627 10455
rect 1869 10421 1903 10455
rect 2329 10421 2363 10455
rect 3065 10421 3099 10455
rect 3249 10421 3283 10455
rect 3893 10421 3927 10455
rect 4813 10421 4847 10455
rect 5457 10421 5491 10455
rect 9413 10421 9447 10455
rect 8033 10217 8067 10251
rect 8401 10217 8435 10251
rect 9137 10217 9171 10251
rect 3433 10149 3467 10183
rect 9413 10149 9447 10183
rect 3709 10081 3743 10115
rect 6101 10081 6135 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 4077 10013 4111 10047
rect 5549 10013 5583 10047
rect 7941 10013 7975 10047
rect 9229 10013 9263 10047
rect 1968 9945 2002 9979
rect 6377 9945 6411 9979
rect 8769 9945 8803 9979
rect 8953 9945 8987 9979
rect 1593 9877 1627 9911
rect 6009 9877 6043 9911
rect 7849 9877 7883 9911
rect 1501 9673 1535 9707
rect 6837 9673 6871 9707
rect 2513 9605 2547 9639
rect 5549 9605 5583 9639
rect 5641 9605 5675 9639
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 2421 9537 2455 9571
rect 3065 9537 3099 9571
rect 4537 9537 4571 9571
rect 5089 9537 5123 9571
rect 5181 9537 5215 9571
rect 5365 9537 5399 9571
rect 5825 9537 5859 9571
rect 6193 9537 6227 9571
rect 6929 9537 6963 9571
rect 9045 9537 9079 9571
rect 2697 9469 2731 9503
rect 7205 9469 7239 9503
rect 7573 9469 7607 9503
rect 5089 9401 5123 9435
rect 7021 9401 7055 9435
rect 2329 9333 2363 9367
rect 4997 9333 5031 9367
rect 6009 9333 6043 9367
rect 9505 9333 9539 9367
rect 1317 9129 1351 9163
rect 2329 9129 2363 9163
rect 2605 9129 2639 9163
rect 3433 9129 3467 9163
rect 3985 9129 4019 9163
rect 4813 9129 4847 9163
rect 5273 9129 5307 9163
rect 9413 9129 9447 9163
rect 2973 9061 3007 9095
rect 5365 8993 5399 9027
rect 1501 8925 1535 8959
rect 1593 8925 1627 8959
rect 2045 8925 2079 8959
rect 2154 8925 2188 8959
rect 2421 8925 2455 8959
rect 2881 8925 2915 8959
rect 3157 8925 3191 8959
rect 3249 8925 3283 8959
rect 3709 8925 3743 8959
rect 3801 8925 3835 8959
rect 4169 8925 4203 8959
rect 5089 8925 5123 8959
rect 7389 8925 7423 8959
rect 8769 8925 8803 8959
rect 4905 8857 4939 8891
rect 5641 8857 5675 8891
rect 8125 8857 8159 8891
rect 1777 8789 1811 8823
rect 1869 8789 1903 8823
rect 2697 8789 2731 8823
rect 3709 8789 3743 8823
rect 7113 8789 7147 8823
rect 9505 8585 9539 8619
rect 1317 8449 1351 8483
rect 1593 8449 1627 8483
rect 6193 8449 6227 8483
rect 7113 8449 7147 8483
rect 7205 8449 7239 8483
rect 9045 8449 9079 8483
rect 2329 8381 2363 8415
rect 2605 8381 2639 8415
rect 4169 8381 4203 8415
rect 4445 8381 4479 8415
rect 5917 8381 5951 8415
rect 7573 8381 7607 8415
rect 1501 8245 1535 8279
rect 2237 8245 2271 8279
rect 4077 8245 4111 8279
rect 6837 8245 6871 8279
rect 6929 8245 6963 8279
rect 1501 8041 1535 8075
rect 4537 8041 4571 8075
rect 4813 8041 4847 8075
rect 8217 8041 8251 8075
rect 8585 7973 8619 8007
rect 5181 7905 5215 7939
rect 5549 7905 5583 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 3617 7837 3651 7871
rect 4353 7837 4387 7871
rect 4905 7837 4939 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 8769 7837 8803 7871
rect 1961 7769 1995 7803
rect 8401 7769 8435 7803
rect 3433 7701 3467 7735
rect 4261 7701 4295 7735
rect 5089 7701 5123 7735
rect 7481 7701 7515 7735
rect 9413 7701 9447 7735
rect 7481 7497 7515 7531
rect 1409 7429 1443 7463
rect 6193 7429 6227 7463
rect 1685 7361 1719 7395
rect 2605 7361 2639 7395
rect 4445 7361 4479 7395
rect 4997 7361 5031 7395
rect 5733 7361 5767 7395
rect 8033 7361 8067 7395
rect 9045 7361 9079 7395
rect 2329 7293 2363 7327
rect 2973 7293 3007 7327
rect 9137 7293 9171 7327
rect 9229 7293 9263 7327
rect 1593 7225 1627 7259
rect 4905 7225 4939 7259
rect 8677 7225 8711 7259
rect 5641 7157 5675 7191
rect 5917 7157 5951 7191
rect 8125 7157 8159 7191
rect 8493 7157 8527 7191
rect 1948 6953 1982 6987
rect 3433 6953 3467 6987
rect 5917 6953 5951 6987
rect 6193 6953 6227 6987
rect 6824 6953 6858 6987
rect 8401 6953 8435 6987
rect 1685 6817 1719 6851
rect 6561 6817 6595 6851
rect 9321 6817 9355 6851
rect 1409 6749 1443 6783
rect 3617 6749 3651 6783
rect 3985 6749 4019 6783
rect 5457 6749 5491 6783
rect 6009 6749 6043 6783
rect 8585 6749 8619 6783
rect 1593 6613 1627 6647
rect 6469 6613 6503 6647
rect 8309 6613 8343 6647
rect 8769 6613 8803 6647
rect 9137 6613 9171 6647
rect 9229 6613 9263 6647
rect 1501 6409 1535 6443
rect 1777 6409 1811 6443
rect 2237 6409 2271 6443
rect 4905 6409 4939 6443
rect 5917 6409 5951 6443
rect 9321 6409 9355 6443
rect 2697 6341 2731 6375
rect 1317 6273 1351 6307
rect 1593 6273 1627 6307
rect 1869 6273 1903 6307
rect 2145 6273 2179 6307
rect 4261 6273 4295 6307
rect 4997 6273 5031 6307
rect 5641 6273 5675 6307
rect 5733 6273 5767 6307
rect 6193 6273 6227 6307
rect 8769 6273 8803 6307
rect 9505 6273 9539 6307
rect 2421 6205 2455 6239
rect 6929 6205 6963 6239
rect 7297 6205 7331 6239
rect 2053 6069 2087 6103
rect 4169 6069 4203 6103
rect 6837 6069 6871 6103
rect 9229 6069 9263 6103
rect 1225 5865 1259 5899
rect 2237 5865 2271 5899
rect 3709 5865 3743 5899
rect 6285 5865 6319 5899
rect 6653 5865 6687 5899
rect 1501 5797 1535 5831
rect 2973 5797 3007 5831
rect 9413 5797 9447 5831
rect 4077 5729 4111 5763
rect 4537 5729 4571 5763
rect 6837 5729 6871 5763
rect 7113 5729 7147 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 2053 5661 2087 5695
rect 2329 5661 2363 5695
rect 2605 5661 2639 5695
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 3617 5661 3651 5695
rect 4261 5661 4295 5695
rect 6193 5661 6227 5695
rect 8769 5661 8803 5695
rect 2789 5593 2823 5627
rect 1777 5525 1811 5559
rect 2513 5525 2547 5559
rect 3433 5525 3467 5559
rect 6009 5525 6043 5559
rect 8585 5525 8619 5559
rect 5089 5321 5123 5355
rect 5549 5253 5583 5287
rect 3341 5185 3375 5219
rect 5365 5185 5399 5219
rect 6193 5185 6227 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 3617 5117 3651 5151
rect 5825 5117 5859 5151
rect 8125 5117 8159 5151
rect 8677 5117 8711 5151
rect 8861 5117 8895 5151
rect 8493 5049 8527 5083
rect 5733 4981 5767 5015
rect 9321 4981 9355 5015
rect 3985 4777 4019 4811
rect 4629 4777 4663 4811
rect 9505 4777 9539 4811
rect 6285 4641 6319 4675
rect 3433 4573 3467 4607
rect 3709 4573 3743 4607
rect 4353 4573 4387 4607
rect 4905 4573 4939 4607
rect 5917 4573 5951 4607
rect 8125 4573 8159 4607
rect 8769 4573 8803 4607
rect 8861 4573 8895 4607
rect 5733 4505 5767 4539
rect 6561 4505 6595 4539
rect 3617 4437 3651 4471
rect 4169 4437 4203 4471
rect 4813 4437 4847 4471
rect 5549 4437 5583 4471
rect 6101 4437 6135 4471
rect 8033 4437 8067 4471
rect 3341 4233 3375 4267
rect 6745 4233 6779 4267
rect 3525 4097 3559 4131
rect 3617 4097 3651 4131
rect 5457 4097 5491 4131
rect 6101 4097 6135 4131
rect 6837 4097 6871 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 9045 4097 9079 4131
rect 3985 4029 4019 4063
rect 7573 4029 7607 4063
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 8033 3961 8067 3995
rect 8493 3961 8527 3995
rect 5917 3893 5951 3927
rect 7481 3893 7515 3927
rect 8677 3893 8711 3927
rect 4261 3689 4295 3723
rect 4353 3689 4387 3723
rect 4721 3689 4755 3723
rect 5457 3689 5491 3723
rect 6101 3689 6135 3723
rect 9045 3689 9079 3723
rect 9505 3689 9539 3723
rect 3341 3621 3375 3655
rect 4997 3621 5031 3655
rect 6929 3553 6963 3587
rect 3525 3485 3559 3519
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 4537 3485 4571 3519
rect 4905 3485 4939 3519
rect 5181 3485 5215 3519
rect 5273 3485 5307 3519
rect 5917 3485 5951 3519
rect 6009 3485 6043 3519
rect 6561 3485 6595 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 9505 3485 9539 3519
rect 3617 3349 3651 3383
rect 5733 3349 5767 3383
rect 6469 3349 6503 3383
rect 8585 3349 8619 3383
rect 8861 3349 8895 3383
rect 9413 3349 9447 3383
rect 3617 3145 3651 3179
rect 3893 3145 3927 3179
rect 9045 3145 9079 3179
rect 7757 3077 7791 3111
rect 3801 3009 3835 3043
rect 4077 3009 4111 3043
rect 4353 3009 4387 3043
rect 4721 3009 4755 3043
rect 6193 3009 6227 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 9137 3009 9171 3043
rect 3525 2941 3559 2975
rect 6653 2941 6687 2975
rect 9321 2941 9355 2975
rect 7481 2873 7515 2907
rect 8493 2873 8527 2907
rect 7941 2805 7975 2839
rect 8677 2805 8711 2839
rect 3709 2601 3743 2635
rect 4261 2601 4295 2635
rect 4629 2601 4663 2635
rect 5457 2601 5491 2635
rect 6469 2601 6503 2635
rect 6653 2601 6687 2635
rect 6929 2601 6963 2635
rect 8861 2601 8895 2635
rect 9321 2601 9355 2635
rect 3893 2533 3927 2567
rect 4905 2533 4939 2567
rect 4077 2397 4111 2431
rect 4537 2397 4571 2431
rect 4813 2397 4847 2431
rect 5089 2397 5123 2431
rect 5273 2397 5307 2431
rect 5733 2397 5767 2431
rect 6009 2397 6043 2431
rect 6285 2397 6319 2431
rect 6837 2397 6871 2431
rect 7113 2397 7147 2431
rect 7665 2397 7699 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8033 2397 8067 2431
rect 8401 2397 8435 2431
rect 8769 2397 8803 2431
rect 9505 2397 9539 2431
rect 7481 2329 7515 2363
rect 4353 2261 4387 2295
rect 5917 2261 5951 2295
rect 6193 2261 6227 2295
rect 8217 2261 8251 2295
rect 8585 2261 8619 2295
rect 9229 2261 9263 2295
rect 3617 2057 3651 2091
rect 3893 2057 3927 2091
rect 4169 2057 4203 2091
rect 4721 2057 4755 2091
rect 7113 1989 7147 2023
rect 3525 1921 3559 1955
rect 3801 1921 3835 1955
rect 4077 1921 4111 1955
rect 4353 1921 4387 1955
rect 4629 1921 4663 1955
rect 4905 1921 4939 1955
rect 5181 1921 5215 1955
rect 7021 1921 7055 1955
rect 8125 1921 8159 1955
rect 8585 1921 8619 1955
rect 8861 1921 8895 1955
rect 9137 1921 9171 1955
rect 9229 1921 9263 1955
rect 7849 1853 7883 1887
rect 4445 1785 4479 1819
rect 4997 1785 5031 1819
rect 8401 1785 8435 1819
rect 8953 1785 8987 1819
rect 9413 1785 9447 1819
rect 3341 1717 3375 1751
rect 7481 1717 7515 1751
rect 7941 1717 7975 1751
rect 8677 1717 8711 1751
rect 7665 1513 7699 1547
rect 8309 1513 8343 1547
rect 9137 1377 9171 1411
rect 3525 1309 3559 1343
rect 7849 1309 7883 1343
rect 8493 1309 8527 1343
rect 8861 1309 8895 1343
rect 8953 1309 8987 1343
rect 9505 1309 9539 1343
rect 3341 1173 3375 1207
rect 9321 1173 9355 1207
<< metal1 >>
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 9490 12220 9496 12232
rect 2464 12192 9496 12220
rect 2464 12180 2470 12192
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 4338 12112 4344 12164
rect 4396 12152 4402 12164
rect 9398 12152 9404 12164
rect 4396 12124 9404 12152
rect 4396 12112 4402 12124
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 5810 12044 5816 12096
rect 5868 12084 5874 12096
rect 9306 12084 9312 12096
rect 5868 12056 9312 12084
rect 5868 12044 5874 12056
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 3050 11976 3056 12028
rect 3108 12016 3114 12028
rect 8754 12016 8760 12028
rect 3108 11988 8760 12016
rect 3108 11976 3114 11988
rect 8754 11976 8760 11988
rect 8812 11976 8818 12028
rect 4798 11908 4804 11960
rect 4856 11948 4862 11960
rect 8662 11948 8668 11960
rect 4856 11920 8668 11948
rect 4856 11908 4862 11920
rect 8662 11908 8668 11920
rect 8720 11908 8726 11960
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 3786 11880 3792 11892
rect 2832 11852 3792 11880
rect 2832 11840 2838 11852
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 8386 11880 8392 11892
rect 5040 11852 8392 11880
rect 5040 11840 5046 11852
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 13538 11880 13544 11892
rect 12406 11852 13544 11880
rect 1486 11772 1492 11824
rect 1544 11812 1550 11824
rect 6638 11812 6644 11824
rect 1544 11784 6644 11812
rect 1544 11772 1550 11784
rect 6638 11772 6644 11784
rect 6696 11772 6702 11824
rect 7006 11772 7012 11824
rect 7064 11812 7070 11824
rect 12406 11812 12434 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 7064 11784 12434 11812
rect 7064 11772 7070 11784
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 5810 11744 5816 11756
rect 2464 11716 5816 11744
rect 2464 11704 2470 11716
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 13814 11744 13820 11756
rect 5960 11716 13820 11744
rect 5960 11704 5966 11716
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 6822 11676 6828 11688
rect 2746 11648 6828 11676
rect 1302 11500 1308 11552
rect 1360 11540 1366 11552
rect 2746 11540 2774 11648
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 2958 11568 2964 11620
rect 3016 11608 3022 11620
rect 8110 11608 8116 11620
rect 3016 11580 8116 11608
rect 3016 11568 3022 11580
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 1360 11512 2774 11540
rect 1360 11500 1366 11512
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 6178 11540 6184 11552
rect 3292 11512 6184 11540
rect 3292 11500 3298 11512
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 8294 11540 8300 11552
rect 6788 11512 8300 11540
rect 6788 11500 6794 11512
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 1302 11336 1308 11348
rect 1263 11308 1308 11336
rect 1302 11296 1308 11308
rect 1360 11296 1366 11348
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11336 1823 11339
rect 3234 11336 3240 11348
rect 1811 11308 3240 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 3344 11308 5273 11336
rect 2041 11271 2099 11277
rect 2041 11237 2053 11271
rect 2087 11237 2099 11271
rect 2041 11231 2099 11237
rect 2056 11200 2084 11231
rect 2222 11228 2228 11280
rect 2280 11268 2286 11280
rect 3344 11268 3372 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 5534 11336 5540 11348
rect 5495 11308 5540 11336
rect 5261 11299 5319 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5902 11336 5908 11348
rect 5863 11308 5908 11336
rect 5902 11296 5908 11308
rect 5960 11296 5966 11348
rect 6086 11296 6092 11348
rect 6144 11336 6150 11348
rect 6273 11339 6331 11345
rect 6273 11336 6285 11339
rect 6144 11308 6285 11336
rect 6144 11296 6150 11308
rect 6273 11305 6285 11308
rect 6319 11336 6331 11339
rect 6638 11336 6644 11348
rect 6319 11308 6500 11336
rect 6599 11308 6644 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 2280 11240 3372 11268
rect 3421 11271 3479 11277
rect 2280 11228 2286 11240
rect 3421 11237 3433 11271
rect 3467 11237 3479 11271
rect 3421 11231 3479 11237
rect 4157 11271 4215 11277
rect 4157 11237 4169 11271
rect 4203 11268 4215 11271
rect 4338 11268 4344 11280
rect 4203 11240 4344 11268
rect 4203 11237 4215 11240
rect 4157 11231 4215 11237
rect 2682 11200 2688 11212
rect 1596 11172 2084 11200
rect 2148 11172 2688 11200
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 1596 11141 1624 11172
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1854 11132 1860 11144
rect 1815 11104 1860 11132
rect 1581 11095 1639 11101
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 2148 11141 2176 11172
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 3436 11200 3464 11231
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 6472 11268 6500 11308
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 7006 11336 7012 11348
rect 6967 11308 7012 11336
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7116 11308 7757 11336
rect 7116 11268 7144 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 8110 11336 8116 11348
rect 8071 11308 8116 11336
rect 7745 11299 7803 11305
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8680 11308 9674 11336
rect 5644 11240 6408 11268
rect 6472 11240 7144 11268
rect 7469 11271 7527 11277
rect 2976 11172 3464 11200
rect 3528 11172 5120 11200
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2314 11092 2320 11144
rect 2372 11092 2378 11144
rect 2406 11092 2412 11144
rect 2464 11132 2470 11144
rect 2593 11135 2651 11141
rect 2464 11104 2544 11132
rect 2464 11092 2470 11104
rect 2332 11064 2360 11092
rect 2516 11064 2544 11104
rect 2593 11101 2605 11135
rect 2639 11132 2651 11135
rect 2866 11132 2872 11144
rect 2639 11104 2774 11132
rect 2827 11104 2872 11132
rect 2639 11101 2651 11104
rect 2593 11095 2651 11101
rect 2746 11064 2774 11104
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 2976 11141 3004 11172
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3418 11132 3424 11144
rect 3283 11104 3424 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3418 11092 3424 11104
rect 3476 11142 3482 11144
rect 3528 11142 3556 11172
rect 3476 11114 3556 11142
rect 3476 11092 3482 11114
rect 3712 11104 4292 11132
rect 3050 11064 3056 11076
rect 2332 11036 2452 11064
rect 2516 11036 2636 11064
rect 2746 11036 3056 11064
rect 2314 10996 2320 11008
rect 2275 10968 2320 10996
rect 2314 10956 2320 10968
rect 2372 10956 2378 11008
rect 2424 11005 2452 11036
rect 2409 10999 2467 11005
rect 2409 10965 2421 10999
rect 2455 10965 2467 10999
rect 2608 10996 2636 11036
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 3510 11024 3516 11076
rect 3568 11064 3574 11076
rect 3605 11067 3663 11073
rect 3605 11064 3617 11067
rect 3568 11036 3617 11064
rect 3568 11024 3574 11036
rect 3605 11033 3617 11036
rect 3651 11033 3663 11067
rect 3605 11027 3663 11033
rect 2685 10999 2743 11005
rect 2685 10996 2697 10999
rect 2608 10968 2697 10996
rect 2409 10959 2467 10965
rect 2685 10965 2697 10968
rect 2731 10965 2743 10999
rect 2685 10959 2743 10965
rect 3145 10999 3203 11005
rect 3145 10965 3157 10999
rect 3191 10996 3203 10999
rect 3712 10996 3740 11104
rect 3789 11067 3847 11073
rect 3789 11033 3801 11067
rect 3835 11033 3847 11067
rect 3970 11064 3976 11076
rect 3931 11036 3976 11064
rect 3789 11027 3847 11033
rect 3191 10968 3740 10996
rect 3804 10996 3832 11027
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 4264 11064 4292 11104
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4617 11135 4675 11141
rect 4396 11104 4441 11132
rect 4396 11092 4402 11104
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4706 11132 4712 11144
rect 4663 11104 4712 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 4982 11132 4988 11144
rect 4943 11104 4988 11132
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5092 11141 5120 11172
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 5644 11132 5672 11240
rect 6380 11200 6408 11240
rect 7469 11237 7481 11271
rect 7515 11237 7527 11271
rect 7469 11231 7527 11237
rect 7374 11200 7380 11212
rect 6380 11172 7380 11200
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7484 11200 7512 11231
rect 8680 11200 8708 11308
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 8846 11268 8852 11280
rect 8803 11240 8852 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 9217 11271 9275 11277
rect 9217 11268 9229 11271
rect 9180 11240 9229 11268
rect 9180 11228 9186 11240
rect 9217 11237 9229 11240
rect 9263 11237 9275 11271
rect 9217 11231 9275 11237
rect 7484 11172 8708 11200
rect 9646 11200 9674 11308
rect 13630 11200 13636 11212
rect 9646 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 5399 11104 5672 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 5776 11104 5821 11132
rect 5776 11092 5782 11104
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 6052 11104 6193 11132
rect 6052 11092 6058 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 7282 11132 7288 11144
rect 7243 11104 7288 11132
rect 6825 11095 6883 11101
rect 6730 11064 6736 11076
rect 4264 11036 6736 11064
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 4062 10996 4068 11008
rect 3804 10968 4068 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 4433 10999 4491 11005
rect 4433 10965 4445 10999
rect 4479 10996 4491 10999
rect 4522 10996 4528 11008
rect 4479 10968 4528 10996
rect 4479 10965 4491 10968
rect 4433 10959 4491 10965
rect 4522 10956 4528 10968
rect 4580 10956 4586 11008
rect 4798 10996 4804 11008
rect 4759 10968 4804 10996
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 6840 10996 6868 11095
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7708 11104 7753 11132
rect 7708 11092 7714 11104
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8352 11104 8397 11132
rect 8352 11092 8358 11104
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 8941 11135 8999 11141
rect 8941 11134 8953 11135
rect 8864 11132 8953 11134
rect 8628 11106 8953 11132
rect 8628 11104 8892 11106
rect 8628 11092 8634 11104
rect 8941 11101 8953 11106
rect 8987 11101 8999 11135
rect 9033 11135 9091 11141
rect 9033 11120 9045 11135
rect 9079 11120 9091 11135
rect 8941 11095 8999 11101
rect 9030 11068 9036 11120
rect 9088 11068 9094 11120
rect 10410 11064 10416 11076
rect 9140 11036 10416 11064
rect 8294 10996 8300 11008
rect 6840 10968 8300 10996
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 8481 10999 8539 11005
rect 8481 10965 8493 10999
rect 8527 10996 8539 10999
rect 9140 10996 9168 11036
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 8527 10968 9168 10996
rect 8527 10965 8539 10968
rect 8481 10959 8539 10965
rect 920 10906 9844 10928
rect 920 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5194 10906
rect 5246 10854 5258 10906
rect 5310 10854 5322 10906
rect 5374 10854 9844 10906
rect 920 10832 9844 10854
rect 1305 10795 1363 10801
rect 1305 10761 1317 10795
rect 1351 10792 1363 10795
rect 1394 10792 1400 10804
rect 1351 10764 1400 10792
rect 1351 10761 1363 10764
rect 1305 10755 1363 10761
rect 1394 10752 1400 10764
rect 1452 10752 1458 10804
rect 2774 10792 2780 10804
rect 1504 10764 2780 10792
rect 1504 10665 1532 10764
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 2924 10764 8064 10792
rect 2924 10752 2930 10764
rect 1946 10684 1952 10736
rect 2004 10724 2010 10736
rect 2004 10696 2452 10724
rect 2004 10684 2010 10696
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 1780 10520 1808 10619
rect 2056 10588 2084 10619
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2424 10665 2452 10696
rect 2498 10684 2504 10736
rect 2556 10724 2562 10736
rect 4709 10727 4767 10733
rect 4709 10724 4721 10727
rect 2556 10696 4721 10724
rect 2556 10684 2562 10696
rect 4709 10693 4721 10696
rect 4755 10693 4767 10727
rect 4709 10687 4767 10693
rect 4798 10684 4804 10736
rect 4856 10724 4862 10736
rect 4856 10696 5304 10724
rect 4856 10684 4862 10696
rect 2409 10659 2467 10665
rect 2188 10628 2233 10656
rect 2188 10616 2194 10628
rect 2409 10625 2421 10659
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 3510 10656 3516 10668
rect 3191 10628 3516 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10656 3847 10659
rect 3878 10656 3884 10668
rect 3835 10628 3884 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 3878 10616 3884 10628
rect 3936 10656 3942 10668
rect 5276 10665 5304 10696
rect 6822 10684 6828 10736
rect 6880 10724 6886 10736
rect 6880 10696 6946 10724
rect 6880 10684 6886 10696
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 3936 10628 4353 10656
rect 3936 10616 3942 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4961 10659 5019 10665
rect 4961 10656 4973 10659
rect 4525 10619 4583 10625
rect 4724 10628 4973 10656
rect 2056 10560 4108 10588
rect 2498 10520 2504 10532
rect 1780 10492 2504 10520
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 2682 10480 2688 10532
rect 2740 10480 2746 10532
rect 3142 10480 3148 10532
rect 3200 10520 3206 10532
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 3200 10492 3617 10520
rect 3200 10480 3206 10492
rect 3605 10489 3617 10492
rect 3651 10489 3663 10523
rect 4080 10520 4108 10560
rect 4249 10523 4307 10529
rect 4249 10520 4261 10523
rect 4080 10492 4261 10520
rect 3605 10483 3663 10489
rect 4249 10489 4261 10492
rect 4295 10489 4307 10523
rect 4249 10483 4307 10489
rect 4540 10520 4568 10619
rect 4724 10600 4752 10628
rect 4961 10625 4973 10628
rect 5007 10625 5019 10659
rect 4961 10619 5019 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 5994 10656 6000 10668
rect 5859 10628 6000 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 4706 10548 4712 10600
rect 4764 10548 4770 10600
rect 5644 10588 5672 10619
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6178 10656 6184 10668
rect 6139 10628 6184 10656
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 8036 10665 8064 10764
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8812 10764 8953 10792
rect 8812 10752 8818 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 8260 10696 8800 10724
rect 8260 10684 8266 10696
rect 8772 10665 8800 10696
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8021 10619 8079 10625
rect 8128 10628 8585 10656
rect 5718 10588 5724 10600
rect 5000 10560 5724 10588
rect 5000 10520 5028 10560
rect 5718 10548 5724 10560
rect 5776 10588 5782 10600
rect 6086 10588 6092 10600
rect 5776 10560 6092 10588
rect 5776 10548 5782 10560
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6546 10588 6552 10600
rect 6507 10560 6552 10588
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 4540 10492 5028 10520
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 1857 10455 1915 10461
rect 1857 10452 1869 10455
rect 1728 10424 1869 10452
rect 1728 10412 1734 10424
rect 1857 10421 1869 10424
rect 1903 10421 1915 10455
rect 1857 10415 1915 10421
rect 2317 10455 2375 10461
rect 2317 10421 2329 10455
rect 2363 10452 2375 10455
rect 2700 10452 2728 10480
rect 3050 10452 3056 10464
rect 2363 10424 2728 10452
rect 3011 10424 3056 10452
rect 2363 10421 2375 10424
rect 2317 10415 2375 10421
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10452 3298 10464
rect 3881 10455 3939 10461
rect 3881 10452 3893 10455
rect 3292 10424 3893 10452
rect 3292 10412 3298 10424
rect 3881 10421 3893 10424
rect 3927 10452 3939 10455
rect 4062 10452 4068 10464
rect 3927 10424 4068 10452
rect 3927 10421 3939 10424
rect 3881 10415 3939 10421
rect 4062 10412 4068 10424
rect 4120 10452 4126 10464
rect 4540 10452 4568 10492
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 5997 10523 6055 10529
rect 5997 10520 6009 10523
rect 5132 10492 6009 10520
rect 5132 10480 5138 10492
rect 5997 10489 6009 10492
rect 6043 10489 6055 10523
rect 5997 10483 6055 10489
rect 7466 10480 7472 10532
rect 7524 10520 7530 10532
rect 8128 10520 8156 10628
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10656 9275 10659
rect 9582 10656 9588 10668
rect 9263 10628 9588 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 7524 10492 8156 10520
rect 8404 10560 9045 10588
rect 7524 10480 7530 10492
rect 4120 10424 4568 10452
rect 4801 10455 4859 10461
rect 4120 10412 4126 10424
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5350 10452 5356 10464
rect 4847 10424 5356 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 8110 10452 8116 10464
rect 5491 10424 8116 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8404 10452 8432 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 8481 10523 8539 10529
rect 8481 10489 8493 10523
rect 8527 10520 8539 10523
rect 9214 10520 9220 10532
rect 8527 10492 9220 10520
rect 8527 10489 8539 10492
rect 8481 10483 8539 10489
rect 9214 10480 9220 10492
rect 9272 10480 9278 10532
rect 8754 10452 8760 10464
rect 8404 10424 8760 10452
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 9030 10412 9036 10464
rect 9088 10452 9094 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9088 10424 9413 10452
rect 9088 10412 9094 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 1636 10220 5580 10248
rect 1636 10208 1642 10220
rect 2958 10140 2964 10192
rect 3016 10180 3022 10192
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 3016 10152 3433 10180
rect 3016 10140 3022 10152
rect 3421 10149 3433 10152
rect 3467 10149 3479 10183
rect 3421 10143 3479 10149
rect 2314 10072 2320 10124
rect 2372 10112 2378 10124
rect 3697 10115 3755 10121
rect 3697 10112 3709 10115
rect 2372 10084 3709 10112
rect 2372 10072 2378 10084
rect 3697 10081 3709 10084
rect 3743 10081 3755 10115
rect 4706 10112 4712 10124
rect 3697 10075 3755 10081
rect 3804 10084 4712 10112
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 3804 10044 3832 10084
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 4062 10044 4068 10056
rect 3252 10016 3832 10044
rect 4023 10016 4068 10044
rect 3252 9988 3280 10016
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 5552 10053 5580 10220
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 6822 10248 6828 10260
rect 6144 10220 6828 10248
rect 6144 10208 6150 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7466 10248 7472 10260
rect 7064 10220 7472 10248
rect 7064 10208 7070 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8021 10251 8079 10257
rect 8021 10248 8033 10251
rect 7576 10220 8033 10248
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 7576 10180 7604 10220
rect 8021 10217 8033 10220
rect 8067 10248 8079 10251
rect 8202 10248 8208 10260
rect 8067 10220 8208 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8386 10248 8392 10260
rect 8347 10220 8392 10248
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8628 10220 9137 10248
rect 8628 10208 8634 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 7432 10152 7604 10180
rect 7432 10140 7438 10152
rect 7926 10140 7932 10192
rect 7984 10180 7990 10192
rect 9401 10183 9459 10189
rect 9401 10180 9413 10183
rect 7984 10152 9413 10180
rect 7984 10140 7990 10152
rect 9401 10149 9413 10152
rect 9447 10149 9459 10183
rect 9401 10143 9459 10149
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6135 10084 8616 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 8588 10056 8616 10084
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 7800 10016 7941 10044
rect 7800 10004 7806 10016
rect 7929 10013 7941 10016
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 8628 10016 9229 10044
rect 8628 10004 8634 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 22278 10044 22284 10056
rect 13872 10016 22284 10044
rect 13872 10004 13878 10016
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 1956 9979 2014 9985
rect 1956 9945 1968 9979
rect 2002 9976 2014 9979
rect 2002 9948 2360 9976
rect 2002 9945 2014 9948
rect 1956 9939 2014 9945
rect 2332 9920 2360 9948
rect 2682 9936 2688 9988
rect 2740 9936 2746 9988
rect 3234 9936 3240 9988
rect 3292 9936 3298 9988
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 2314 9868 2320 9920
rect 2372 9868 2378 9920
rect 2590 9868 2596 9920
rect 2648 9908 2654 9920
rect 4448 9908 4476 9962
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6365 9979 6423 9985
rect 6365 9976 6377 9979
rect 5868 9948 6377 9976
rect 5868 9936 5874 9948
rect 6365 9945 6377 9948
rect 6411 9945 6423 9979
rect 6365 9939 6423 9945
rect 6822 9936 6828 9988
rect 6880 9936 6886 9988
rect 7650 9936 7656 9988
rect 7708 9976 7714 9988
rect 8757 9979 8815 9985
rect 8757 9976 8769 9979
rect 7708 9948 8769 9976
rect 7708 9936 7714 9948
rect 8757 9945 8769 9948
rect 8803 9945 8815 9979
rect 8757 9939 8815 9945
rect 8941 9979 8999 9985
rect 8941 9945 8953 9979
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 2648 9880 4476 9908
rect 2648 9868 2654 9880
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 5997 9911 6055 9917
rect 5997 9908 6009 9911
rect 4764 9880 6009 9908
rect 4764 9868 4770 9880
rect 5997 9877 6009 9880
rect 6043 9877 6055 9911
rect 5997 9871 6055 9877
rect 6178 9868 6184 9920
rect 6236 9908 6242 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 6236 9880 7849 9908
rect 6236 9868 6242 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 8956 9908 8984 9939
rect 8260 9880 8984 9908
rect 8260 9868 8266 9880
rect 920 9818 9844 9840
rect 920 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5194 9818
rect 5246 9766 5258 9818
rect 5310 9766 5322 9818
rect 5374 9766 9844 9818
rect 920 9744 9844 9766
rect 1489 9707 1547 9713
rect 1489 9673 1501 9707
rect 1535 9704 1547 9707
rect 2130 9704 2136 9716
rect 1535 9676 2136 9704
rect 1535 9673 1547 9676
rect 1489 9667 1547 9673
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 2314 9664 2320 9716
rect 2372 9704 2378 9716
rect 6178 9704 6184 9716
rect 2372 9676 6184 9704
rect 2372 9664 2378 9676
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6604 9676 6837 9704
rect 6604 9664 6610 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 7650 9704 7656 9716
rect 7248 9676 7656 9704
rect 7248 9664 7254 9676
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 1596 9608 1808 9636
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9568 1455 9571
rect 1596 9568 1624 9608
rect 1443 9540 1624 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 1596 9364 1624 9540
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1780 9568 1808 9608
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 2501 9639 2559 9645
rect 2501 9636 2513 9639
rect 1912 9608 2513 9636
rect 1912 9596 1918 9608
rect 2501 9605 2513 9608
rect 2547 9605 2559 9639
rect 2501 9599 2559 9605
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 5534 9636 5540 9648
rect 3384 9608 3450 9636
rect 5495 9608 5540 9636
rect 3384 9596 3390 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5629 9639 5687 9645
rect 5629 9605 5641 9639
rect 5675 9636 5687 9639
rect 6086 9636 6092 9648
rect 5675 9608 6092 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 6086 9596 6092 9608
rect 6144 9596 6150 9648
rect 2406 9568 2412 9580
rect 1780 9540 2412 9568
rect 1673 9531 1731 9537
rect 1688 9432 1716 9531
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 3050 9568 3056 9580
rect 3011 9540 3056 9568
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4396 9540 4537 9568
rect 4396 9528 4402 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 5123 9540 5181 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5316 9540 5365 9568
rect 5316 9528 5322 9540
rect 5353 9537 5365 9540
rect 5399 9568 5411 9571
rect 5718 9568 5724 9580
rect 5399 9540 5724 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5718 9528 5724 9540
rect 5776 9568 5782 9580
rect 6196 9577 6224 9664
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 9306 9636 9312 9648
rect 6420 9608 7236 9636
rect 8694 9608 9312 9636
rect 6420 9596 6426 9608
rect 5813 9571 5871 9577
rect 5813 9568 5825 9571
rect 5776 9540 5825 9568
rect 5776 9528 5782 9540
rect 5813 9537 5825 9540
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6914 9568 6920 9580
rect 6181 9531 6239 9537
rect 6656 9540 6920 9568
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2372 9472 2697 9500
rect 2372 9460 2378 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2958 9500 2964 9512
rect 2685 9463 2743 9469
rect 2792 9472 2964 9500
rect 2792 9432 2820 9472
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 6656 9500 6684 9540
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7208 9568 7236 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 7650 9568 7656 9580
rect 7208 9540 7656 9568
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9490 9568 9496 9580
rect 9079 9540 9496 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 4908 9472 6684 9500
rect 1688 9404 2820 9432
rect 1854 9364 1860 9376
rect 1596 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 2004 9336 2329 9364
rect 2004 9324 2010 9336
rect 2317 9333 2329 9336
rect 2363 9333 2375 9367
rect 2317 9327 2375 9333
rect 2406 9324 2412 9376
rect 2464 9364 2470 9376
rect 4908 9364 4936 9472
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6788 9472 7205 9500
rect 6788 9460 6794 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 8202 9500 8208 9512
rect 7607 9472 8208 9500
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 5123 9404 5488 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 2464 9336 4936 9364
rect 4985 9367 5043 9373
rect 2464 9324 2470 9336
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5350 9364 5356 9376
rect 5031 9336 5356 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 5460 9364 5488 9404
rect 5718 9392 5724 9444
rect 5776 9432 5782 9444
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 5776 9404 7021 9432
rect 5776 9392 5782 9404
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 5902 9364 5908 9376
rect 5460 9336 5908 9364
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 7098 9364 7104 9376
rect 6043 9336 7104 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 8352 9336 9505 9364
rect 8352 9324 8358 9336
rect 9493 9333 9505 9336
rect 9539 9333 9551 9367
rect 9493 9327 9551 9333
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 1210 9120 1216 9172
rect 1268 9160 1274 9172
rect 1305 9163 1363 9169
rect 1305 9160 1317 9163
rect 1268 9132 1317 9160
rect 1268 9120 1274 9132
rect 1305 9129 1317 9132
rect 1351 9129 1363 9163
rect 2130 9160 2136 9172
rect 1305 9123 1363 9129
rect 1596 9132 2136 9160
rect 1026 8916 1032 8968
rect 1084 8956 1090 8968
rect 1596 8965 1624 9132
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 2593 9163 2651 9169
rect 2593 9160 2605 9163
rect 2424 9132 2605 9160
rect 1946 9052 1952 9104
rect 2004 9052 2010 9104
rect 1489 8959 1547 8965
rect 1489 8956 1501 8959
rect 1084 8928 1501 8956
rect 1084 8916 1090 8928
rect 1489 8925 1501 8928
rect 1535 8925 1547 8959
rect 1489 8919 1547 8925
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 1971 8956 1999 9052
rect 2424 9024 2452 9132
rect 2593 9129 2605 9132
rect 2639 9129 2651 9163
rect 3418 9160 3424 9172
rect 2593 9123 2651 9129
rect 2700 9132 3424 9160
rect 2332 8996 2452 9024
rect 2033 8959 2091 8965
rect 2033 8956 2045 8959
rect 1971 8928 2045 8956
rect 2033 8925 2045 8928
rect 2079 8925 2091 8959
rect 2033 8919 2091 8925
rect 2142 8959 2200 8965
rect 2142 8925 2154 8959
rect 2188 8956 2200 8959
rect 2332 8956 2360 8996
rect 2188 8928 2360 8956
rect 2409 8959 2467 8965
rect 2188 8925 2200 8928
rect 2142 8919 2200 8925
rect 2409 8925 2421 8959
rect 2455 8956 2467 8959
rect 2498 8956 2504 8968
rect 2455 8928 2504 8956
rect 2455 8925 2467 8928
rect 2409 8919 2467 8925
rect 2498 8916 2504 8928
rect 2556 8956 2562 8968
rect 2700 8956 2728 9132
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 3973 9163 4031 9169
rect 3973 9160 3985 9163
rect 3660 9132 3985 9160
rect 3660 9120 3666 9132
rect 3973 9129 3985 9132
rect 4019 9129 4031 9163
rect 3973 9123 4031 9129
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4801 9163 4859 9169
rect 4801 9160 4813 9163
rect 4120 9132 4813 9160
rect 4120 9120 4126 9132
rect 4801 9129 4813 9132
rect 4847 9129 4859 9163
rect 4801 9123 4859 9129
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 5261 9163 5319 9169
rect 5261 9160 5273 9163
rect 4948 9132 5273 9160
rect 4948 9120 4954 9132
rect 5261 9129 5273 9132
rect 5307 9129 5319 9163
rect 5261 9123 5319 9129
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5408 9132 6684 9160
rect 5408 9120 5414 9132
rect 2961 9095 3019 9101
rect 2961 9061 2973 9095
rect 3007 9092 3019 9095
rect 3326 9092 3332 9104
rect 3007 9064 3332 9092
rect 3007 9061 3019 9064
rect 2961 9055 3019 9061
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 4154 9092 4160 9104
rect 3844 9064 4160 9092
rect 3844 9052 3850 9064
rect 4154 9052 4160 9064
rect 4212 9052 4218 9104
rect 6656 9092 6684 9132
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 8260 9132 9413 9160
rect 8260 9120 8266 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 8754 9092 8760 9104
rect 6656 9064 8760 9092
rect 8754 9052 8760 9064
rect 8812 9092 8818 9104
rect 9306 9092 9312 9104
rect 8812 9064 9312 9092
rect 8812 9052 8818 9064
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 3970 9024 3976 9036
rect 2884 8996 3976 9024
rect 2884 8965 2912 8996
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 8570 9024 8576 9036
rect 5399 8996 8576 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 2556 8928 2728 8956
rect 2869 8959 2927 8965
rect 2556 8916 2562 8928
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 2869 8919 2927 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3697 8959 3755 8965
rect 3292 8928 3337 8956
rect 3292 8916 3298 8928
rect 3697 8925 3709 8959
rect 3743 8956 3755 8959
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3743 8928 3801 8956
rect 3743 8925 3755 8928
rect 3697 8919 3755 8925
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 4120 8928 4169 8956
rect 4120 8916 4126 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5258 8956 5264 8968
rect 5123 8928 5264 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7282 8956 7288 8968
rect 6788 8928 7288 8956
rect 6788 8916 6794 8928
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 8754 8956 8760 8968
rect 7423 8928 8616 8956
rect 8715 8928 8760 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 1780 8888 1808 8916
rect 2222 8888 2228 8900
rect 1780 8860 2228 8888
rect 2222 8848 2228 8860
rect 2280 8848 2286 8900
rect 3326 8888 3332 8900
rect 2332 8860 3332 8888
rect 1118 8780 1124 8832
rect 1176 8820 1182 8832
rect 1486 8820 1492 8832
rect 1176 8792 1492 8820
rect 1176 8780 1182 8792
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8820 1915 8823
rect 2332 8820 2360 8860
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 4338 8888 4344 8900
rect 3620 8860 4344 8888
rect 1903 8792 2360 8820
rect 2685 8823 2743 8829
rect 1903 8789 1915 8792
rect 1857 8783 1915 8789
rect 2685 8789 2697 8823
rect 2731 8820 2743 8823
rect 3620 8820 3648 8860
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 4893 8891 4951 8897
rect 4893 8888 4905 8891
rect 4856 8860 4905 8888
rect 4856 8848 4862 8860
rect 4893 8857 4905 8860
rect 4939 8857 4951 8891
rect 4893 8851 4951 8857
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5902 8888 5908 8900
rect 5675 8860 5908 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 6932 8860 7604 8888
rect 2731 8792 3648 8820
rect 3697 8823 3755 8829
rect 2731 8789 2743 8792
rect 2685 8783 2743 8789
rect 3697 8789 3709 8823
rect 3743 8820 3755 8823
rect 6932 8820 6960 8860
rect 3743 8792 6960 8820
rect 7101 8823 7159 8829
rect 3743 8789 3755 8792
rect 3697 8783 3755 8789
rect 7101 8789 7113 8823
rect 7147 8820 7159 8823
rect 7466 8820 7472 8832
rect 7147 8792 7472 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 7576 8820 7604 8860
rect 7650 8848 7656 8900
rect 7708 8888 7714 8900
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 7708 8860 8125 8888
rect 7708 8848 7714 8860
rect 8113 8857 8125 8860
rect 8159 8888 8171 8891
rect 8202 8888 8208 8900
rect 8159 8860 8208 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 8588 8888 8616 8928
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 9674 8888 9680 8900
rect 8588 8860 9680 8888
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 8386 8820 8392 8832
rect 7576 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 920 8730 9844 8752
rect 920 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5194 8730
rect 5246 8678 5258 8730
rect 5310 8678 5322 8730
rect 5374 8678 9844 8730
rect 920 8656 9844 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1820 8588 7236 8616
rect 1820 8576 1826 8588
rect 1486 8508 1492 8560
rect 1544 8548 1550 8560
rect 2498 8548 2504 8560
rect 1544 8520 2504 8548
rect 1544 8508 1550 8520
rect 2498 8508 2504 8520
rect 2556 8508 2562 8560
rect 4430 8548 4436 8560
rect 3818 8520 4436 8548
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 6730 8548 6736 8560
rect 5658 8534 6736 8548
rect 5644 8520 6736 8534
rect 1305 8483 1363 8489
rect 1305 8449 1317 8483
rect 1351 8449 1363 8483
rect 1305 8443 1363 8449
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 1946 8480 1952 8492
rect 1627 8452 1952 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 1320 8412 1348 8443
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2222 8440 2228 8492
rect 2280 8440 2286 8492
rect 1762 8412 1768 8424
rect 1320 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2240 8412 2268 8440
rect 2096 8384 2268 8412
rect 2317 8415 2375 8421
rect 2096 8372 2102 8384
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 2958 8412 2964 8424
rect 2639 8384 2964 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 2332 8344 2360 8375
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 3620 8384 4169 8412
rect 1728 8316 2360 8344
rect 1728 8304 1734 8316
rect 1302 8236 1308 8288
rect 1360 8276 1366 8288
rect 1489 8279 1547 8285
rect 1489 8276 1501 8279
rect 1360 8248 1501 8276
rect 1360 8236 1366 8248
rect 1489 8245 1501 8248
rect 1535 8245 1547 8279
rect 2222 8276 2228 8288
rect 2183 8248 2228 8276
rect 1489 8239 1547 8245
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 2332 8276 2360 8316
rect 3620 8276 3648 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4890 8412 4896 8424
rect 4479 8384 4896 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 5644 8412 5672 8520
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5920 8452 6193 8480
rect 5920 8424 5948 8452
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 7098 8480 7104 8492
rect 7059 8452 7104 8480
rect 6181 8443 6239 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7208 8489 7236 8588
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 8536 8588 9505 8616
rect 8536 8576 8542 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 8662 8508 8668 8560
rect 8720 8508 8726 8560
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9398 8480 9404 8492
rect 9079 8452 9404 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 5902 8412 5908 8424
rect 5132 8384 5672 8412
rect 5863 8384 5908 8412
rect 5132 8372 5138 8384
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 5994 8372 6000 8424
rect 6052 8372 6058 8424
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 8202 8412 8208 8424
rect 7607 8384 8208 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 6012 8344 6040 8372
rect 5644 8316 6040 8344
rect 5644 8288 5672 8316
rect 2332 8248 3648 8276
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4120 8248 4165 8276
rect 4120 8236 4126 8248
rect 5626 8236 5632 8288
rect 5684 8236 5690 8288
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6052 8248 6837 8276
rect 6052 8236 6058 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 7006 8276 7012 8288
rect 6963 8248 7012 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 3234 8072 3240 8084
rect 1535 8044 3240 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 4488 8044 4537 8072
rect 4488 8032 4494 8044
rect 4525 8041 4537 8044
rect 4571 8041 4583 8075
rect 4525 8035 4583 8041
rect 4540 8004 4568 8035
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4672 8044 4813 8072
rect 4672 8032 4678 8044
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 8205 8075 8263 8081
rect 8205 8041 8217 8075
rect 8251 8072 8263 8075
rect 8754 8072 8760 8084
rect 8251 8044 8760 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 5074 8004 5080 8016
rect 4540 7976 5080 8004
rect 5074 7964 5080 7976
rect 5132 7964 5138 8016
rect 8570 8004 8576 8016
rect 8531 7976 8576 8004
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 1578 7896 1584 7948
rect 1636 7936 1642 7948
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 1636 7908 5181 7936
rect 1636 7896 1642 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7936 5595 7939
rect 5994 7936 6000 7948
rect 5583 7908 6000 7936
rect 5583 7905 5595 7908
rect 5537 7899 5595 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7837 1455 7871
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1397 7831 1455 7837
rect 1412 7800 1440 7831
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4120 7840 4353 7868
rect 4120 7828 4126 7840
rect 4341 7837 4353 7840
rect 4387 7868 4399 7871
rect 4798 7868 4804 7880
rect 4387 7840 4804 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 4893 7831 4951 7837
rect 1854 7800 1860 7812
rect 1412 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 1949 7803 2007 7809
rect 1949 7769 1961 7803
rect 1995 7769 2007 7803
rect 3234 7800 3240 7812
rect 3174 7772 3240 7800
rect 1949 7763 2007 7769
rect 934 7692 940 7744
rect 992 7732 998 7744
rect 1578 7732 1584 7744
rect 992 7704 1584 7732
rect 992 7692 998 7704
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 1964 7732 1992 7763
rect 3234 7760 3240 7772
rect 3292 7760 3298 7812
rect 3694 7760 3700 7812
rect 3752 7800 3758 7812
rect 4908 7800 4936 7831
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7524 7840 7573 7868
rect 7524 7828 7530 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8720 7840 8769 7868
rect 8720 7828 8726 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 8386 7800 8392 7812
rect 3752 7772 4936 7800
rect 6670 7772 8248 7800
rect 8347 7772 8392 7800
rect 3752 7760 3758 7772
rect 2590 7732 2596 7744
rect 1964 7704 2596 7732
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 3421 7735 3479 7741
rect 3421 7732 3433 7735
rect 2740 7704 3433 7732
rect 2740 7692 2746 7704
rect 3421 7701 3433 7704
rect 3467 7701 3479 7735
rect 3421 7695 3479 7701
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 4430 7732 4436 7744
rect 4295 7704 4436 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 5077 7735 5135 7741
rect 5077 7732 5089 7735
rect 4672 7704 5089 7732
rect 4672 7692 4678 7704
rect 5077 7701 5089 7704
rect 5123 7701 5135 7735
rect 5077 7695 5135 7701
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 7432 7704 7481 7732
rect 7432 7692 7438 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 8220 7732 8248 7772
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 8294 7732 8300 7744
rect 8220 7704 8300 7732
rect 7469 7695 7527 7701
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 8812 7704 9413 7732
rect 8812 7692 8818 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 920 7642 9844 7664
rect 920 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5194 7642
rect 5246 7590 5258 7642
rect 5310 7590 5322 7642
rect 5374 7590 9844 7642
rect 920 7568 9844 7590
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 1412 7500 7481 7528
rect 1412 7469 1440 7500
rect 7469 7497 7481 7500
rect 7515 7528 7527 7531
rect 8386 7528 8392 7540
rect 7515 7500 8392 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 1397 7463 1455 7469
rect 1397 7429 1409 7463
rect 1443 7429 1455 7463
rect 2222 7460 2228 7472
rect 1397 7423 1455 7429
rect 1688 7432 2228 7460
rect 1688 7401 1716 7432
rect 2222 7420 2228 7432
rect 2280 7420 2286 7472
rect 3326 7420 3332 7472
rect 3384 7420 3390 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 6181 7463 6239 7469
rect 4304 7432 6040 7460
rect 4304 7420 4310 7432
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 1673 7355 1731 7361
rect 2056 7364 2605 7392
rect 1302 7284 1308 7336
rect 1360 7324 1366 7336
rect 2056 7324 2084 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4522 7392 4528 7404
rect 4479 7364 4528 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 5902 7392 5908 7404
rect 5767 7364 5908 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 1360 7296 2084 7324
rect 2317 7327 2375 7333
rect 1360 7284 1366 7296
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2363 7296 2973 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 5000 7324 5028 7355
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6012 7392 6040 7432
rect 6181 7429 6193 7463
rect 6227 7460 6239 7463
rect 6822 7460 6828 7472
rect 6227 7432 6828 7460
rect 6227 7429 6239 7432
rect 6181 7423 6239 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 6012 7364 8033 7392
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8021 7355 8079 7361
rect 8312 7364 9045 7392
rect 2961 7287 3019 7293
rect 4632 7296 5028 7324
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 1670 7256 1676 7268
rect 1627 7228 1676 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 1670 7216 1676 7228
rect 1728 7216 1734 7268
rect 1946 7216 1952 7268
rect 2004 7256 2010 7268
rect 2682 7256 2688 7268
rect 2004 7228 2688 7256
rect 2004 7216 2010 7228
rect 2682 7216 2688 7228
rect 2740 7216 2746 7268
rect 4632 7200 4660 7296
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 6730 7324 6736 7336
rect 6236 7296 6736 7324
rect 6236 7284 6242 7296
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 8312 7324 8340 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 7064 7296 8340 7324
rect 7064 7284 7070 7296
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 8444 7296 9137 7324
rect 8444 7284 8450 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9272 7296 9317 7324
rect 9272 7284 9278 7296
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 6454 7256 6460 7268
rect 4939 7228 6460 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 8665 7259 8723 7265
rect 8665 7256 8677 7259
rect 7248 7228 8677 7256
rect 7248 7216 7254 7228
rect 8665 7225 8677 7228
rect 8711 7225 8723 7259
rect 8665 7219 8723 7225
rect 4614 7148 4620 7200
rect 4672 7148 4678 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5629 7191 5687 7197
rect 5629 7188 5641 7191
rect 5040 7160 5641 7188
rect 5040 7148 5046 7160
rect 5629 7157 5641 7160
rect 5675 7157 5687 7191
rect 5629 7151 5687 7157
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 6638 7188 6644 7200
rect 5951 7160 6644 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 8110 7188 8116 7200
rect 8071 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8481 7191 8539 7197
rect 8481 7157 8493 7191
rect 8527 7188 8539 7191
rect 9398 7188 9404 7200
rect 8527 7160 9404 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 1946 6993 1952 6996
rect 1936 6987 1952 6993
rect 1936 6953 1948 6987
rect 1936 6947 1952 6953
rect 1946 6944 1952 6947
rect 2004 6944 2010 6996
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 3016 6956 3433 6984
rect 3016 6944 3022 6956
rect 3421 6953 3433 6956
rect 3467 6984 3479 6987
rect 3602 6984 3608 6996
rect 3467 6956 3608 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 5902 6984 5908 6996
rect 5863 6956 5908 6984
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 6178 6984 6184 6996
rect 6139 6956 6184 6984
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 6812 6987 6870 6993
rect 6812 6953 6824 6987
rect 6858 6984 6870 6987
rect 7466 6984 7472 6996
rect 6858 6956 7472 6984
rect 6858 6953 6870 6956
rect 6812 6947 6870 6953
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 8352 6956 8401 6984
rect 8352 6944 8358 6956
rect 8389 6953 8401 6956
rect 8435 6953 8447 6987
rect 8389 6947 8447 6953
rect 7834 6876 7840 6928
rect 7892 6916 7898 6928
rect 8110 6916 8116 6928
rect 7892 6888 8116 6916
rect 7892 6876 7898 6888
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 8570 6876 8576 6928
rect 8628 6876 8634 6928
rect 1670 6848 1676 6860
rect 1631 6820 1676 6848
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 4338 6848 4344 6860
rect 2004 6820 4344 6848
rect 2004 6808 2010 6820
rect 4338 6808 4344 6820
rect 4396 6848 4402 6860
rect 4522 6848 4528 6860
rect 4396 6820 4528 6848
rect 4396 6808 4402 6820
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6914 6848 6920 6860
rect 6595 6820 6920 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6914 6808 6920 6820
rect 6972 6848 6978 6860
rect 8588 6848 8616 6876
rect 6972 6820 8616 6848
rect 6972 6808 6978 6820
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9272 6820 9321 6848
rect 9272 6808 9278 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 1486 6780 1492 6792
rect 1443 6752 1492 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 3602 6780 3608 6792
rect 3563 6752 3608 6780
rect 3602 6740 3608 6752
rect 3660 6740 3666 6792
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 8573 6783 8631 6789
rect 8573 6780 8585 6783
rect 8128 6752 8585 6780
rect 3234 6712 3240 6724
rect 3174 6684 3240 6712
rect 3234 6672 3240 6684
rect 3292 6672 3298 6724
rect 1210 6604 1216 6656
rect 1268 6644 1274 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1268 6616 1593 6644
rect 1268 6604 1274 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 4356 6644 4384 6698
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 7098 6712 7104 6724
rect 6604 6684 7104 6712
rect 6604 6672 6610 6684
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 7834 6672 7840 6724
rect 7892 6672 7898 6724
rect 2280 6616 4384 6644
rect 6457 6647 6515 6653
rect 2280 6604 2286 6616
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 8128 6644 8156 6752
rect 8573 6749 8585 6752
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 8536 6684 8800 6712
rect 8536 6672 8542 6684
rect 8294 6644 8300 6656
rect 6503 6616 8156 6644
rect 8255 6616 8300 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 8294 6604 8300 6616
rect 8352 6644 8358 6656
rect 8662 6644 8668 6656
rect 8352 6616 8668 6644
rect 8352 6604 8358 6616
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 8772 6653 8800 6684
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8996 6616 9137 6644
rect 8996 6604 9002 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9272 6616 9317 6644
rect 9272 6604 9278 6616
rect 920 6554 9844 6576
rect 920 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5194 6554
rect 5246 6502 5258 6554
rect 5310 6502 5322 6554
rect 5374 6502 9844 6554
rect 920 6480 9844 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1489 6443 1547 6449
rect 1489 6440 1501 6443
rect 1452 6412 1501 6440
rect 1452 6400 1458 6412
rect 1489 6409 1501 6412
rect 1535 6409 1547 6443
rect 1762 6440 1768 6452
rect 1723 6412 1768 6440
rect 1489 6403 1547 6409
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 1854 6400 1860 6452
rect 1912 6440 1918 6452
rect 2225 6443 2283 6449
rect 1912 6412 2176 6440
rect 1912 6400 1918 6412
rect 1305 6307 1363 6313
rect 1305 6273 1317 6307
rect 1351 6273 1363 6307
rect 1305 6267 1363 6273
rect 1320 6168 1348 6267
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1544 6276 1593 6304
rect 1544 6264 1550 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 1946 6304 1952 6316
rect 1903 6276 1952 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2148 6313 2176 6412
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 3694 6440 3700 6452
rect 2271 6412 3700 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 4028 6412 4905 6440
rect 4028 6400 4034 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 5902 6440 5908 6452
rect 5863 6412 5908 6440
rect 4893 6403 4951 6409
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 7190 6440 7196 6452
rect 6012 6412 7196 6440
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6372 2743 6375
rect 2958 6372 2964 6384
rect 2731 6344 2964 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 4798 6372 4804 6384
rect 3988 6344 4804 6372
rect 3988 6316 4016 6344
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 3752 6276 3818 6304
rect 3752 6264 3758 6276
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4430 6304 4436 6316
rect 4295 6276 4436 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 4982 6304 4988 6316
rect 4943 6276 4988 6304
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5592 6276 5641 6304
rect 5592 6264 5598 6276
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6012 6304 6040 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8938 6440 8944 6452
rect 8168 6412 8944 6440
rect 8168 6400 8174 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6409 9367 6443
rect 9309 6403 9367 6409
rect 9324 6372 9352 6403
rect 8418 6344 9352 6372
rect 5767 6276 6040 6304
rect 6181 6307 6239 6313
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6730 6304 6736 6316
rect 6227 6276 6736 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 8846 6304 8852 6316
rect 8803 6276 8852 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9490 6304 9496 6316
rect 9451 6276 9496 6304
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 2406 6236 2412 6248
rect 1728 6208 2412 6236
rect 1728 6196 1734 6208
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 3476 6208 6929 6236
rect 3476 6196 3482 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 7282 6236 7288 6248
rect 7243 6208 7288 6236
rect 6917 6199 6975 6205
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 5718 6168 5724 6180
rect 1320 6140 2268 6168
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 2130 6100 2136 6112
rect 2087 6072 2136 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 2240 6100 2268 6140
rect 4080 6140 5724 6168
rect 4080 6100 4108 6140
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 2240 6072 4108 6100
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 4614 6100 4620 6112
rect 4203 6072 4620 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6236 6072 6837 6100
rect 6236 6060 6242 6072
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 9030 6060 9036 6112
rect 9088 6100 9094 6112
rect 9217 6103 9275 6109
rect 9217 6100 9229 6103
rect 9088 6072 9229 6100
rect 9088 6060 9094 6072
rect 9217 6069 9229 6072
rect 9263 6069 9275 6103
rect 9217 6063 9275 6069
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 1213 5899 1271 5905
rect 1213 5865 1225 5899
rect 1259 5896 1271 5899
rect 1854 5896 1860 5908
rect 1259 5868 1860 5896
rect 1259 5865 1271 5868
rect 1213 5859 1271 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2225 5899 2283 5905
rect 2225 5865 2237 5899
rect 2271 5896 2283 5899
rect 3602 5896 3608 5908
rect 2271 5868 3608 5896
rect 2271 5865 2283 5868
rect 2225 5859 2283 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 5994 5896 6000 5908
rect 3752 5868 3797 5896
rect 3988 5868 6000 5896
rect 3752 5856 3758 5868
rect 1302 5788 1308 5840
rect 1360 5828 1366 5840
rect 1489 5831 1547 5837
rect 1489 5828 1501 5831
rect 1360 5800 1501 5828
rect 1360 5788 1366 5800
rect 1489 5797 1501 5800
rect 1535 5797 1547 5831
rect 2958 5828 2964 5840
rect 2919 5800 2964 5828
rect 1489 5791 1547 5797
rect 2958 5788 2964 5800
rect 3016 5788 3022 5840
rect 3712 5828 3740 5856
rect 3252 5800 3740 5828
rect 1688 5732 2544 5760
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 1578 5692 1584 5704
rect 1443 5664 1584 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 1688 5701 1716 5732
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1946 5692 1952 5704
rect 1907 5664 1952 5692
rect 1673 5655 1731 5661
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 1210 5584 1216 5636
rect 1268 5624 1274 5636
rect 2056 5624 2084 5655
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2188 5664 2329 5692
rect 2188 5652 2194 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 1268 5596 2084 5624
rect 2516 5624 2544 5732
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2958 5692 2964 5704
rect 2639 5664 2964 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 3252 5701 3280 5800
rect 3418 5760 3424 5772
rect 3344 5732 3424 5760
rect 3237 5695 3295 5701
rect 3108 5664 3153 5692
rect 3108 5652 3114 5664
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 2777 5627 2835 5633
rect 2777 5624 2789 5627
rect 2516 5596 2789 5624
rect 1268 5584 1274 5596
rect 2777 5593 2789 5596
rect 2823 5624 2835 5627
rect 3252 5624 3280 5655
rect 2823 5596 3280 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5556 1823 5559
rect 2222 5556 2228 5568
rect 1811 5528 2228 5556
rect 1811 5525 1823 5528
rect 1765 5519 1823 5525
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 3344 5556 3372 5732
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 3436 5680 3617 5692
rect 3418 5628 3424 5680
rect 3476 5664 3617 5680
rect 3476 5628 3482 5664
rect 3605 5661 3617 5664
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 3988 5692 4016 5868
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 6641 5899 6699 5905
rect 6641 5865 6653 5899
rect 6687 5896 6699 5899
rect 9490 5896 9496 5908
rect 6687 5868 9496 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4154 5760 4160 5772
rect 4111 5732 4160 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 4522 5760 4528 5772
rect 4483 5732 4528 5760
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 6288 5760 6316 5859
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 9401 5831 9459 5837
rect 9401 5828 9413 5831
rect 8260 5800 9413 5828
rect 8260 5788 8266 5800
rect 9401 5797 9413 5800
rect 9447 5797 9459 5831
rect 9401 5791 9459 5797
rect 6822 5760 6828 5772
rect 5644 5732 6684 5760
rect 6783 5732 6828 5760
rect 4246 5692 4252 5704
rect 3752 5664 4016 5692
rect 4207 5664 4252 5692
rect 3752 5652 3758 5664
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5644 5692 5672 5732
rect 5592 5678 5672 5692
rect 5592 5664 5658 5678
rect 5592 5652 5598 5664
rect 6086 5652 6092 5704
rect 6144 5692 6150 5704
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 6144 5664 6193 5692
rect 6144 5652 6150 5664
rect 6181 5661 6193 5664
rect 6227 5692 6239 5695
rect 6546 5692 6552 5704
rect 6227 5664 6552 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 6454 5624 6460 5636
rect 5920 5596 6460 5624
rect 2547 5528 3372 5556
rect 3421 5559 3479 5565
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 5920 5556 5948 5596
rect 6454 5584 6460 5596
rect 6512 5584 6518 5636
rect 6656 5624 6684 5732
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 8294 5760 8300 5772
rect 7147 5732 8300 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 16942 5760 16948 5772
rect 13872 5732 16948 5760
rect 13872 5720 13878 5732
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 8754 5692 8760 5704
rect 8715 5664 8760 5692
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 7558 5624 7564 5636
rect 6656 5596 7564 5624
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 3467 5528 5948 5556
rect 5997 5559 6055 5565
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 5997 5525 6009 5559
rect 6043 5556 6055 5559
rect 6546 5556 6552 5568
rect 6043 5528 6552 5556
rect 6043 5525 6055 5528
rect 5997 5519 6055 5525
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7190 5556 7196 5568
rect 6880 5528 7196 5556
rect 6880 5516 6886 5528
rect 7190 5516 7196 5528
rect 7248 5556 7254 5568
rect 8573 5559 8631 5565
rect 8573 5556 8585 5559
rect 7248 5528 8585 5556
rect 7248 5516 7254 5528
rect 8573 5525 8585 5528
rect 8619 5525 8631 5559
rect 8573 5519 8631 5525
rect 920 5466 9844 5488
rect 920 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 5194 5466
rect 5246 5414 5258 5466
rect 5310 5414 5322 5466
rect 5374 5414 9844 5466
rect 920 5392 9844 5414
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 4948 5324 5089 5352
rect 4948 5312 4954 5324
rect 5077 5321 5089 5324
rect 5123 5321 5135 5355
rect 5077 5315 5135 5321
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 9306 5352 9312 5364
rect 8812 5324 9312 5352
rect 8812 5312 8818 5324
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 1118 5244 1124 5296
rect 1176 5284 1182 5296
rect 2682 5284 2688 5296
rect 1176 5256 2688 5284
rect 1176 5244 1182 5256
rect 2682 5244 2688 5256
rect 2740 5244 2746 5296
rect 5534 5284 5540 5296
rect 4830 5256 5540 5284
rect 4908 5228 4936 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 7466 5284 7472 5296
rect 7314 5256 7472 5284
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 2406 5176 2412 5228
rect 2464 5216 2470 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 2464 5188 3341 5216
rect 2464 5176 2470 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2774 5148 2780 5160
rect 2096 5120 2780 5148
rect 2096 5108 2102 5120
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 3344 5012 3372 5179
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 5350 5216 5356 5228
rect 5311 5188 5356 5216
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5552 5216 5580 5244
rect 5994 5216 6000 5228
rect 5552 5188 6000 5216
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6178 5216 6184 5228
rect 6139 5188 6184 5216
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7156 5188 7665 5216
rect 7156 5176 7162 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7653 5179 7711 5185
rect 8128 5188 8309 5216
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 4614 5148 4620 5160
rect 3651 5120 4620 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5810 5148 5816 5160
rect 5771 5120 5816 5148
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 8128 5157 8156 5188
rect 8297 5185 8309 5188
rect 8343 5216 8355 5219
rect 8386 5216 8392 5228
rect 8343 5188 8392 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5117 8171 5151
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8113 5111 8171 5117
rect 8220 5120 8677 5148
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 8220 5080 8248 5120
rect 8665 5117 8677 5120
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9398 5148 9404 5160
rect 8895 5120 9404 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 7248 5052 8248 5080
rect 8481 5083 8539 5089
rect 7248 5040 7254 5052
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 13814 5080 13820 5092
rect 8527 5052 13820 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 4246 5012 4252 5024
rect 3344 4984 4252 5012
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5592 4984 5733 5012
rect 5592 4972 5598 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 9306 5012 9312 5024
rect 9267 4984 9312 5012
rect 5721 4975 5779 4981
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 3602 4768 3608 4820
rect 3660 4808 3666 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3660 4780 3985 4808
rect 3660 4768 3666 4780
rect 3973 4777 3985 4780
rect 4019 4808 4031 4811
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4019 4780 4629 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 4617 4777 4629 4780
rect 4663 4808 4675 4811
rect 4890 4808 4896 4820
rect 4663 4780 4896 4808
rect 4663 4777 4675 4780
rect 4617 4771 4675 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 7340 4780 9505 4808
rect 7340 4768 7346 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 5350 4740 5356 4752
rect 3712 4712 5356 4740
rect 1026 4564 1032 4616
rect 1084 4604 1090 4616
rect 3142 4604 3148 4616
rect 1084 4576 3148 4604
rect 1084 4564 1090 4576
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3418 4604 3424 4616
rect 3379 4576 3424 4604
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3712 4613 3740 4712
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 4614 4632 4620 4684
rect 4672 4672 4678 4684
rect 5626 4672 5632 4684
rect 4672 4644 5632 4672
rect 4672 4632 4678 4644
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6914 4672 6920 4684
rect 6319 4644 6920 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 8018 4672 8024 4684
rect 7892 4644 8024 4672
rect 7892 4632 7898 4644
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 3697 4607 3755 4613
rect 3697 4573 3709 4607
rect 3743 4573 3755 4607
rect 3697 4567 3755 4573
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 3712 4536 3740 4567
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 4304 4576 4353 4604
rect 4304 4564 4310 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5074 4604 5080 4616
rect 4939 4576 5080 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 2924 4508 3740 4536
rect 4356 4536 4384 4567
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 5994 4604 6000 4616
rect 5951 4576 6000 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 8036 4576 8125 4604
rect 5721 4539 5779 4545
rect 5721 4536 5733 4539
rect 4356 4508 5733 4536
rect 2924 4496 2930 4508
rect 5721 4505 5733 4508
rect 5767 4505 5779 4539
rect 6012 4536 6040 4564
rect 6546 4536 6552 4548
rect 6012 4508 6408 4536
rect 6507 4508 6552 4536
rect 5721 4499 5779 4505
rect 3602 4468 3608 4480
rect 3563 4440 3608 4468
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4522 4468 4528 4480
rect 4203 4440 4528 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 4798 4468 4804 4480
rect 4759 4440 4804 4468
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 5537 4471 5595 4477
rect 5537 4468 5549 4471
rect 5040 4440 5549 4468
rect 5040 4428 5046 4440
rect 5537 4437 5549 4440
rect 5583 4437 5595 4471
rect 6086 4468 6092 4480
rect 6047 4440 6092 4468
rect 5537 4431 5595 4437
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6380 4468 6408 4508
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 7024 4468 7052 4522
rect 8036 4480 8064 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 8803 4576 8861 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 7282 4468 7288 4480
rect 6380 4440 7288 4468
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 8018 4468 8024 4480
rect 7979 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 3036 4378 9844 4400
rect 3036 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 5194 4378
rect 5246 4326 5258 4378
rect 5310 4326 5322 4378
rect 5374 4326 9844 4378
rect 3036 4304 9844 4326
rect 3329 4267 3387 4273
rect 3329 4233 3341 4267
rect 3375 4264 3387 4267
rect 4246 4264 4252 4276
rect 3375 4236 4252 4264
rect 3375 4233 3387 4236
rect 3329 4227 3387 4233
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 6730 4264 6736 4276
rect 4764 4236 5212 4264
rect 6691 4236 6736 4264
rect 4764 4224 4770 4236
rect 4430 4156 4436 4208
rect 4488 4156 4494 4208
rect 5184 4196 5212 4236
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 9766 4264 9772 4276
rect 7524 4236 9772 4264
rect 7524 4224 7530 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 5258 4196 5264 4208
rect 5184 4168 5264 4196
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 8846 4156 8852 4208
rect 8904 4196 8910 4208
rect 8904 4168 9352 4196
rect 8904 4156 8910 4168
rect 3510 4128 3516 4140
rect 3471 4100 3516 4128
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 5442 4128 5448 4140
rect 3660 4100 3705 4128
rect 5403 4100 5448 4128
rect 3660 4088 3666 4100
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6546 4128 6552 4140
rect 6135 4100 6552 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6788 4100 6837 4128
rect 6788 4088 6794 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 7524 4100 8125 4128
rect 7524 4088 7530 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8570 4128 8576 4140
rect 8343 4100 8576 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8996 4100 9045 4128
rect 8996 4088 9002 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 3973 4063 4031 4069
rect 3973 4029 3985 4063
rect 4019 4060 4031 4063
rect 4614 4060 4620 4072
rect 4019 4032 4620 4060
rect 4019 4029 4031 4032
rect 3973 4023 4031 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 7561 4063 7619 4069
rect 7561 4029 7573 4063
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 7576 3992 7604 4023
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9324 4069 9352 4168
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8720 4032 9137 4060
rect 8720 4020 8726 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9582 4060 9588 4072
rect 9355 4032 9588 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 7742 3992 7748 4004
rect 7576 3964 7748 3992
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 7834 3952 7840 4004
rect 7892 3992 7898 4004
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 7892 3964 8033 3992
rect 7892 3952 7898 3964
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 13814 3992 13820 4004
rect 8527 3964 13820 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 5224 3896 5917 3924
rect 5224 3884 5230 3896
rect 5905 3893 5917 3896
rect 5951 3893 5963 3927
rect 5905 3887 5963 3893
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 6972 3896 7481 3924
rect 6972 3884 6978 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3924 8723 3927
rect 9214 3924 9220 3936
rect 8711 3896 9220 3924
rect 8711 3893 8723 3896
rect 8665 3887 8723 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 3476 3692 4261 3720
rect 3476 3680 3482 3692
rect 4249 3689 4261 3692
rect 4295 3689 4307 3723
rect 4249 3683 4307 3689
rect 4341 3723 4399 3729
rect 4341 3689 4353 3723
rect 4387 3720 4399 3723
rect 4430 3720 4436 3732
rect 4387 3692 4436 3720
rect 4387 3689 4399 3692
rect 4341 3683 4399 3689
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 4706 3720 4712 3732
rect 4667 3692 4712 3720
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3689 5503 3723
rect 5445 3683 5503 3689
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3652 3387 3655
rect 3602 3652 3608 3664
rect 3375 3624 3608 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 4614 3612 4620 3664
rect 4672 3652 4678 3664
rect 4985 3655 5043 3661
rect 4985 3652 4997 3655
rect 4672 3624 4997 3652
rect 4672 3612 4678 3624
rect 4985 3621 4997 3624
rect 5031 3621 5043 3655
rect 4985 3615 5043 3621
rect 5460 3596 5488 3683
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 6089 3723 6147 3729
rect 6089 3720 6101 3723
rect 6052 3692 6101 3720
rect 6052 3680 6058 3692
rect 6089 3689 6101 3692
rect 6135 3689 6147 3723
rect 6089 3683 6147 3689
rect 6196 3692 7880 3720
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 6196 3652 6224 3692
rect 5684 3624 6224 3652
rect 7852 3652 7880 3692
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8260 3692 8800 3720
rect 8260 3680 8266 3692
rect 8772 3652 8800 3692
rect 8956 3692 9045 3720
rect 8956 3652 8984 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 9493 3723 9551 3729
rect 9493 3720 9505 3723
rect 9272 3692 9505 3720
rect 9272 3680 9278 3692
rect 9493 3689 9505 3692
rect 9539 3689 9551 3723
rect 9493 3683 9551 3689
rect 13722 3652 13728 3664
rect 7852 3624 8708 3652
rect 8772 3624 8984 3652
rect 9048 3624 13728 3652
rect 5684 3612 5690 3624
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 3292 3556 3832 3584
rect 3292 3544 3298 3556
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3694 3516 3700 3528
rect 3559 3488 3700 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 3804 3525 3832 3556
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 4430 3584 4436 3596
rect 4304 3556 4436 3584
rect 4304 3544 4310 3556
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 4856 3556 5212 3584
rect 4856 3544 4862 3556
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 4338 3516 4344 3528
rect 4111 3488 4344 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 5184 3525 5212 3556
rect 5442 3544 5448 3596
rect 5500 3544 5506 3596
rect 6086 3584 6092 3596
rect 5920 3556 6092 3584
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 4908 3448 4936 3479
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5718 3516 5724 3528
rect 5316 3488 5361 3516
rect 5644 3488 5724 3516
rect 5316 3476 5322 3488
rect 5534 3448 5540 3460
rect 3620 3420 4752 3448
rect 4908 3420 5540 3448
rect 3620 3389 3648 3420
rect 3605 3383 3663 3389
rect 3605 3349 3617 3383
rect 3651 3349 3663 3383
rect 3605 3343 3663 3349
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 4062 3380 4068 3392
rect 3752 3352 4068 3380
rect 3752 3340 3758 3352
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4724 3380 4752 3420
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 5644 3380 5672 3488
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 5920 3525 5948 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6914 3584 6920 3596
rect 6875 3556 6920 3584
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 8680 3584 8708 3624
rect 9048 3584 9076 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 8680 3556 9076 3584
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 16574 3584 16580 3596
rect 9916 3556 16580 3584
rect 9916 3544 9922 3556
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 6546 3516 6552 3528
rect 6052 3488 6097 3516
rect 6507 3488 6552 3516
rect 6052 3476 6058 3488
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8404 3448 8432 3479
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 8941 3519 8999 3525
rect 8628 3488 8892 3516
rect 8628 3476 8634 3488
rect 8754 3448 8760 3460
rect 7392 3392 7420 3434
rect 8404 3420 8760 3448
rect 8754 3408 8760 3420
rect 8812 3408 8818 3460
rect 4724 3352 5672 3380
rect 5721 3383 5779 3389
rect 5721 3349 5733 3383
rect 5767 3380 5779 3383
rect 6178 3380 6184 3392
rect 5767 3352 6184 3380
rect 5767 3349 5779 3352
rect 5721 3343 5779 3349
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 6822 3380 6828 3392
rect 6503 3352 6828 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 7374 3340 7380 3392
rect 7432 3340 7438 3392
rect 8570 3380 8576 3392
rect 8531 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 8864 3389 8892 3488
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 8987 3488 9505 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 8849 3383 8907 3389
rect 8849 3349 8861 3383
rect 8895 3349 8907 3383
rect 8849 3343 8907 3349
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9490 3380 9496 3392
rect 9447 3352 9496 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 3036 3290 9844 3312
rect 3036 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 5194 3290
rect 5246 3238 5258 3290
rect 5310 3238 5322 3290
rect 5374 3238 9844 3290
rect 13814 3272 13820 3324
rect 13872 3312 13878 3324
rect 16758 3312 16764 3324
rect 13872 3284 16764 3312
rect 13872 3272 13878 3284
rect 16758 3272 16764 3284
rect 16816 3272 16822 3324
rect 3036 3216 9844 3238
rect 3605 3179 3663 3185
rect 3605 3145 3617 3179
rect 3651 3176 3663 3179
rect 3694 3176 3700 3188
rect 3651 3148 3700 3176
rect 3651 3145 3663 3148
rect 3605 3139 3663 3145
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 3844 3148 3893 3176
rect 3844 3136 3850 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 3881 3139 3939 3145
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4120 3148 7880 3176
rect 4120 3136 4126 3148
rect 3050 3068 3056 3120
rect 3108 3108 3114 3120
rect 3108 3080 4200 3108
rect 3108 3068 3114 3080
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 3804 2972 3832 3003
rect 3970 3000 3976 3052
rect 4028 3040 4034 3052
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 4028 3012 4077 3040
rect 4028 3000 4034 3012
rect 4065 3009 4077 3012
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 3559 2944 3832 2972
rect 4172 2972 4200 3080
rect 4982 3068 4988 3120
rect 5040 3108 5046 3120
rect 5040 3080 5106 3108
rect 5040 3068 5046 3080
rect 5994 3068 6000 3120
rect 6052 3108 6058 3120
rect 6052 3080 6960 3108
rect 6052 3068 6058 3080
rect 4338 3040 4344 3052
rect 4299 3012 4344 3040
rect 4338 3000 4344 3012
rect 4396 3000 4402 3052
rect 4522 3000 4528 3052
rect 4580 3040 4586 3052
rect 4709 3043 4767 3049
rect 4709 3040 4721 3043
rect 4580 3012 4721 3040
rect 4580 3000 4586 3012
rect 4709 3009 4721 3012
rect 4755 3009 4767 3043
rect 6178 3040 6184 3052
rect 6139 3012 6184 3040
rect 4709 3003 4767 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6932 3040 6960 3080
rect 7466 3068 7472 3120
rect 7524 3108 7530 3120
rect 7745 3111 7803 3117
rect 7745 3108 7757 3111
rect 7524 3080 7757 3108
rect 7524 3068 7530 3080
rect 7745 3077 7757 3080
rect 7791 3077 7803 3111
rect 7852 3108 7880 3148
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 9033 3179 9091 3185
rect 9033 3176 9045 3179
rect 8628 3148 9045 3176
rect 8628 3136 8634 3148
rect 9033 3145 9045 3148
rect 9079 3145 9091 3179
rect 13446 3176 13452 3188
rect 9033 3139 9091 3145
rect 9140 3148 13452 3176
rect 9140 3108 9168 3148
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 16850 3176 16856 3188
rect 13688 3148 16856 3176
rect 13688 3136 13694 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 7852 3080 9168 3108
rect 7745 3071 7803 3077
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 6932 3012 7573 3040
rect 6825 3003 6883 3009
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8260 3012 8309 3040
rect 8260 3000 8266 3012
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 8938 3040 8944 3052
rect 8628 3012 8944 3040
rect 8628 3000 8634 3012
rect 8938 3000 8944 3012
rect 8996 3044 9002 3052
rect 9125 3044 9183 3049
rect 8996 3043 9183 3044
rect 8996 3016 9137 3043
rect 8996 3000 9002 3016
rect 9125 3009 9137 3016
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 9232 3012 22094 3040
rect 5166 2972 5172 2984
rect 4172 2944 5172 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3804 2836 3832 2944
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 8110 2972 8116 2984
rect 6687 2944 8116 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 9232 2972 9260 3012
rect 8220 2944 9260 2972
rect 9309 2975 9367 2981
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 7469 2907 7527 2913
rect 7469 2904 7481 2907
rect 6512 2876 7481 2904
rect 6512 2864 6518 2876
rect 7469 2873 7481 2876
rect 7515 2873 7527 2907
rect 8220 2904 8248 2944
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 9766 2972 9772 2984
rect 9355 2944 9772 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 7469 2867 7527 2873
rect 7576 2876 8248 2904
rect 8481 2907 8539 2913
rect 7576 2836 7604 2876
rect 8481 2873 8493 2907
rect 8527 2904 8539 2907
rect 13814 2904 13820 2916
rect 8527 2876 13820 2904
rect 8527 2873 8539 2876
rect 8481 2867 8539 2873
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 22066 2904 22094 3012
rect 22186 2904 22192 2916
rect 22066 2876 22192 2904
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 3804 2808 7604 2836
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2836 7987 2839
rect 8202 2836 8208 2848
rect 7975 2808 8208 2836
rect 7975 2805 7987 2808
rect 7929 2799 7987 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8662 2836 8668 2848
rect 8623 2808 8668 2836
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 3510 2592 3516 2644
rect 3568 2632 3574 2644
rect 3697 2635 3755 2641
rect 3697 2632 3709 2635
rect 3568 2604 3709 2632
rect 3568 2592 3574 2604
rect 3697 2601 3709 2604
rect 3743 2632 3755 2635
rect 3970 2632 3976 2644
rect 3743 2604 3976 2632
rect 3743 2601 3755 2604
rect 3697 2595 3755 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4249 2635 4307 2641
rect 4249 2632 4261 2635
rect 4172 2604 4261 2632
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4062 2564 4068 2576
rect 3927 2536 4068 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4172 2428 4200 2604
rect 4249 2601 4261 2604
rect 4295 2632 4307 2635
rect 4522 2632 4528 2644
rect 4295 2604 4528 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 5166 2632 5172 2644
rect 4663 2604 5172 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5810 2632 5816 2644
rect 5491 2604 5816 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 6457 2635 6515 2641
rect 6457 2601 6469 2635
rect 6503 2632 6515 2635
rect 6546 2632 6552 2644
rect 6503 2604 6552 2632
rect 6503 2601 6515 2604
rect 6457 2595 6515 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 6641 2635 6699 2641
rect 6641 2601 6653 2635
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7098 2632 7104 2644
rect 6963 2604 7104 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 4430 2524 4436 2576
rect 4488 2564 4494 2576
rect 4798 2564 4804 2576
rect 4488 2536 4804 2564
rect 4488 2524 4494 2536
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 4893 2567 4951 2573
rect 4893 2533 4905 2567
rect 4939 2564 4951 2567
rect 5994 2564 6000 2576
rect 4939 2536 6000 2564
rect 4939 2533 4951 2536
rect 4893 2527 4951 2533
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 6270 2524 6276 2576
rect 6328 2524 6334 2576
rect 6656 2564 6684 2595
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 8849 2635 8907 2641
rect 8849 2632 8861 2635
rect 8312 2604 8861 2632
rect 7374 2564 7380 2576
rect 6656 2536 7380 2564
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 8018 2564 8024 2576
rect 7760 2536 8024 2564
rect 4338 2456 4344 2508
rect 4396 2496 4402 2508
rect 4396 2468 5764 2496
rect 4396 2456 4402 2468
rect 4111 2400 4200 2428
rect 4525 2431 4583 2437
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4614 2428 4620 2440
rect 4571 2400 4620 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5166 2428 5172 2440
rect 5123 2400 5172 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 4430 2360 4436 2372
rect 3016 2332 4436 2360
rect 3016 2320 3022 2332
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 4246 2292 4252 2304
rect 2924 2264 4252 2292
rect 2924 2252 2930 2264
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 4522 2292 4528 2304
rect 4387 2264 4528 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 4816 2292 4844 2391
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5736 2437 5764 2468
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6288 2496 6316 2524
rect 5868 2468 6316 2496
rect 5868 2456 5874 2468
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 6696 2468 7144 2496
rect 6696 2456 6702 2468
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5767 2400 6009 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 5997 2397 6009 2400
rect 6043 2397 6055 2431
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 5997 2391 6055 2397
rect 6196 2400 6285 2428
rect 5276 2360 5304 2391
rect 5276 2332 5948 2360
rect 5810 2292 5816 2304
rect 4816 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 5920 2301 5948 2332
rect 6196 2301 6224 2400
rect 6273 2397 6285 2400
rect 6319 2397 6331 2431
rect 6822 2428 6828 2440
rect 6783 2400 6828 2428
rect 6273 2391 6331 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 7116 2437 7144 2468
rect 7760 2437 7788 2536
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 8312 2496 8340 2604
rect 8849 2601 8861 2604
rect 8895 2632 8907 2635
rect 9030 2632 9036 2644
rect 8895 2604 9036 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9674 2632 9680 2644
rect 9355 2604 9680 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 8386 2524 8392 2576
rect 8444 2564 8450 2576
rect 8444 2536 8800 2564
rect 8444 2524 8450 2536
rect 8036 2468 8340 2496
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 7469 2363 7527 2369
rect 7469 2329 7481 2363
rect 7515 2360 7527 2363
rect 7668 2360 7696 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8036 2437 8064 2468
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7892 2400 7941 2428
rect 7892 2388 7898 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8772 2437 8800 2536
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9766 2496 9772 2508
rect 9088 2468 9772 2496
rect 9088 2456 9094 2468
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8168 2400 8401 2428
rect 8168 2388 8174 2400
rect 8389 2397 8401 2400
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9582 2428 9588 2440
rect 9539 2400 9588 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 7515 2332 8432 2360
rect 7515 2329 7527 2332
rect 7469 2323 7527 2329
rect 8404 2304 8432 2332
rect 8588 2332 12572 2360
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2261 5963 2295
rect 5905 2255 5963 2261
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2261 6239 2295
rect 6181 2255 6239 2261
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 8076 2264 8217 2292
rect 8076 2252 8082 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 8588 2301 8616 2332
rect 8573 2295 8631 2301
rect 8573 2261 8585 2295
rect 8619 2261 8631 2295
rect 8573 2255 8631 2261
rect 8846 2252 8852 2304
rect 8904 2292 8910 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8904 2264 9229 2292
rect 8904 2252 8910 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 12544 2292 12572 2332
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 16850 2360 16856 2372
rect 13872 2332 16856 2360
rect 13872 2320 13878 2332
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 16758 2292 16764 2304
rect 12544 2264 16764 2292
rect 9217 2255 9275 2261
rect 16758 2252 16764 2264
rect 16816 2252 16822 2304
rect 3036 2202 9844 2224
rect 3036 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 5194 2202
rect 5246 2150 5258 2202
rect 5310 2150 5322 2202
rect 5374 2150 9844 2202
rect 3036 2128 9844 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 3605 2091 3663 2097
rect 3605 2088 3617 2091
rect 3292 2060 3617 2088
rect 3292 2048 3298 2060
rect 3605 2057 3617 2060
rect 3651 2057 3663 2091
rect 3878 2088 3884 2100
rect 3839 2060 3884 2088
rect 3605 2051 3663 2057
rect 3878 2048 3884 2060
rect 3936 2048 3942 2100
rect 4154 2088 4160 2100
rect 4115 2060 4160 2088
rect 4154 2048 4160 2060
rect 4212 2048 4218 2100
rect 4246 2048 4252 2100
rect 4304 2088 4310 2100
rect 4709 2091 4767 2097
rect 4709 2088 4721 2091
rect 4304 2060 4721 2088
rect 4304 2048 4310 2060
rect 4709 2057 4721 2060
rect 4755 2057 4767 2091
rect 9122 2088 9128 2100
rect 4709 2051 4767 2057
rect 5184 2060 9128 2088
rect 2682 1980 2688 2032
rect 2740 2020 2746 2032
rect 2740 1992 3832 2020
rect 2740 1980 2746 1992
rect 3510 1952 3516 1964
rect 3471 1924 3516 1952
rect 3510 1912 3516 1924
rect 3568 1912 3574 1964
rect 3804 1961 3832 1992
rect 3789 1955 3847 1961
rect 3789 1921 3801 1955
rect 3835 1921 3847 1955
rect 3789 1915 3847 1921
rect 4065 1955 4123 1961
rect 4065 1921 4077 1955
rect 4111 1921 4123 1955
rect 4065 1915 4123 1921
rect 4341 1955 4399 1961
rect 4341 1921 4353 1955
rect 4387 1921 4399 1955
rect 4341 1915 4399 1921
rect 4617 1955 4675 1961
rect 4617 1921 4629 1955
rect 4663 1952 4675 1955
rect 4706 1952 4712 1964
rect 4663 1924 4712 1952
rect 4663 1921 4675 1924
rect 4617 1915 4675 1921
rect 2774 1844 2780 1896
rect 2832 1884 2838 1896
rect 4080 1884 4108 1915
rect 2832 1856 4108 1884
rect 2832 1844 2838 1856
rect 4356 1816 4384 1915
rect 4706 1912 4712 1924
rect 4764 1912 4770 1964
rect 4798 1912 4804 1964
rect 4856 1952 4862 1964
rect 5184 1961 5212 2060
rect 9122 2048 9128 2060
rect 9180 2048 9186 2100
rect 7101 2023 7159 2029
rect 7101 1989 7113 2023
rect 7147 2020 7159 2023
rect 7466 2020 7472 2032
rect 7147 1992 7472 2020
rect 7147 1989 7159 1992
rect 7101 1983 7159 1989
rect 7466 1980 7472 1992
rect 7524 1980 7530 2032
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 8260 1992 8984 2020
rect 8260 1980 8266 1992
rect 4893 1955 4951 1961
rect 4893 1952 4905 1955
rect 4856 1924 4905 1952
rect 4856 1912 4862 1924
rect 4893 1921 4905 1924
rect 4939 1921 4951 1955
rect 4893 1915 4951 1921
rect 5169 1955 5227 1961
rect 5169 1921 5181 1955
rect 5215 1921 5227 1955
rect 7006 1952 7012 1964
rect 6967 1924 7012 1952
rect 5169 1915 5227 1921
rect 7006 1912 7012 1924
rect 7064 1912 7070 1964
rect 8113 1955 8171 1961
rect 8113 1921 8125 1955
rect 8159 1921 8171 1955
rect 8113 1915 8171 1921
rect 4522 1844 4528 1896
rect 4580 1884 4586 1896
rect 6086 1884 6092 1896
rect 4580 1856 6092 1884
rect 4580 1844 4586 1856
rect 6086 1844 6092 1856
rect 6144 1844 6150 1896
rect 7837 1887 7895 1893
rect 7837 1853 7849 1887
rect 7883 1884 7895 1887
rect 8128 1884 8156 1915
rect 8478 1912 8484 1964
rect 8536 1952 8542 1964
rect 8573 1955 8631 1961
rect 8573 1952 8585 1955
rect 8536 1924 8585 1952
rect 8536 1912 8542 1924
rect 8573 1921 8585 1924
rect 8619 1921 8631 1955
rect 8846 1952 8852 1964
rect 8807 1924 8852 1952
rect 8573 1915 8631 1921
rect 8846 1912 8852 1924
rect 8904 1912 8910 1964
rect 8956 1952 8984 1992
rect 9125 1955 9183 1961
rect 9125 1952 9137 1955
rect 8956 1924 9137 1952
rect 9125 1921 9137 1924
rect 9171 1921 9183 1955
rect 9125 1915 9183 1921
rect 9214 1912 9220 1964
rect 9272 1952 9278 1964
rect 9272 1924 9317 1952
rect 9272 1912 9278 1924
rect 16666 1884 16672 1896
rect 7883 1856 9076 1884
rect 7883 1853 7895 1856
rect 7837 1847 7895 1853
rect 2746 1788 4384 1816
rect 2498 1504 2504 1556
rect 2556 1544 2562 1556
rect 2746 1544 2774 1788
rect 4430 1776 4436 1828
rect 4488 1816 4494 1828
rect 4985 1819 5043 1825
rect 4488 1788 4533 1816
rect 4488 1776 4494 1788
rect 4985 1785 4997 1819
rect 5031 1816 5043 1819
rect 5626 1816 5632 1828
rect 5031 1788 5632 1816
rect 5031 1785 5043 1788
rect 4985 1779 5043 1785
rect 5626 1776 5632 1788
rect 5684 1776 5690 1828
rect 8294 1776 8300 1828
rect 8352 1816 8358 1828
rect 8389 1819 8447 1825
rect 8389 1816 8401 1819
rect 8352 1788 8401 1816
rect 8352 1776 8358 1788
rect 8389 1785 8401 1788
rect 8435 1785 8447 1819
rect 8389 1779 8447 1785
rect 8754 1776 8760 1828
rect 8812 1816 8818 1828
rect 8941 1819 8999 1825
rect 8941 1816 8953 1819
rect 8812 1788 8953 1816
rect 8812 1776 8818 1788
rect 8941 1785 8953 1788
rect 8987 1785 8999 1819
rect 8941 1779 8999 1785
rect 3329 1751 3387 1757
rect 3329 1748 3341 1751
rect 2556 1516 2774 1544
rect 2976 1720 3341 1748
rect 2976 1544 3004 1720
rect 3329 1717 3341 1720
rect 3375 1717 3387 1751
rect 7466 1748 7472 1760
rect 7427 1720 7472 1748
rect 3329 1711 3387 1717
rect 7466 1708 7472 1720
rect 7524 1708 7530 1760
rect 7929 1751 7987 1757
rect 7929 1717 7941 1751
rect 7975 1748 7987 1751
rect 8570 1748 8576 1760
rect 7975 1720 8576 1748
rect 7975 1717 7987 1720
rect 7929 1711 7987 1717
rect 8570 1708 8576 1720
rect 8628 1708 8634 1760
rect 8665 1751 8723 1757
rect 8665 1717 8677 1751
rect 8711 1748 8723 1751
rect 8846 1748 8852 1760
rect 8711 1720 8852 1748
rect 8711 1717 8723 1720
rect 8665 1711 8723 1717
rect 8846 1708 8852 1720
rect 8904 1708 8910 1760
rect 9048 1748 9076 1856
rect 12406 1856 16672 1884
rect 9401 1819 9459 1825
rect 9401 1785 9413 1819
rect 9447 1816 9459 1819
rect 12406 1816 12434 1856
rect 16666 1844 16672 1856
rect 16724 1844 16730 1896
rect 16574 1816 16580 1828
rect 9447 1788 12434 1816
rect 9447 1785 9459 1788
rect 9401 1779 9459 1785
rect 16546 1776 16580 1816
rect 16632 1776 16638 1828
rect 16546 1748 16574 1776
rect 9048 1720 16574 1748
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 6914 1544 6920 1556
rect 2976 1516 6920 1544
rect 2556 1504 2562 1516
rect 6914 1504 6920 1516
rect 6972 1504 6978 1556
rect 7006 1504 7012 1556
rect 7064 1544 7070 1556
rect 7653 1547 7711 1553
rect 7653 1544 7665 1547
rect 7064 1516 7665 1544
rect 7064 1504 7070 1516
rect 7653 1513 7665 1516
rect 7699 1513 7711 1547
rect 7653 1507 7711 1513
rect 8297 1547 8355 1553
rect 8297 1513 8309 1547
rect 8343 1544 8355 1547
rect 8662 1544 8668 1556
rect 8343 1516 8668 1544
rect 8343 1513 8355 1516
rect 8297 1507 8355 1513
rect 8662 1504 8668 1516
rect 8720 1504 8726 1556
rect 16942 1544 16948 1556
rect 16546 1516 16948 1544
rect 7466 1436 7472 1488
rect 7524 1476 7530 1488
rect 16546 1476 16574 1516
rect 16942 1504 16948 1516
rect 17000 1504 17006 1556
rect 7524 1448 16574 1476
rect 7524 1436 7530 1448
rect 7852 1349 7880 1448
rect 8386 1368 8392 1420
rect 8444 1408 8450 1420
rect 9122 1408 9128 1420
rect 8444 1380 8892 1408
rect 9083 1380 9128 1408
rect 8444 1368 8450 1380
rect 8864 1349 8892 1380
rect 9122 1368 9128 1380
rect 9180 1368 9186 1420
rect 3513 1343 3571 1349
rect 3513 1309 3525 1343
rect 3559 1309 3571 1343
rect 3513 1303 3571 1309
rect 7837 1343 7895 1349
rect 7837 1309 7849 1343
rect 7883 1309 7895 1343
rect 7837 1303 7895 1309
rect 8481 1343 8539 1349
rect 8481 1309 8493 1343
rect 8527 1309 8539 1343
rect 8481 1303 8539 1309
rect 8849 1343 8907 1349
rect 8849 1309 8861 1343
rect 8895 1340 8907 1343
rect 8938 1340 8944 1352
rect 8895 1312 8944 1340
rect 8895 1309 8907 1312
rect 8849 1303 8907 1309
rect 3528 1272 3556 1303
rect 7926 1272 7932 1284
rect 3528 1244 7932 1272
rect 7926 1232 7932 1244
rect 7984 1232 7990 1284
rect 8496 1272 8524 1303
rect 8938 1300 8944 1312
rect 8996 1300 9002 1352
rect 9490 1340 9496 1352
rect 9451 1312 9496 1340
rect 9490 1300 9496 1312
rect 9548 1300 9554 1352
rect 16574 1340 16580 1352
rect 16546 1300 16580 1340
rect 16632 1300 16638 1352
rect 16546 1272 16574 1300
rect 8496 1244 16574 1272
rect 3326 1204 3332 1216
rect 3287 1176 3332 1204
rect 3326 1164 3332 1176
rect 3384 1164 3390 1216
rect 9309 1207 9367 1213
rect 9309 1173 9321 1207
rect 9355 1204 9367 1207
rect 9398 1204 9404 1216
rect 9355 1176 9404 1204
rect 9355 1173 9367 1176
rect 9309 1167 9367 1173
rect 9398 1164 9404 1176
rect 9456 1164 9462 1216
rect 3036 1114 9844 1136
rect 3036 1062 5066 1114
rect 5118 1062 5130 1114
rect 5182 1062 5194 1114
rect 5246 1062 5258 1114
rect 5310 1062 5322 1114
rect 5374 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 2412 12180 2464 12232
rect 9496 12180 9548 12232
rect 4344 12112 4396 12164
rect 9404 12112 9456 12164
rect 5816 12044 5868 12096
rect 9312 12044 9364 12096
rect 3056 11976 3108 12028
rect 8760 11976 8812 12028
rect 4804 11908 4856 11960
rect 8668 11908 8720 11960
rect 2780 11840 2832 11892
rect 3792 11840 3844 11892
rect 4988 11840 5040 11892
rect 8392 11840 8444 11892
rect 1492 11772 1544 11824
rect 6644 11772 6696 11824
rect 7012 11772 7064 11824
rect 13544 11840 13596 11892
rect 2412 11704 2464 11756
rect 5816 11704 5868 11756
rect 5908 11704 5960 11756
rect 13820 11704 13872 11756
rect 1308 11500 1360 11552
rect 6828 11636 6880 11688
rect 2964 11568 3016 11620
rect 8116 11568 8168 11620
rect 3240 11500 3292 11552
rect 6184 11500 6236 11552
rect 6736 11500 6788 11552
rect 8300 11500 8352 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 1308 11339 1360 11348
rect 1308 11305 1317 11339
rect 1317 11305 1351 11339
rect 1351 11305 1360 11339
rect 1308 11296 1360 11305
rect 3240 11296 3292 11348
rect 2228 11228 2280 11280
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 5908 11339 5960 11348
rect 5908 11305 5917 11339
rect 5917 11305 5951 11339
rect 5951 11305 5960 11339
rect 5908 11296 5960 11305
rect 6092 11296 6144 11348
rect 6644 11339 6696 11348
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 2688 11160 2740 11212
rect 4344 11228 4396 11280
rect 6644 11305 6653 11339
rect 6653 11305 6687 11339
rect 6687 11305 6696 11339
rect 6644 11296 6696 11305
rect 7012 11339 7064 11348
rect 7012 11305 7021 11339
rect 7021 11305 7055 11339
rect 7055 11305 7064 11339
rect 7012 11296 7064 11305
rect 8116 11339 8168 11348
rect 8116 11305 8125 11339
rect 8125 11305 8159 11339
rect 8159 11305 8168 11339
rect 8116 11296 8168 11305
rect 2320 11092 2372 11144
rect 2412 11092 2464 11144
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3424 11092 3476 11144
rect 2320 10999 2372 11008
rect 2320 10965 2329 10999
rect 2329 10965 2363 10999
rect 2363 10965 2372 10999
rect 2320 10956 2372 10965
rect 3056 11024 3108 11076
rect 3516 11024 3568 11076
rect 3976 11067 4028 11076
rect 3976 11033 3985 11067
rect 3985 11033 4019 11067
rect 4019 11033 4028 11067
rect 3976 11024 4028 11033
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 4712 11092 4764 11144
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 7380 11160 7432 11212
rect 8852 11228 8904 11280
rect 9128 11228 9180 11280
rect 13636 11160 13688 11212
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6000 11092 6052 11144
rect 7288 11135 7340 11144
rect 6736 11024 6788 11076
rect 4068 10956 4120 11008
rect 4528 10956 4580 11008
rect 4804 10999 4856 11008
rect 4804 10965 4813 10999
rect 4813 10965 4847 10999
rect 4847 10965 4856 10999
rect 4804 10956 4856 10965
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 8576 11092 8628 11144
rect 9036 11101 9045 11120
rect 9045 11101 9079 11120
rect 9079 11101 9088 11120
rect 9036 11068 9088 11101
rect 8300 10956 8352 11008
rect 10416 11024 10468 11076
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5194 10854 5246 10906
rect 5258 10854 5310 10906
rect 5322 10854 5374 10906
rect 1400 10752 1452 10804
rect 2780 10752 2832 10804
rect 2872 10752 2924 10804
rect 1952 10684 2004 10736
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2504 10684 2556 10736
rect 4804 10684 4856 10736
rect 2136 10616 2188 10625
rect 3516 10616 3568 10668
rect 3884 10616 3936 10668
rect 6828 10684 6880 10736
rect 2504 10480 2556 10532
rect 2688 10480 2740 10532
rect 3148 10480 3200 10532
rect 4712 10548 4764 10600
rect 6000 10616 6052 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 8760 10752 8812 10804
rect 8208 10684 8260 10736
rect 5724 10548 5776 10600
rect 6092 10548 6144 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 1676 10412 1728 10464
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 4068 10412 4120 10464
rect 5080 10480 5132 10532
rect 7472 10480 7524 10532
rect 9588 10616 9640 10668
rect 5356 10412 5408 10464
rect 8116 10412 8168 10464
rect 9220 10480 9272 10532
rect 8760 10412 8812 10464
rect 9036 10412 9088 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 1584 10208 1636 10260
rect 2964 10140 3016 10192
rect 2320 10072 2372 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 4712 10072 4764 10124
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 6092 10208 6144 10260
rect 6828 10208 6880 10260
rect 7012 10208 7064 10260
rect 7472 10208 7524 10260
rect 7380 10140 7432 10192
rect 8208 10208 8260 10260
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 8576 10208 8628 10260
rect 7932 10140 7984 10192
rect 7748 10004 7800 10056
rect 8576 10004 8628 10056
rect 13820 10004 13872 10056
rect 22284 10004 22336 10056
rect 2688 9936 2740 9988
rect 3240 9936 3292 9988
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2320 9868 2372 9920
rect 2596 9868 2648 9920
rect 5816 9936 5868 9988
rect 6828 9936 6880 9988
rect 7656 9936 7708 9988
rect 4712 9868 4764 9920
rect 6184 9868 6236 9920
rect 8208 9868 8260 9920
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5194 9766 5246 9818
rect 5258 9766 5310 9818
rect 5322 9766 5374 9818
rect 2136 9664 2188 9716
rect 2320 9664 2372 9716
rect 6184 9664 6236 9716
rect 6552 9664 6604 9716
rect 7196 9664 7248 9716
rect 7656 9664 7708 9716
rect 1860 9596 1912 9648
rect 3332 9596 3384 9648
rect 5540 9639 5592 9648
rect 5540 9605 5549 9639
rect 5549 9605 5583 9639
rect 5583 9605 5592 9639
rect 5540 9596 5592 9605
rect 6092 9596 6144 9648
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 4344 9528 4396 9580
rect 5264 9528 5316 9580
rect 5724 9528 5776 9580
rect 6368 9596 6420 9648
rect 6920 9571 6972 9580
rect 2320 9460 2372 9512
rect 2964 9460 3016 9512
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 9312 9596 9364 9648
rect 7656 9528 7708 9580
rect 9496 9528 9548 9580
rect 1860 9324 1912 9376
rect 1952 9324 2004 9376
rect 2412 9324 2464 9376
rect 6736 9460 6788 9512
rect 8208 9460 8260 9512
rect 5356 9324 5408 9376
rect 5724 9392 5776 9444
rect 5908 9324 5960 9376
rect 7104 9324 7156 9376
rect 8300 9324 8352 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 1216 9120 1268 9172
rect 1032 8916 1084 8968
rect 2136 9120 2188 9172
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 1952 9052 2004 9104
rect 1768 8916 1820 8968
rect 3424 9163 3476 9172
rect 2504 8916 2556 8968
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 3608 9120 3660 9172
rect 4068 9120 4120 9172
rect 4896 9120 4948 9172
rect 5356 9120 5408 9172
rect 3332 9052 3384 9104
rect 3792 9052 3844 9104
rect 4160 9052 4212 9104
rect 8208 9120 8260 9172
rect 8760 9052 8812 9104
rect 9312 9052 9364 9104
rect 3976 8984 4028 9036
rect 8576 8984 8628 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4068 8916 4120 8968
rect 5264 8916 5316 8968
rect 6736 8916 6788 8968
rect 7288 8916 7340 8968
rect 8760 8959 8812 8968
rect 2228 8848 2280 8900
rect 1124 8780 1176 8832
rect 1492 8780 1544 8832
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 3332 8848 3384 8900
rect 4344 8848 4396 8900
rect 4804 8848 4856 8900
rect 5908 8848 5960 8900
rect 7472 8780 7524 8832
rect 7656 8848 7708 8900
rect 8208 8848 8260 8900
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 9680 8848 9732 8900
rect 8392 8780 8444 8832
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5194 8678 5246 8730
rect 5258 8678 5310 8730
rect 5322 8678 5374 8730
rect 1768 8576 1820 8628
rect 1492 8508 1544 8560
rect 2504 8508 2556 8560
rect 4436 8508 4488 8560
rect 1952 8440 2004 8492
rect 2228 8440 2280 8492
rect 1768 8372 1820 8424
rect 2044 8372 2096 8424
rect 1676 8304 1728 8356
rect 2964 8372 3016 8424
rect 1308 8236 1360 8288
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 4896 8372 4948 8424
rect 5080 8372 5132 8424
rect 6736 8508 6788 8560
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 8484 8576 8536 8628
rect 8668 8508 8720 8560
rect 9404 8440 9456 8492
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 6000 8372 6052 8424
rect 8208 8372 8260 8424
rect 4068 8279 4120 8288
rect 4068 8245 4077 8279
rect 4077 8245 4111 8279
rect 4111 8245 4120 8279
rect 4068 8236 4120 8245
rect 5632 8236 5684 8288
rect 6000 8236 6052 8288
rect 7012 8236 7064 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 3240 8032 3292 8084
rect 4436 8032 4488 8084
rect 4620 8032 4672 8084
rect 8760 8032 8812 8084
rect 5080 7964 5132 8016
rect 8576 8007 8628 8016
rect 8576 7973 8585 8007
rect 8585 7973 8619 8007
rect 8619 7973 8628 8007
rect 8576 7964 8628 7973
rect 1584 7896 1636 7948
rect 6000 7896 6052 7948
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 4068 7828 4120 7880
rect 4804 7828 4856 7880
rect 7012 7871 7064 7880
rect 1860 7760 1912 7812
rect 940 7692 992 7744
rect 1584 7692 1636 7744
rect 3240 7760 3292 7812
rect 3700 7760 3752 7812
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 7472 7828 7524 7880
rect 8668 7828 8720 7880
rect 8392 7803 8444 7812
rect 2596 7692 2648 7744
rect 2688 7692 2740 7744
rect 4436 7692 4488 7744
rect 4620 7692 4672 7744
rect 7380 7692 7432 7744
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 8300 7692 8352 7744
rect 8760 7692 8812 7744
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5194 7590 5246 7642
rect 5258 7590 5310 7642
rect 5322 7590 5374 7642
rect 8392 7488 8444 7540
rect 2228 7420 2280 7472
rect 3332 7420 3384 7472
rect 4252 7420 4304 7472
rect 1308 7284 1360 7336
rect 4528 7352 4580 7404
rect 5908 7352 5960 7404
rect 6828 7420 6880 7472
rect 1676 7216 1728 7268
rect 1952 7216 2004 7268
rect 2688 7216 2740 7268
rect 6184 7284 6236 7336
rect 6736 7284 6788 7336
rect 7012 7284 7064 7336
rect 8392 7284 8444 7336
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 6460 7216 6512 7268
rect 7196 7216 7248 7268
rect 4620 7148 4672 7200
rect 4988 7148 5040 7200
rect 6644 7148 6696 7200
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 9404 7148 9456 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 1952 6987 2004 6996
rect 1952 6953 1982 6987
rect 1982 6953 2004 6987
rect 1952 6944 2004 6953
rect 2964 6944 3016 6996
rect 3608 6944 3660 6996
rect 5908 6987 5960 6996
rect 5908 6953 5917 6987
rect 5917 6953 5951 6987
rect 5951 6953 5960 6987
rect 5908 6944 5960 6953
rect 6184 6987 6236 6996
rect 6184 6953 6193 6987
rect 6193 6953 6227 6987
rect 6227 6953 6236 6987
rect 6184 6944 6236 6953
rect 7472 6944 7524 6996
rect 8300 6944 8352 6996
rect 7840 6876 7892 6928
rect 8116 6876 8168 6928
rect 8576 6876 8628 6928
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 1952 6808 2004 6860
rect 4344 6808 4396 6860
rect 4528 6808 4580 6860
rect 6920 6808 6972 6860
rect 9220 6808 9272 6860
rect 1492 6740 1544 6792
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 3240 6672 3292 6724
rect 1216 6604 1268 6656
rect 2228 6604 2280 6656
rect 6552 6672 6604 6724
rect 7104 6672 7156 6724
rect 7840 6672 7892 6724
rect 8484 6672 8536 6724
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 8668 6604 8720 6656
rect 8944 6604 8996 6656
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5194 6502 5246 6554
rect 5258 6502 5310 6554
rect 5322 6502 5374 6554
rect 1400 6400 1452 6452
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 1860 6400 1912 6452
rect 1492 6264 1544 6316
rect 1952 6264 2004 6316
rect 3700 6400 3752 6452
rect 3976 6400 4028 6452
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 2964 6332 3016 6384
rect 4804 6332 4856 6384
rect 3700 6264 3752 6316
rect 3976 6264 4028 6316
rect 4436 6264 4488 6316
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5540 6264 5592 6316
rect 7196 6400 7248 6452
rect 8116 6400 8168 6452
rect 8944 6400 8996 6452
rect 6736 6264 6788 6316
rect 8852 6264 8904 6316
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 9496 6264 9548 6273
rect 1676 6196 1728 6248
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 3424 6196 3476 6248
rect 7288 6239 7340 6248
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 2136 6060 2188 6112
rect 5724 6128 5776 6180
rect 4620 6060 4672 6112
rect 6184 6060 6236 6112
rect 9036 6060 9088 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 1860 5856 1912 5908
rect 3608 5856 3660 5908
rect 3700 5899 3752 5908
rect 3700 5865 3709 5899
rect 3709 5865 3743 5899
rect 3743 5865 3752 5899
rect 3700 5856 3752 5865
rect 1308 5788 1360 5840
rect 2964 5831 3016 5840
rect 2964 5797 2973 5831
rect 2973 5797 3007 5831
rect 3007 5797 3016 5831
rect 2964 5788 3016 5797
rect 1584 5652 1636 5704
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 1216 5584 1268 5636
rect 2136 5652 2188 5704
rect 2964 5652 3016 5704
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 2228 5516 2280 5568
rect 3424 5720 3476 5772
rect 3424 5628 3476 5680
rect 3700 5652 3752 5704
rect 6000 5856 6052 5908
rect 4160 5720 4212 5772
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 9496 5856 9548 5908
rect 8208 5788 8260 5840
rect 6828 5763 6880 5772
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 5540 5652 5592 5704
rect 6092 5652 6144 5704
rect 6552 5652 6604 5704
rect 6460 5584 6512 5636
rect 6828 5729 6837 5763
rect 6837 5729 6871 5763
rect 6871 5729 6880 5763
rect 6828 5720 6880 5729
rect 8300 5720 8352 5772
rect 13820 5720 13872 5772
rect 16948 5720 17000 5772
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 7564 5584 7616 5636
rect 6552 5516 6604 5568
rect 6828 5516 6880 5568
rect 7196 5516 7248 5568
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5194 5414 5246 5466
rect 5258 5414 5310 5466
rect 5322 5414 5374 5466
rect 4896 5312 4948 5364
rect 8760 5312 8812 5364
rect 9312 5312 9364 5364
rect 1124 5244 1176 5296
rect 2688 5244 2740 5296
rect 5540 5287 5592 5296
rect 5540 5253 5549 5287
rect 5549 5253 5583 5287
rect 5583 5253 5592 5287
rect 5540 5244 5592 5253
rect 7472 5244 7524 5296
rect 2412 5176 2464 5228
rect 2044 5108 2096 5160
rect 2780 5108 2832 5160
rect 4896 5176 4948 5228
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 6000 5176 6052 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 7104 5176 7156 5228
rect 4620 5108 4672 5160
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 8392 5176 8444 5228
rect 7196 5040 7248 5092
rect 9404 5108 9456 5160
rect 13820 5040 13872 5092
rect 4252 4972 4304 5024
rect 5540 4972 5592 5024
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 3608 4768 3660 4820
rect 4896 4768 4948 4820
rect 7288 4768 7340 4820
rect 1032 4564 1084 4616
rect 3148 4564 3200 4616
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 5356 4700 5408 4752
rect 4620 4632 4672 4684
rect 5632 4632 5684 4684
rect 6920 4632 6972 4684
rect 7840 4632 7892 4684
rect 8024 4632 8076 4684
rect 2872 4496 2924 4548
rect 4252 4564 4304 4616
rect 5080 4564 5132 4616
rect 6000 4564 6052 4616
rect 6552 4539 6604 4548
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 4528 4428 4580 4480
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 4988 4428 5040 4480
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 6552 4505 6561 4539
rect 6561 4505 6595 4539
rect 6595 4505 6604 4539
rect 6552 4496 6604 4505
rect 7288 4428 7340 4480
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5194 4326 5246 4378
rect 5258 4326 5310 4378
rect 5322 4326 5374 4378
rect 4252 4224 4304 4276
rect 4712 4224 4764 4276
rect 6736 4267 6788 4276
rect 4436 4156 4488 4208
rect 6736 4233 6745 4267
rect 6745 4233 6779 4267
rect 6779 4233 6788 4267
rect 6736 4224 6788 4233
rect 7472 4224 7524 4276
rect 9772 4224 9824 4276
rect 5264 4156 5316 4208
rect 8852 4156 8904 4208
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 5448 4131 5500 4140
rect 3608 4088 3660 4097
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 6552 4088 6604 4140
rect 6736 4088 6788 4140
rect 7472 4088 7524 4140
rect 8576 4088 8628 4140
rect 8944 4088 8996 4140
rect 4620 4020 4672 4072
rect 8668 4020 8720 4072
rect 9588 4020 9640 4072
rect 7748 3952 7800 4004
rect 7840 3952 7892 4004
rect 13820 3952 13872 4004
rect 5172 3884 5224 3936
rect 6920 3884 6972 3936
rect 9220 3884 9272 3936
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 3424 3680 3476 3732
rect 4436 3680 4488 3732
rect 4712 3723 4764 3732
rect 4712 3689 4721 3723
rect 4721 3689 4755 3723
rect 4755 3689 4764 3723
rect 4712 3680 4764 3689
rect 3608 3612 3660 3664
rect 4620 3612 4672 3664
rect 6000 3680 6052 3732
rect 5632 3612 5684 3664
rect 8208 3680 8260 3732
rect 9220 3680 9272 3732
rect 3240 3544 3292 3596
rect 3700 3476 3752 3528
rect 4252 3544 4304 3596
rect 4436 3544 4488 3596
rect 4804 3544 4856 3596
rect 4344 3476 4396 3528
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 5448 3544 5500 3596
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 3700 3340 3752 3392
rect 4068 3340 4120 3392
rect 5540 3408 5592 3460
rect 5724 3476 5776 3528
rect 6092 3544 6144 3596
rect 6920 3587 6972 3596
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 13728 3612 13780 3664
rect 9864 3544 9916 3596
rect 16580 3544 16632 3596
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6552 3519 6604 3528
rect 6000 3476 6052 3485
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 8576 3476 8628 3528
rect 8760 3408 8812 3460
rect 6184 3340 6236 3392
rect 6828 3340 6880 3392
rect 7380 3340 7432 3392
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9496 3340 9548 3392
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5194 3238 5246 3290
rect 5258 3238 5310 3290
rect 5322 3238 5374 3290
rect 13820 3272 13872 3324
rect 16764 3272 16816 3324
rect 3700 3136 3752 3188
rect 3792 3136 3844 3188
rect 4068 3136 4120 3188
rect 3056 3068 3108 3120
rect 3976 3000 4028 3052
rect 4988 3068 5040 3120
rect 6000 3068 6052 3120
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 4528 3000 4580 3052
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 6736 3000 6788 3052
rect 7472 3068 7524 3120
rect 8576 3136 8628 3188
rect 13452 3136 13504 3188
rect 13636 3136 13688 3188
rect 16856 3136 16908 3188
rect 8208 3000 8260 3052
rect 8576 3000 8628 3052
rect 8944 3000 8996 3052
rect 5172 2932 5224 2984
rect 8116 2932 8168 2984
rect 6460 2864 6512 2916
rect 9772 2932 9824 2984
rect 13820 2864 13872 2916
rect 22192 2864 22244 2916
rect 8208 2796 8260 2848
rect 8668 2839 8720 2848
rect 8668 2805 8677 2839
rect 8677 2805 8711 2839
rect 8711 2805 8720 2839
rect 8668 2796 8720 2805
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 3516 2592 3568 2644
rect 3976 2592 4028 2644
rect 4068 2524 4120 2576
rect 4528 2592 4580 2644
rect 5172 2592 5224 2644
rect 5816 2592 5868 2644
rect 6552 2592 6604 2644
rect 4436 2524 4488 2576
rect 4804 2524 4856 2576
rect 6000 2524 6052 2576
rect 6276 2524 6328 2576
rect 7104 2592 7156 2644
rect 7380 2524 7432 2576
rect 4344 2456 4396 2508
rect 4620 2388 4672 2440
rect 2964 2320 3016 2372
rect 4436 2320 4488 2372
rect 2872 2252 2924 2304
rect 4252 2252 4304 2304
rect 4528 2252 4580 2304
rect 5172 2388 5224 2440
rect 5816 2456 5868 2508
rect 6644 2456 6696 2508
rect 5816 2252 5868 2304
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 8024 2524 8076 2576
rect 9036 2592 9088 2644
rect 9680 2592 9732 2644
rect 8392 2524 8444 2576
rect 7840 2388 7892 2440
rect 8116 2388 8168 2440
rect 9036 2456 9088 2508
rect 9772 2456 9824 2508
rect 9588 2388 9640 2440
rect 8024 2252 8076 2304
rect 8392 2252 8444 2304
rect 8852 2252 8904 2304
rect 13820 2320 13872 2372
rect 16856 2320 16908 2372
rect 16764 2252 16816 2304
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 5194 2150 5246 2202
rect 5258 2150 5310 2202
rect 5322 2150 5374 2202
rect 3240 2048 3292 2100
rect 3884 2091 3936 2100
rect 3884 2057 3893 2091
rect 3893 2057 3927 2091
rect 3927 2057 3936 2091
rect 3884 2048 3936 2057
rect 4160 2091 4212 2100
rect 4160 2057 4169 2091
rect 4169 2057 4203 2091
rect 4203 2057 4212 2091
rect 4160 2048 4212 2057
rect 4252 2048 4304 2100
rect 2688 1980 2740 2032
rect 3516 1955 3568 1964
rect 3516 1921 3525 1955
rect 3525 1921 3559 1955
rect 3559 1921 3568 1955
rect 3516 1912 3568 1921
rect 2780 1844 2832 1896
rect 4712 1912 4764 1964
rect 4804 1912 4856 1964
rect 9128 2048 9180 2100
rect 7472 1980 7524 2032
rect 8208 1980 8260 2032
rect 7012 1955 7064 1964
rect 7012 1921 7021 1955
rect 7021 1921 7055 1955
rect 7055 1921 7064 1955
rect 7012 1912 7064 1921
rect 4528 1844 4580 1896
rect 6092 1844 6144 1896
rect 8484 1912 8536 1964
rect 8852 1955 8904 1964
rect 8852 1921 8861 1955
rect 8861 1921 8895 1955
rect 8895 1921 8904 1955
rect 8852 1912 8904 1921
rect 9220 1955 9272 1964
rect 9220 1921 9229 1955
rect 9229 1921 9263 1955
rect 9263 1921 9272 1955
rect 9220 1912 9272 1921
rect 2504 1504 2556 1556
rect 4436 1819 4488 1828
rect 4436 1785 4445 1819
rect 4445 1785 4479 1819
rect 4479 1785 4488 1819
rect 4436 1776 4488 1785
rect 5632 1776 5684 1828
rect 8300 1776 8352 1828
rect 8760 1776 8812 1828
rect 7472 1751 7524 1760
rect 7472 1717 7481 1751
rect 7481 1717 7515 1751
rect 7515 1717 7524 1751
rect 7472 1708 7524 1717
rect 8576 1708 8628 1760
rect 8852 1708 8904 1760
rect 16672 1844 16724 1896
rect 16580 1776 16632 1828
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 6920 1504 6972 1556
rect 7012 1504 7064 1556
rect 8668 1504 8720 1556
rect 7472 1436 7524 1488
rect 16948 1504 17000 1556
rect 8392 1368 8444 1420
rect 9128 1411 9180 1420
rect 9128 1377 9137 1411
rect 9137 1377 9171 1411
rect 9171 1377 9180 1411
rect 9128 1368 9180 1377
rect 8944 1343 8996 1352
rect 7932 1232 7984 1284
rect 8944 1309 8953 1343
rect 8953 1309 8987 1343
rect 8987 1309 8996 1343
rect 8944 1300 8996 1309
rect 9496 1343 9548 1352
rect 9496 1309 9505 1343
rect 9505 1309 9539 1343
rect 9539 1309 9548 1343
rect 9496 1300 9548 1309
rect 16580 1300 16632 1352
rect 3332 1207 3384 1216
rect 3332 1173 3341 1207
rect 3341 1173 3375 1207
rect 3375 1173 3384 1207
rect 3332 1164 3384 1173
rect 9404 1164 9456 1216
rect 5066 1062 5118 1114
rect 5130 1062 5182 1114
rect 5194 1062 5246 1114
rect 5258 1062 5310 1114
rect 5322 1062 5374 1114
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 1858 12200 1914 13000
rect 2056 12294 2268 12322
rect 952 7750 980 12200
rect 1308 11552 1360 11558
rect 1308 11494 1360 11500
rect 1320 11354 1348 11494
rect 1308 11348 1360 11354
rect 1308 11290 1360 11296
rect 1412 10962 1440 12200
rect 1492 11824 1544 11830
rect 1492 11766 1544 11772
rect 1504 11150 1532 11766
rect 1872 11234 1900 12200
rect 1780 11206 1900 11234
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1412 10934 1532 10962
rect 1398 10840 1454 10849
rect 1398 10775 1400 10784
rect 1452 10775 1454 10784
rect 1400 10746 1452 10752
rect 1214 10704 1270 10713
rect 1214 10639 1270 10648
rect 1228 9178 1256 10639
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1306 9480 1362 9489
rect 1306 9415 1362 9424
rect 1216 9172 1268 9178
rect 1216 9114 1268 9120
rect 1032 8968 1084 8974
rect 1032 8910 1084 8916
rect 940 7744 992 7750
rect 940 7686 992 7692
rect 1044 4622 1072 8910
rect 1124 8832 1176 8838
rect 1124 8774 1176 8780
rect 1136 5302 1164 8774
rect 1320 8378 1348 9415
rect 1228 8350 1348 8378
rect 1228 6746 1256 8350
rect 1308 8288 1360 8294
rect 1308 8230 1360 8236
rect 1320 7342 1348 8230
rect 1308 7336 1360 7342
rect 1308 7278 1360 7284
rect 1228 6718 1348 6746
rect 1216 6656 1268 6662
rect 1216 6598 1268 6604
rect 1228 5642 1256 6598
rect 1320 5846 1348 6718
rect 1412 6458 1440 9998
rect 1504 8838 1532 10934
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1596 10266 1624 10406
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1688 10169 1716 10406
rect 1674 10160 1730 10169
rect 1674 10095 1730 10104
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1492 8560 1544 8566
rect 1492 8502 1544 8508
rect 1504 6798 1532 8502
rect 1596 7954 1624 9862
rect 1688 8362 1716 9998
rect 1780 8974 1808 11206
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1872 9654 1900 11086
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1964 9382 1992 10678
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8634 1808 8774
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1688 7886 1716 8298
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1504 6322 1532 6734
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1308 5840 1360 5846
rect 1308 5782 1360 5788
rect 1596 5710 1624 7686
rect 1688 7274 1716 7822
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1688 6866 1716 7210
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1688 6254 1716 6802
rect 1780 6458 1808 8366
rect 1872 7818 1900 9318
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 2056 9058 2084 12294
rect 2240 12152 2268 12294
rect 2318 12200 2374 13000
rect 2412 12232 2464 12238
rect 2332 12152 2360 12200
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6104 12294 6316 12322
rect 2412 12174 2464 12180
rect 2240 12124 2360 12152
rect 2424 12016 2452 12174
rect 2332 11988 2452 12016
rect 2228 11280 2280 11286
rect 2228 11222 2280 11228
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 9722 2176 10610
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2136 9172 2188 9178
rect 2240 9160 2268 11222
rect 2332 11150 2360 11988
rect 2792 11898 2820 12200
rect 3056 12028 3108 12034
rect 3056 11970 3108 11976
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2424 11150 2452 11698
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10130 2360 10950
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2516 10538 2544 10678
rect 2700 10538 2728 11154
rect 2872 11144 2924 11150
rect 2976 11132 3004 11562
rect 2924 11104 3004 11132
rect 2872 11086 2924 11092
rect 3068 11082 3096 11970
rect 3252 11642 3280 12200
rect 3252 11614 3372 11642
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11354 3280 11494
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2870 10840 2926 10849
rect 2780 10804 2832 10810
rect 2870 10775 2872 10784
rect 2780 10746 2832 10752
rect 2924 10775 2926 10784
rect 2872 10746 2924 10752
rect 2792 10577 2820 10746
rect 2778 10568 2834 10577
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2688 10532 2740 10538
rect 2778 10503 2834 10512
rect 3148 10532 3200 10538
rect 2688 10474 2740 10480
rect 3148 10474 3200 10480
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2964 10192 3016 10198
rect 2594 10160 2650 10169
rect 2320 10124 2372 10130
rect 2594 10095 2650 10104
rect 2778 10160 2834 10169
rect 2964 10134 3016 10140
rect 2778 10095 2834 10104
rect 2320 10066 2372 10072
rect 2608 9926 2636 10095
rect 2688 9988 2740 9994
rect 2792 9976 2820 10095
rect 2740 9948 2820 9976
rect 2688 9930 2740 9936
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2332 9722 2360 9862
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2332 9178 2360 9454
rect 2424 9382 2452 9522
rect 2976 9518 3004 10134
rect 3068 9586 3096 10406
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2188 9132 2268 9160
rect 2320 9172 2372 9178
rect 2136 9114 2188 9120
rect 2320 9114 2372 9120
rect 1964 8616 1992 9046
rect 2056 9030 2176 9058
rect 1964 8588 2084 8616
rect 2056 8537 2084 8588
rect 2042 8528 2098 8537
rect 1952 8492 2004 8498
rect 2042 8463 2098 8472
rect 1952 8434 2004 8440
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 6458 1900 7754
rect 1964 7274 1992 8434
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2148 8378 2176 9030
rect 2504 8968 2556 8974
rect 2410 8936 2466 8945
rect 2228 8900 2280 8906
rect 2504 8910 2556 8916
rect 2410 8871 2466 8880
rect 2228 8842 2280 8848
rect 2240 8498 2268 8842
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 1964 7002 1992 7210
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1858 6352 1914 6361
rect 1964 6322 1992 6802
rect 1858 6287 1914 6296
rect 1952 6316 2004 6322
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1872 5914 1900 6287
rect 1952 6258 2004 6264
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1950 5808 2006 5817
rect 1950 5743 2006 5752
rect 1964 5710 1992 5743
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1216 5636 1268 5642
rect 1216 5578 1268 5584
rect 1124 5296 1176 5302
rect 1124 5238 1176 5244
rect 2056 5166 2084 8366
rect 2148 8350 2360 8378
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2240 7478 2268 8230
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5710 2176 6054
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2240 5574 2268 6598
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2332 5114 2360 8350
rect 2424 6984 2452 8871
rect 2516 8566 2544 8910
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2976 8430 3004 9454
rect 3054 9072 3110 9081
rect 3054 9007 3110 9016
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2594 7984 2650 7993
rect 2594 7919 2650 7928
rect 2608 7750 2636 7919
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2700 7274 2728 7686
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2964 6996 3016 7002
rect 2424 6956 2544 6984
rect 2412 6248 2464 6254
rect 2516 6225 2544 6956
rect 2964 6938 3016 6944
rect 2976 6390 3004 6938
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3068 6236 3096 9007
rect 3160 8974 3188 10474
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 10169 3280 10406
rect 3238 10160 3294 10169
rect 3238 10095 3294 10104
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 3252 9081 3280 9930
rect 3344 9761 3372 11614
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3344 9110 3372 9590
rect 3436 9178 3464 11086
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3528 10674 3556 11018
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3332 9104 3384 9110
rect 3238 9072 3294 9081
rect 3528 9058 3556 10610
rect 3606 10160 3662 10169
rect 3606 10095 3662 10104
rect 3620 9178 3648 10095
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3332 9046 3384 9052
rect 3238 9007 3294 9016
rect 3436 9030 3556 9058
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3146 8392 3202 8401
rect 3146 8327 3202 8336
rect 2412 6190 2464 6196
rect 2502 6216 2558 6225
rect 2424 5234 2452 6190
rect 2502 6151 2558 6160
rect 2976 6208 3096 6236
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 2976 5846 3004 6208
rect 3054 5944 3110 5953
rect 3054 5879 3110 5888
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 3068 5710 3096 5879
rect 3160 5794 3188 8327
rect 3252 8090 3280 8910
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3252 6730 3280 7754
rect 3344 7478 3372 8842
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3436 7290 3464 9030
rect 3712 8242 3740 12200
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3804 9217 3832 11834
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3790 9208 3846 9217
rect 3790 9143 3846 9152
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3344 7262 3464 7290
rect 3528 8214 3740 8242
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3252 6225 3280 6666
rect 3238 6216 3294 6225
rect 3238 6151 3294 6160
rect 3160 5766 3280 5794
rect 2964 5704 3016 5710
rect 2962 5672 2964 5681
rect 3056 5704 3108 5710
rect 3016 5672 3018 5681
rect 3056 5646 3108 5652
rect 2962 5607 3018 5616
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2332 5086 2544 5114
rect 1032 4616 1084 4622
rect 1032 4558 1084 4564
rect 2516 1562 2544 5086
rect 2700 2038 2728 5238
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2688 2032 2740 2038
rect 2688 1974 2740 1980
rect 2792 1902 2820 5102
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2884 2310 2912 4490
rect 2976 2378 3004 5607
rect 3068 3126 3096 5646
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3160 2417 3188 4558
rect 3252 3602 3280 5766
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3344 2774 3372 7262
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3436 5778 3464 6190
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3424 5681 3476 5686
rect 3422 5680 3478 5681
rect 3422 5672 3424 5680
rect 3476 5672 3478 5680
rect 3422 5607 3478 5616
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3436 3738 3464 4558
rect 3528 4146 3556 8214
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3620 7002 3648 7822
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3620 5914 3648 6734
rect 3712 6458 3740 7754
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3712 6225 3740 6258
rect 3698 6216 3754 6225
rect 3698 6151 3754 6160
rect 3712 5914 3740 6151
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3712 5794 3740 5850
rect 3620 5766 3740 5794
rect 3620 4826 3648 5766
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 4146 3648 4422
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3712 4026 3740 5646
rect 3620 3998 3740 4026
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3620 3670 3648 3998
rect 3608 3664 3660 3670
rect 3804 3618 3832 9046
rect 3896 8922 3924 10610
rect 3988 9042 4016 11018
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10470 4108 10950
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9178 4108 9998
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4172 9110 4200 12200
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4356 11286 4384 12106
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10441 4384 11086
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4342 10432 4398 10441
rect 4342 10367 4398 10376
rect 4250 9616 4306 9625
rect 4250 9551 4306 9560
rect 4344 9580 4396 9586
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4068 8968 4120 8974
rect 3896 8894 4016 8922
rect 4264 8956 4292 9551
rect 4344 9522 4396 9528
rect 4068 8910 4120 8916
rect 4172 8928 4292 8956
rect 3988 7562 4016 8894
rect 4080 8294 4108 8910
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7993 4108 8230
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3608 3606 3660 3612
rect 3712 3590 3832 3618
rect 3896 7534 4016 7562
rect 3712 3534 3740 3590
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3712 3194 3740 3334
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3804 3097 3832 3130
rect 3790 3088 3846 3097
rect 3790 3023 3846 3032
rect 3252 2746 3372 2774
rect 3146 2408 3202 2417
rect 2964 2372 3016 2378
rect 3146 2343 3202 2352
rect 2964 2314 3016 2320
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 3252 2106 3280 2746
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 3528 1970 3556 2586
rect 3896 2106 3924 7534
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 6458 4016 6734
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3988 3058 4016 6258
rect 4080 5658 4108 7822
rect 4172 6225 4200 8928
rect 4356 8906 4384 9522
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4448 8090 4476 8502
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4158 6216 4214 6225
rect 4158 6151 4214 6160
rect 4264 5953 4292 7414
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4250 5944 4306 5953
rect 4250 5879 4306 5888
rect 4158 5808 4214 5817
rect 4158 5743 4160 5752
rect 4212 5743 4214 5752
rect 4160 5714 4212 5720
rect 4252 5704 4304 5710
rect 4080 5630 4200 5658
rect 4252 5646 4304 5652
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 4080 3398 4108 5199
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4080 2774 4108 3130
rect 3988 2746 4108 2774
rect 3988 2650 4016 2746
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4068 2576 4120 2582
rect 4066 2544 4068 2553
rect 4120 2544 4122 2553
rect 4066 2479 4122 2488
rect 4172 2106 4200 5630
rect 4264 5030 4292 5646
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4282 4292 4558
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4250 4176 4306 4185
rect 4250 4111 4306 4120
rect 4264 3602 4292 4111
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4356 3534 4384 6802
rect 4448 6322 4476 7686
rect 4540 7410 4568 10950
rect 4632 8401 4660 12200
rect 4804 11960 4856 11966
rect 4804 11902 4856 11908
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4724 10826 4752 11086
rect 4816 11014 4844 11902
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5000 11150 5028 11834
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4804 11008 4856 11014
rect 5092 10996 5120 12200
rect 5552 11744 5580 12200
rect 6012 12152 6040 12200
rect 6104 12152 6132 12294
rect 6012 12124 6132 12152
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 11762 5856 12038
rect 5816 11756 5868 11762
rect 5552 11716 5672 11744
rect 5538 11656 5594 11665
rect 5538 11591 5594 11600
rect 5552 11354 5580 11591
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 4804 10950 4856 10956
rect 5000 10968 5120 10996
rect 4724 10798 4936 10826
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 10130 4752 10542
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4618 8392 4674 8401
rect 4618 8327 4674 8336
rect 4618 8256 4674 8265
rect 4618 8191 4674 8200
rect 4632 8090 4660 8191
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4632 7290 4660 7686
rect 4540 7262 4660 7290
rect 4540 6866 4568 7262
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4434 6216 4490 6225
rect 4434 6151 4490 6160
rect 4448 4321 4476 6151
rect 4632 6118 4660 7142
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4526 5944 4582 5953
rect 4526 5879 4582 5888
rect 4540 5778 4568 5879
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4632 5166 4660 6054
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4434 4312 4490 4321
rect 4434 4247 4490 4256
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4448 3738 4476 4150
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4356 3058 4384 3470
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4356 2514 4384 2994
rect 4448 2582 4476 3538
rect 4540 3534 4568 4422
rect 4632 4078 4660 4626
rect 4724 4282 4752 9862
rect 4816 9489 4844 10678
rect 4802 9480 4858 9489
rect 4802 9415 4858 9424
rect 4908 9178 4936 10798
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4816 7886 4844 8842
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4802 7304 4858 7313
rect 4802 7239 4858 7248
rect 4816 6390 4844 7239
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4802 6080 4858 6089
rect 4802 6015 4858 6024
rect 4816 4706 4844 6015
rect 4908 5370 4936 8366
rect 5000 7313 5028 10968
rect 5066 10908 5374 10928
rect 5066 10906 5072 10908
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5368 10906 5374 10908
rect 5128 10854 5130 10906
rect 5310 10854 5312 10906
rect 5066 10852 5072 10854
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5368 10852 5374 10854
rect 5066 10832 5374 10852
rect 5078 10568 5134 10577
rect 5078 10503 5080 10512
rect 5132 10503 5134 10512
rect 5080 10474 5132 10480
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5538 10432 5594 10441
rect 5368 9908 5396 10406
rect 5538 10367 5594 10376
rect 5368 9880 5488 9908
rect 5066 9820 5374 9840
rect 5066 9818 5072 9820
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5368 9818 5374 9820
rect 5128 9766 5130 9818
rect 5310 9766 5312 9818
rect 5066 9764 5072 9766
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5368 9764 5374 9766
rect 5066 9744 5374 9764
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 8974 5304 9522
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 9178 5396 9318
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5066 8732 5374 8752
rect 5066 8730 5072 8732
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5368 8730 5374 8732
rect 5128 8678 5130 8730
rect 5310 8678 5312 8730
rect 5066 8676 5072 8678
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5368 8676 5374 8678
rect 5066 8656 5374 8676
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5092 8022 5120 8366
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5066 7644 5374 7664
rect 5066 7642 5072 7644
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5368 7642 5374 7644
rect 5128 7590 5130 7642
rect 5310 7590 5312 7642
rect 5066 7588 5072 7590
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5368 7588 5374 7590
rect 5066 7568 5374 7588
rect 4986 7304 5042 7313
rect 4986 7239 5042 7248
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6322 5028 7142
rect 5460 6798 5488 9880
rect 5552 9654 5580 10367
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5644 8378 5672 11716
rect 5816 11698 5868 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5920 11354 5948 11698
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5736 10713 5764 11086
rect 5722 10704 5778 10713
rect 6012 10674 6040 11086
rect 5722 10639 5778 10648
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5736 9586 5764 10542
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5552 8350 5672 8378
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5552 6644 5580 8350
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5460 6616 5580 6644
rect 5066 6556 5374 6576
rect 5066 6554 5072 6556
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5368 6554 5374 6556
rect 5128 6502 5130 6554
rect 5310 6502 5312 6554
rect 5066 6500 5072 6502
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5368 6500 5374 6502
rect 5066 6480 5374 6500
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5066 5468 5374 5488
rect 5066 5466 5072 5468
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5368 5466 5374 5468
rect 5128 5414 5130 5466
rect 5310 5414 5312 5466
rect 5066 5412 5072 5414
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5368 5412 5374 5414
rect 5066 5392 5374 5412
rect 4896 5364 4948 5370
rect 4948 5324 5120 5352
rect 4896 5306 4948 5312
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4826 4936 5170
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4816 4678 4936 4706
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4710 3768 4766 3777
rect 4710 3703 4712 3712
rect 4764 3703 4766 3712
rect 4712 3674 4764 3680
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4526 3360 4582 3369
rect 4526 3295 4582 3304
rect 4540 3058 4568 3295
rect 4632 3233 4660 3606
rect 4816 3602 4844 4422
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4908 3482 4936 4678
rect 5092 4622 5120 5324
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5368 4758 5396 5170
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5000 3641 5028 4422
rect 5066 4380 5374 4400
rect 5066 4378 5072 4380
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5368 4378 5374 4380
rect 5128 4326 5130 4378
rect 5310 4326 5312 4378
rect 5066 4324 5072 4326
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5368 4324 5374 4326
rect 5066 4304 5374 4324
rect 5460 4264 5488 6616
rect 5644 6361 5672 8230
rect 5630 6352 5686 6361
rect 5540 6316 5592 6322
rect 5630 6287 5686 6296
rect 5540 6258 5592 6264
rect 5552 5794 5580 6258
rect 5736 6186 5764 9386
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5722 6080 5778 6089
rect 5722 6015 5778 6024
rect 5552 5766 5672 5794
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5302 5580 5646
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5368 4236 5488 4264
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 4986 3632 5042 3641
rect 4986 3567 5042 3576
rect 5184 3505 5212 3878
rect 5276 3534 5304 4150
rect 5264 3528 5316 3534
rect 4724 3454 4936 3482
rect 5170 3496 5226 3505
rect 4618 3224 4674 3233
rect 4618 3159 4674 3168
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4618 2816 4674 2825
rect 4618 2751 4674 2760
rect 4526 2680 4582 2689
rect 4526 2615 4528 2624
rect 4580 2615 4582 2624
rect 4528 2586 4580 2592
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4632 2446 4660 2751
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4264 2106 4292 2246
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 4448 1834 4476 2314
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 1902 4568 2246
rect 4724 1970 4752 3454
rect 5264 3470 5316 3476
rect 5368 3482 5396 4236
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3777 5488 4082
rect 5446 3768 5502 3777
rect 5446 3703 5502 3712
rect 5446 3632 5502 3641
rect 5446 3567 5448 3576
rect 5500 3567 5502 3576
rect 5448 3538 5500 3544
rect 5368 3454 5488 3482
rect 5552 3466 5580 4966
rect 5644 4690 5672 5766
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5170 3431 5226 3440
rect 5066 3292 5374 3312
rect 5066 3290 5072 3292
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5368 3290 5374 3292
rect 5128 3238 5130 3290
rect 5310 3238 5312 3290
rect 5066 3236 5072 3238
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5368 3236 5374 3238
rect 4894 3224 4950 3233
rect 5066 3216 5374 3236
rect 4894 3159 4950 3168
rect 4908 3108 4936 3159
rect 4988 3120 5040 3126
rect 4908 3080 4988 3108
rect 4988 3062 5040 3068
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5262 2952 5318 2961
rect 5184 2650 5212 2926
rect 5262 2887 5318 2896
rect 5276 2689 5304 2887
rect 5460 2836 5488 3454
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5368 2808 5488 2836
rect 5262 2680 5318 2689
rect 5172 2644 5224 2650
rect 5262 2615 5318 2624
rect 5172 2586 5224 2592
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4816 1970 4844 2518
rect 5172 2440 5224 2446
rect 5368 2428 5396 2808
rect 5224 2400 5396 2428
rect 5172 2382 5224 2388
rect 5066 2204 5374 2224
rect 5066 2202 5072 2204
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5368 2202 5374 2204
rect 5128 2150 5130 2202
rect 5310 2150 5312 2202
rect 5066 2148 5072 2150
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5368 2148 5374 2150
rect 5066 2128 5374 2148
rect 4712 1964 4764 1970
rect 4712 1906 4764 1912
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 5644 1834 5672 3606
rect 5736 3534 5764 6015
rect 5828 5273 5856 9930
rect 5908 9376 5960 9382
rect 5906 9344 5908 9353
rect 5960 9344 5962 9353
rect 5906 9279 5962 9288
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5920 8430 5948 8842
rect 6012 8430 6040 10610
rect 6104 10606 6132 11290
rect 6196 10674 6224 11494
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6104 10266 6132 10542
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 9722 6224 9862
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7954 6040 8230
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6104 7834 6132 9590
rect 6182 9344 6238 9353
rect 6182 9279 6238 9288
rect 6012 7806 6132 7834
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 7002 5948 7346
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5906 6896 5962 6905
rect 5906 6831 5962 6840
rect 5920 6458 5948 6831
rect 6012 6798 6040 7806
rect 6196 7732 6224 9279
rect 6104 7704 6224 7732
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6012 5914 6040 6734
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6104 5794 6132 7704
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6196 7002 6224 7278
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 5920 5766 6132 5794
rect 5814 5264 5870 5273
rect 5814 5199 5870 5208
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5736 2553 5764 3295
rect 5828 2650 5856 5102
rect 5920 3097 5948 5766
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6012 4622 6040 5170
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6104 4570 6132 5646
rect 6196 5234 6224 6054
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6012 3738 6040 4558
rect 6104 4542 6224 4570
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6104 3602 6132 4422
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6000 3528 6052 3534
rect 6196 3482 6224 4542
rect 6000 3470 6052 3476
rect 6012 3126 6040 3470
rect 6104 3454 6224 3482
rect 6000 3120 6052 3126
rect 5906 3088 5962 3097
rect 6000 3062 6052 3068
rect 5906 3023 5962 3032
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6012 2582 6040 3062
rect 6000 2576 6052 2582
rect 5722 2544 5778 2553
rect 6000 2518 6052 2524
rect 5722 2479 5778 2488
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5828 2310 5856 2450
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6104 1902 6132 3454
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6196 3058 6224 3334
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6288 2582 6316 12294
rect 6458 12200 6514 13000
rect 16578 12608 16634 12617
rect 16578 12543 16634 12552
rect 9496 12232 9548 12238
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6380 9353 6408 9590
rect 6366 9344 6422 9353
rect 6366 9279 6422 9288
rect 6472 8378 6500 12200
rect 9496 12174 9548 12180
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 8760 12028 8812 12034
rect 8760 11970 8812 11976
rect 8668 11960 8720 11966
rect 8668 11902 8720 11908
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6656 11354 6684 11766
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6748 11234 6776 11494
rect 6656 11206 6776 11234
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 9722 6592 10542
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6380 8350 6500 8378
rect 6380 2825 6408 8350
rect 6656 7290 6684 11206
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6748 9518 6776 11018
rect 6840 10742 6868 11630
rect 7024 11354 7052 11766
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 7566 11452 7874 11472
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11376 7874 11396
rect 8128 11354 8156 11562
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7380 11212 7432 11218
rect 7576 11206 8064 11234
rect 7576 11200 7604 11206
rect 7432 11172 7604 11200
rect 7380 11154 7432 11160
rect 7288 11144 7340 11150
rect 7656 11144 7708 11150
rect 7288 11086 7340 11092
rect 7484 11104 7656 11132
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6918 10704 6974 10713
rect 6918 10639 6974 10648
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6840 9994 6868 10202
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6840 9897 6868 9930
rect 6826 9888 6882 9897
rect 6826 9823 6882 9832
rect 6932 9586 6960 10639
rect 7300 10577 7328 11086
rect 7286 10568 7342 10577
rect 7484 10538 7512 11104
rect 7656 11086 7708 11092
rect 7286 10503 7342 10512
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7484 10266 7512 10474
rect 7566 10364 7874 10384
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10288 7874 10308
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6736 9512 6788 9518
rect 7024 9466 7052 10202
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7932 10192 7984 10198
rect 7932 10134 7984 10140
rect 7392 9897 7420 10134
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7378 9888 7434 9897
rect 7378 9823 7434 9832
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 6736 9454 6788 9460
rect 6932 9438 7052 9466
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8566 6776 8910
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6748 7342 6776 8502
rect 6826 7712 6882 7721
rect 6826 7647 6882 7656
rect 6840 7478 6868 7647
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6460 7268 6512 7274
rect 6564 7262 6684 7290
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6564 7256 6592 7262
rect 6512 7228 6592 7256
rect 6460 7210 6512 7216
rect 6472 5817 6500 7210
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6458 5808 6514 5817
rect 6458 5743 6514 5752
rect 6564 5710 6592 6666
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6472 4026 6500 5578
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 4554 6592 5510
rect 6656 5409 6684 7142
rect 6932 7018 6960 9438
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 8498 7144 9318
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7886 7052 8230
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7208 7426 7236 9658
rect 7288 8968 7340 8974
rect 7392 8956 7420 9823
rect 7668 9722 7696 9930
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7656 9580 7708 9586
rect 7760 9568 7788 9998
rect 7708 9540 7788 9568
rect 7656 9522 7708 9528
rect 7566 9276 7874 9296
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9200 7874 9220
rect 7340 8928 7420 8956
rect 7288 8910 7340 8916
rect 7392 8922 7420 8928
rect 7392 8906 7696 8922
rect 7392 8900 7708 8906
rect 7392 8894 7656 8900
rect 7656 8842 7708 8848
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 7886 7512 8774
rect 7566 8188 7874 8208
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8112 7874 8132
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7116 7398 7236 7426
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6840 6990 6960 7018
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6642 5400 6698 5409
rect 6642 5335 6698 5344
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6564 4146 6592 4490
rect 6748 4282 6776 6258
rect 6840 6089 6868 6990
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6826 6080 6882 6089
rect 6826 6015 6882 6024
rect 6932 5794 6960 6802
rect 6840 5778 6960 5794
rect 6828 5772 6960 5778
rect 6880 5766 6960 5772
rect 6828 5714 6880 5720
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6472 3998 6684 4026
rect 6458 3768 6514 3777
rect 6458 3703 6514 3712
rect 6472 2922 6500 3703
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6366 2816 6422 2825
rect 6366 2751 6422 2760
rect 6564 2650 6592 3470
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6276 2576 6328 2582
rect 6276 2518 6328 2524
rect 6656 2514 6684 3998
rect 6748 3777 6776 4082
rect 6734 3768 6790 3777
rect 6734 3703 6790 3712
rect 6840 3482 6868 5510
rect 6932 4690 6960 5766
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3602 6960 3878
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6748 3454 6868 3482
rect 6748 3058 6776 3454
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6840 2446 6868 3334
rect 7024 2774 7052 7278
rect 7116 6730 7144 7398
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7208 6458 7236 7210
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7194 5944 7250 5953
rect 7194 5879 7250 5888
rect 7208 5574 7236 5879
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6932 2746 7052 2774
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6092 1896 6144 1902
rect 6092 1838 6144 1844
rect 4436 1828 4488 1834
rect 4436 1770 4488 1776
rect 5632 1828 5684 1834
rect 5632 1770 5684 1776
rect 6932 1562 6960 2746
rect 7116 2650 7144 5170
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7208 1986 7236 5034
rect 7300 4826 7328 6190
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 3618 7328 4422
rect 7392 4185 7420 7686
rect 7484 7002 7512 7822
rect 7566 7100 7874 7120
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7024 7874 7044
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7852 6730 7880 6870
rect 7840 6724 7892 6730
rect 7484 6684 7840 6712
rect 7484 5624 7512 6684
rect 7840 6666 7892 6672
rect 7566 6012 7874 6032
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5936 7874 5956
rect 7564 5636 7616 5642
rect 7484 5596 7564 5624
rect 7564 5578 7616 5584
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7484 4282 7512 5238
rect 7566 4924 7874 4944
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4848 7874 4868
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7378 4176 7434 4185
rect 7378 4111 7434 4120
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 3720 7512 4082
rect 7746 4040 7802 4049
rect 7852 4010 7880 4626
rect 7746 3975 7748 3984
rect 7800 3975 7802 3984
rect 7840 4004 7892 4010
rect 7748 3946 7800 3952
rect 7840 3946 7892 3952
rect 7566 3836 7874 3856
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3760 7874 3780
rect 7484 3692 7696 3720
rect 7300 3590 7512 3618
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 2582 7420 3334
rect 7484 3126 7512 3590
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7668 2836 7696 3692
rect 7838 3632 7894 3641
rect 7838 3567 7894 3576
rect 7852 3233 7880 3567
rect 7838 3224 7894 3233
rect 7838 3159 7894 3168
rect 7484 2808 7696 2836
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7484 2038 7512 2808
rect 7566 2748 7874 2768
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2672 7874 2692
rect 7840 2440 7892 2446
rect 7838 2408 7840 2417
rect 7892 2408 7894 2417
rect 7838 2343 7894 2352
rect 7024 1970 7236 1986
rect 7472 2032 7524 2038
rect 7472 1974 7524 1980
rect 7012 1964 7236 1970
rect 7064 1958 7236 1964
rect 7012 1906 7064 1912
rect 7024 1562 7052 1906
rect 7472 1760 7524 1766
rect 7472 1702 7524 1708
rect 2504 1556 2556 1562
rect 2504 1498 2556 1504
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 7012 1556 7064 1562
rect 7012 1498 7064 1504
rect 7484 1494 7512 1702
rect 7566 1660 7874 1680
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1584 7874 1604
rect 7472 1488 7524 1494
rect 7472 1430 7524 1436
rect 7944 1290 7972 10134
rect 8036 4690 8064 11206
rect 8312 11150 8340 11494
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 8673 8156 10406
rect 8220 10266 8248 10678
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8220 9926 8248 10202
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 9178 8248 9454
rect 8312 9382 8340 10950
rect 8404 10266 8432 11834
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8482 10568 8538 10577
rect 8482 10503 8538 10512
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8114 8664 8170 8673
rect 8114 8599 8170 8608
rect 8220 8514 8248 8842
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8128 8486 8248 8514
rect 8128 7206 8156 8486
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8404 8378 8432 8774
rect 8496 8634 8524 10503
rect 8588 10266 8616 11086
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9042 8616 9998
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6934 8156 7142
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 2582 8064 4422
rect 8128 3369 8156 6394
rect 8220 5846 8248 8366
rect 8404 8350 8524 8378
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7002 8340 7686
rect 8404 7546 8432 7754
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8312 5778 8340 6598
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8206 5672 8262 5681
rect 8206 5607 8262 5616
rect 8220 3738 8248 5607
rect 8404 5386 8432 7278
rect 8496 6730 8524 8350
rect 8588 8022 8616 8978
rect 8680 8566 8708 11902
rect 8772 10810 8800 11970
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8772 9110 8800 10406
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8772 8090 8800 8910
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8588 6934 8616 7958
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8680 6662 8708 7822
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8772 5710 8800 7686
rect 8864 6322 8892 11222
rect 9036 11120 9088 11126
rect 9036 11062 9088 11068
rect 9048 10713 9076 11062
rect 9034 10704 9090 10713
rect 9034 10639 9090 10648
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6458 8984 6598
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9048 6236 9076 10406
rect 8956 6208 9076 6236
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8956 5522 8984 6208
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 8312 5358 8432 5386
rect 8496 5494 8984 5522
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8206 3632 8262 3641
rect 8206 3567 8262 3576
rect 8114 3360 8170 3369
rect 8114 3295 8170 3304
rect 8220 3058 8248 3567
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 8128 2446 8156 2926
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8116 2440 8168 2446
rect 8022 2408 8078 2417
rect 8116 2382 8168 2388
rect 8022 2343 8078 2352
rect 8036 2310 8064 2343
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8220 2038 8248 2790
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8312 1834 8340 5358
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8404 2582 8432 5170
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 8404 1426 8432 2246
rect 8496 1970 8524 5494
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8588 3534 8616 4082
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8588 3194 8616 3334
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 8588 1766 8616 2994
rect 8680 2854 8708 4014
rect 8772 3777 8800 5306
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8666 2544 8722 2553
rect 8666 2479 8722 2488
rect 8576 1760 8628 1766
rect 8576 1702 8628 1708
rect 8680 1562 8708 2479
rect 8772 1834 8800 3402
rect 8864 2553 8892 4150
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8956 3058 8984 4082
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 9048 2650 9076 6054
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8850 2544 8906 2553
rect 8850 2479 8906 2488
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8864 1970 8892 2246
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 9048 1884 9076 2450
rect 9140 2106 9168 11222
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 9232 7342 9260 10474
rect 9324 9654 9352 12038
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 6866 9260 7278
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 3942 9260 6598
rect 9324 5370 9352 9046
rect 9416 8498 9444 12106
rect 9508 9586 9536 12174
rect 13450 11928 13506 11937
rect 13450 11863 13506 11872
rect 13544 11892 13596 11898
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9416 5250 9444 7142
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9508 5914 9536 6258
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9416 5222 9536 5250
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9218 3768 9274 3777
rect 9218 3703 9220 3712
rect 9272 3703 9274 3712
rect 9220 3674 9272 3680
rect 9218 3360 9274 3369
rect 9218 3295 9274 3304
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 9232 1970 9260 3295
rect 9220 1964 9272 1970
rect 9220 1906 9272 1912
rect 8956 1856 9076 1884
rect 8956 1850 8984 1856
rect 8760 1828 8812 1834
rect 8760 1770 8812 1776
rect 8864 1822 8984 1850
rect 8864 1766 8892 1822
rect 8852 1760 8904 1766
rect 8852 1702 8904 1708
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 9128 1420 9180 1426
rect 9128 1362 9180 1368
rect 8944 1352 8996 1358
rect 8942 1320 8944 1329
rect 8996 1320 8998 1329
rect 7932 1284 7984 1290
rect 8942 1255 8998 1264
rect 7932 1226 7984 1232
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 3344 241 3372 1158
rect 5066 1116 5374 1136
rect 5066 1114 5072 1116
rect 5128 1114 5152 1116
rect 5208 1114 5232 1116
rect 5288 1114 5312 1116
rect 5368 1114 5374 1116
rect 5128 1062 5130 1114
rect 5310 1062 5312 1114
rect 5066 1060 5072 1062
rect 5128 1060 5152 1062
rect 5208 1060 5232 1062
rect 5288 1060 5312 1062
rect 5368 1060 5374 1062
rect 5066 1040 5374 1060
rect 9140 513 9168 1362
rect 9324 921 9352 4966
rect 9416 1222 9444 5102
rect 9508 3482 9536 5222
rect 9600 4078 9628 10610
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8265 9720 8842
rect 9678 8256 9734 8265
rect 9678 8191 9734 8200
rect 10428 6225 10456 11018
rect 10414 6216 10470 6225
rect 10414 6151 10470 6160
rect 9678 4992 9734 5001
rect 9678 4927 9734 4936
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9692 3641 9720 4927
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9678 3632 9734 3641
rect 9678 3567 9734 3576
rect 9784 3482 9812 4218
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9508 3454 9628 3482
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 1358 9536 3334
rect 9600 2446 9628 3454
rect 9692 3454 9812 3482
rect 9692 2650 9720 3454
rect 9772 2984 9824 2990
rect 9876 2961 9904 3538
rect 13464 3194 13492 11863
rect 13544 11834 13596 11840
rect 13556 7585 13584 11834
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 7857 13676 11154
rect 13726 11112 13782 11121
rect 13726 11047 13782 11056
rect 13634 7848 13690 7857
rect 13634 7783 13690 7792
rect 13542 7576 13598 7585
rect 13542 7511 13598 7520
rect 13634 4584 13690 4593
rect 13634 4519 13690 4528
rect 13648 3194 13676 4519
rect 13740 3670 13768 11047
rect 13832 10305 13860 11698
rect 13818 10296 13874 10305
rect 13818 10231 13874 10240
rect 13818 10160 13874 10169
rect 13818 10095 13874 10104
rect 13832 10062 13860 10095
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13818 9072 13874 9081
rect 13818 9007 13874 9016
rect 13832 7721 13860 9007
rect 13818 7712 13874 7721
rect 13818 7647 13874 7656
rect 13818 5808 13874 5817
rect 13818 5743 13820 5752
rect 13872 5743 13874 5752
rect 13820 5714 13872 5720
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4185 13860 5034
rect 13818 4176 13874 4185
rect 13818 4111 13874 4120
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13832 3777 13860 3946
rect 13818 3768 13874 3777
rect 13818 3703 13874 3712
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 16592 3602 16620 12543
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22190 9888 22246 9897
rect 22190 9823 22246 9832
rect 22098 9480 22154 9489
rect 22098 9415 22154 9424
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 13818 3360 13874 3369
rect 13818 3295 13820 3304
rect 13872 3295 13874 3304
rect 16764 3324 16816 3330
rect 13820 3266 13872 3272
rect 16764 3266 16816 3272
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 9772 2926 9824 2932
rect 9862 2952 9918 2961
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9784 2514 9812 2926
rect 9862 2887 9918 2896
rect 13818 2952 13874 2961
rect 13818 2887 13820 2896
rect 13872 2887 13874 2896
rect 13820 2858 13872 2864
rect 16670 2544 16726 2553
rect 9772 2508 9824 2514
rect 16670 2479 16726 2488
rect 9772 2450 9824 2456
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 13818 2408 13874 2417
rect 13818 2343 13820 2352
rect 13872 2343 13874 2352
rect 13820 2314 13872 2320
rect 16578 2136 16634 2145
rect 16578 2071 16634 2080
rect 16592 1834 16620 2071
rect 16684 1902 16712 2479
rect 16776 2310 16804 3266
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16868 2378 16896 3130
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16672 1896 16724 1902
rect 16672 1838 16724 1844
rect 16580 1828 16632 1834
rect 16580 1770 16632 1776
rect 16578 1728 16634 1737
rect 16578 1663 16634 1672
rect 16592 1358 16620 1663
rect 16960 1562 16988 5714
rect 16948 1556 17000 1562
rect 16948 1498 17000 1504
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9310 912 9366 921
rect 9310 847 9366 856
rect 9126 504 9182 513
rect 9126 439 9182 448
rect 22112 241 22140 9415
rect 22204 2922 22232 9823
rect 22296 6633 22324 9998
rect 22282 6624 22338 6633
rect 22282 6559 22338 6568
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 3330 232 3386 241
rect 3330 167 3386 176
rect 22098 232 22154 241
rect 22098 167 22154 176
<< via2 >>
rect 1398 10804 1454 10840
rect 1398 10784 1400 10804
rect 1400 10784 1452 10804
rect 1452 10784 1454 10804
rect 1214 10648 1270 10704
rect 1306 9424 1362 9480
rect 1674 10104 1730 10160
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2870 10804 2926 10840
rect 2870 10784 2872 10804
rect 2872 10784 2924 10804
rect 2924 10784 2926 10804
rect 2778 10512 2834 10568
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2594 10104 2650 10160
rect 2778 10104 2834 10160
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2042 8472 2098 8528
rect 2410 8880 2466 8936
rect 1858 6296 1914 6352
rect 1950 5752 2006 5808
rect 3054 9016 3110 9072
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2594 7928 2650 7984
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 3238 10104 3294 10160
rect 3330 9696 3386 9752
rect 3238 9016 3294 9072
rect 3606 10104 3662 10160
rect 3146 8336 3202 8392
rect 2502 6160 2558 6216
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 3054 5888 3110 5944
rect 3790 9152 3846 9208
rect 3238 6160 3294 6216
rect 2962 5652 2964 5672
rect 2964 5652 3016 5672
rect 3016 5652 3018 5672
rect 2962 5616 3018 5652
rect 3422 5628 3424 5672
rect 3424 5628 3476 5672
rect 3476 5628 3478 5672
rect 3422 5616 3478 5628
rect 3698 6160 3754 6216
rect 4342 10376 4398 10432
rect 4250 9560 4306 9616
rect 4066 7928 4122 7984
rect 3790 3032 3846 3088
rect 3146 2352 3202 2408
rect 4158 6160 4214 6216
rect 4250 5888 4306 5944
rect 4158 5772 4214 5808
rect 4158 5752 4160 5772
rect 4160 5752 4212 5772
rect 4212 5752 4214 5772
rect 4066 5208 4122 5264
rect 4066 2524 4068 2544
rect 4068 2524 4120 2544
rect 4120 2524 4122 2544
rect 4066 2488 4122 2524
rect 4250 4120 4306 4176
rect 5538 11600 5594 11656
rect 4618 8336 4674 8392
rect 4618 8200 4674 8256
rect 4434 6160 4490 6216
rect 4526 5888 4582 5944
rect 4434 4256 4490 4312
rect 4802 9424 4858 9480
rect 4802 7248 4858 7304
rect 4802 6024 4858 6080
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5118 10906
rect 5118 10854 5128 10906
rect 5152 10854 5182 10906
rect 5182 10854 5194 10906
rect 5194 10854 5208 10906
rect 5232 10854 5246 10906
rect 5246 10854 5258 10906
rect 5258 10854 5288 10906
rect 5312 10854 5322 10906
rect 5322 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 5078 10532 5134 10568
rect 5078 10512 5080 10532
rect 5080 10512 5132 10532
rect 5132 10512 5134 10532
rect 5538 10376 5594 10432
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5118 9818
rect 5118 9766 5128 9818
rect 5152 9766 5182 9818
rect 5182 9766 5194 9818
rect 5194 9766 5208 9818
rect 5232 9766 5246 9818
rect 5246 9766 5258 9818
rect 5258 9766 5288 9818
rect 5312 9766 5322 9818
rect 5322 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5118 8730
rect 5118 8678 5128 8730
rect 5152 8678 5182 8730
rect 5182 8678 5194 8730
rect 5194 8678 5208 8730
rect 5232 8678 5246 8730
rect 5246 8678 5258 8730
rect 5258 8678 5288 8730
rect 5312 8678 5322 8730
rect 5322 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5118 7642
rect 5118 7590 5128 7642
rect 5152 7590 5182 7642
rect 5182 7590 5194 7642
rect 5194 7590 5208 7642
rect 5232 7590 5246 7642
rect 5246 7590 5258 7642
rect 5258 7590 5288 7642
rect 5312 7590 5322 7642
rect 5322 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 4986 7248 5042 7304
rect 5722 10648 5778 10704
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5118 6554
rect 5118 6502 5128 6554
rect 5152 6502 5182 6554
rect 5182 6502 5194 6554
rect 5194 6502 5208 6554
rect 5232 6502 5246 6554
rect 5246 6502 5258 6554
rect 5258 6502 5288 6554
rect 5312 6502 5322 6554
rect 5322 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5118 5466
rect 5118 5414 5128 5466
rect 5152 5414 5182 5466
rect 5182 5414 5194 5466
rect 5194 5414 5208 5466
rect 5232 5414 5246 5466
rect 5246 5414 5258 5466
rect 5258 5414 5288 5466
rect 5312 5414 5322 5466
rect 5322 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 4710 3732 4766 3768
rect 4710 3712 4712 3732
rect 4712 3712 4764 3732
rect 4764 3712 4766 3732
rect 4526 3304 4582 3360
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5118 4378
rect 5118 4326 5128 4378
rect 5152 4326 5182 4378
rect 5182 4326 5194 4378
rect 5194 4326 5208 4378
rect 5232 4326 5246 4378
rect 5246 4326 5258 4378
rect 5258 4326 5288 4378
rect 5312 4326 5322 4378
rect 5322 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 5630 6296 5686 6352
rect 5722 6024 5778 6080
rect 4986 3576 5042 3632
rect 4618 3168 4674 3224
rect 4618 2760 4674 2816
rect 4526 2644 4582 2680
rect 4526 2624 4528 2644
rect 4528 2624 4580 2644
rect 4580 2624 4582 2644
rect 5170 3440 5226 3496
rect 5446 3712 5502 3768
rect 5446 3596 5502 3632
rect 5446 3576 5448 3596
rect 5448 3576 5500 3596
rect 5500 3576 5502 3596
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5118 3290
rect 5118 3238 5128 3290
rect 5152 3238 5182 3290
rect 5182 3238 5194 3290
rect 5194 3238 5208 3290
rect 5232 3238 5246 3290
rect 5246 3238 5258 3290
rect 5258 3238 5288 3290
rect 5312 3238 5322 3290
rect 5322 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 4894 3168 4950 3224
rect 5262 2896 5318 2952
rect 5262 2624 5318 2680
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5118 2202
rect 5118 2150 5128 2202
rect 5152 2150 5182 2202
rect 5182 2150 5194 2202
rect 5194 2150 5208 2202
rect 5232 2150 5246 2202
rect 5246 2150 5258 2202
rect 5258 2150 5288 2202
rect 5312 2150 5322 2202
rect 5322 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 5906 9324 5908 9344
rect 5908 9324 5960 9344
rect 5960 9324 5962 9344
rect 5906 9288 5962 9324
rect 6182 9288 6238 9344
rect 5906 6840 5962 6896
rect 5814 5208 5870 5264
rect 5722 3304 5778 3360
rect 5906 3032 5962 3088
rect 5722 2488 5778 2544
rect 16578 12552 16634 12608
rect 6366 9288 6422 9344
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 6918 10648 6974 10704
rect 6826 9832 6882 9888
rect 7286 10512 7342 10568
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 7378 9832 7434 9888
rect 6826 7656 6882 7712
rect 6458 5752 6514 5808
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 6642 5344 6698 5400
rect 6826 6024 6882 6080
rect 6458 3712 6514 3768
rect 6366 2760 6422 2816
rect 6734 3712 6790 3768
rect 7194 5888 7250 5944
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7378 4120 7434 4176
rect 7746 4004 7802 4040
rect 7746 3984 7748 4004
rect 7748 3984 7800 4004
rect 7800 3984 7802 4004
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 7838 3576 7894 3632
rect 7838 3168 7894 3224
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 7838 2388 7840 2408
rect 7840 2388 7892 2408
rect 7892 2388 7894 2408
rect 7838 2352 7894 2388
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 8482 10512 8538 10568
rect 8114 8608 8170 8664
rect 8206 5616 8262 5672
rect 9034 10648 9090 10704
rect 8206 3576 8262 3632
rect 8114 3304 8170 3360
rect 8022 2352 8078 2408
rect 8758 3712 8814 3768
rect 8666 2488 8722 2544
rect 8850 2488 8906 2544
rect 13450 11872 13506 11928
rect 9218 3732 9274 3768
rect 9218 3712 9220 3732
rect 9220 3712 9272 3732
rect 9272 3712 9274 3732
rect 9218 3304 9274 3360
rect 8942 1300 8944 1320
rect 8944 1300 8996 1320
rect 8996 1300 8998 1320
rect 8942 1264 8998 1300
rect 5072 1114 5128 1116
rect 5152 1114 5208 1116
rect 5232 1114 5288 1116
rect 5312 1114 5368 1116
rect 5072 1062 5118 1114
rect 5118 1062 5128 1114
rect 5152 1062 5182 1114
rect 5182 1062 5194 1114
rect 5194 1062 5208 1114
rect 5232 1062 5246 1114
rect 5246 1062 5258 1114
rect 5258 1062 5288 1114
rect 5312 1062 5322 1114
rect 5322 1062 5368 1114
rect 5072 1060 5128 1062
rect 5152 1060 5208 1062
rect 5232 1060 5288 1062
rect 5312 1060 5368 1062
rect 9678 8200 9734 8256
rect 10414 6160 10470 6216
rect 9678 4936 9734 4992
rect 9678 3576 9734 3632
rect 13726 11056 13782 11112
rect 13634 7792 13690 7848
rect 13542 7520 13598 7576
rect 13634 4528 13690 4584
rect 13818 10240 13874 10296
rect 13818 10104 13874 10160
rect 13818 9016 13874 9072
rect 13818 7656 13874 7712
rect 13818 5772 13874 5808
rect 13818 5752 13820 5772
rect 13820 5752 13872 5772
rect 13872 5752 13874 5772
rect 13818 4120 13874 4176
rect 13818 3712 13874 3768
rect 22190 9832 22246 9888
rect 22098 9424 22154 9480
rect 13818 3324 13874 3360
rect 13818 3304 13820 3324
rect 13820 3304 13872 3324
rect 13872 3304 13874 3324
rect 9862 2896 9918 2952
rect 13818 2916 13874 2952
rect 13818 2896 13820 2916
rect 13820 2896 13872 2916
rect 13872 2896 13874 2916
rect 16670 2488 16726 2544
rect 13818 2372 13874 2408
rect 13818 2352 13820 2372
rect 13820 2352 13872 2372
rect 13872 2352 13874 2372
rect 16578 2080 16634 2136
rect 16578 1672 16634 1728
rect 9310 856 9366 912
rect 9126 448 9182 504
rect 22282 6568 22338 6624
rect 3330 176 3386 232
rect 22098 176 22154 232
<< metal3 >>
rect 16573 12610 16639 12613
rect 13862 12608 16639 12610
rect 13862 12552 16578 12608
rect 16634 12552 16639 12608
rect 13862 12550 16639 12552
rect 13862 12338 13922 12550
rect 16573 12547 16639 12550
rect 14000 12338 34000 12368
rect 13862 12278 34000 12338
rect 14000 12248 34000 12278
rect 13445 11930 13511 11933
rect 14000 11930 34000 11960
rect 13445 11928 34000 11930
rect 13445 11872 13450 11928
rect 13506 11872 34000 11928
rect 13445 11870 34000 11872
rect 13445 11867 13511 11870
rect 14000 11840 34000 11870
rect 5533 11658 5599 11661
rect 5533 11656 12450 11658
rect 5533 11600 5538 11656
rect 5594 11600 12450 11656
rect 5533 11598 12450 11600
rect 5533 11595 5599 11598
rect 12390 11522 12450 11598
rect 14000 11522 34000 11552
rect 12390 11462 34000 11522
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 7560 11456 7880 11457
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 14000 11432 34000 11462
rect 7560 11391 7880 11392
rect 13721 11114 13787 11117
rect 14000 11114 34000 11144
rect 13721 11112 34000 11114
rect 13721 11056 13726 11112
rect 13782 11056 34000 11112
rect 13721 11054 34000 11056
rect 13721 11051 13787 11054
rect 14000 11024 34000 11054
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10847 5380 10848
rect 1393 10842 1459 10845
rect 2865 10842 2931 10845
rect 1393 10840 2931 10842
rect 1393 10784 1398 10840
rect 1454 10784 2870 10840
rect 2926 10784 2931 10840
rect 1393 10782 2931 10784
rect 1393 10779 1459 10782
rect 2865 10779 2931 10782
rect 1209 10706 1275 10709
rect 5717 10706 5783 10709
rect 1209 10704 5783 10706
rect 1209 10648 1214 10704
rect 1270 10648 5722 10704
rect 5778 10648 5783 10704
rect 1209 10646 5783 10648
rect 1209 10643 1275 10646
rect 5717 10643 5783 10646
rect 6913 10706 6979 10709
rect 9029 10706 9095 10709
rect 14000 10706 34000 10736
rect 6913 10704 34000 10706
rect 6913 10648 6918 10704
rect 6974 10648 9034 10704
rect 9090 10648 34000 10704
rect 6913 10646 34000 10648
rect 6913 10643 6979 10646
rect 9029 10643 9095 10646
rect 14000 10616 34000 10646
rect 2773 10570 2839 10573
rect 5073 10570 5139 10573
rect 2773 10568 5139 10570
rect 2773 10512 2778 10568
rect 2834 10512 5078 10568
rect 5134 10512 5139 10568
rect 2773 10510 5139 10512
rect 2773 10507 2839 10510
rect 5073 10507 5139 10510
rect 7281 10570 7347 10573
rect 8477 10570 8543 10573
rect 7281 10568 8543 10570
rect 7281 10512 7286 10568
rect 7342 10512 8482 10568
rect 8538 10512 8543 10568
rect 7281 10510 8543 10512
rect 7281 10507 7347 10510
rect 8477 10507 8543 10510
rect 4337 10434 4403 10437
rect 5533 10434 5599 10437
rect 4337 10432 5599 10434
rect 4337 10376 4342 10432
rect 4398 10376 5538 10432
rect 5594 10376 5599 10432
rect 4337 10374 5599 10376
rect 4337 10371 4403 10374
rect 5533 10371 5599 10374
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 7560 10368 7880 10369
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 10303 7880 10304
rect 13813 10298 13879 10301
rect 14000 10298 34000 10328
rect 13813 10296 34000 10298
rect 13813 10240 13818 10296
rect 13874 10240 34000 10296
rect 13813 10238 34000 10240
rect 13813 10235 13879 10238
rect 14000 10208 34000 10238
rect 1669 10162 1735 10165
rect 2589 10162 2655 10165
rect 1669 10160 2655 10162
rect 1669 10104 1674 10160
rect 1730 10104 2594 10160
rect 2650 10104 2655 10160
rect 1669 10102 2655 10104
rect 1669 10099 1735 10102
rect 2589 10099 2655 10102
rect 2773 10162 2839 10165
rect 3233 10162 3299 10165
rect 2773 10160 3299 10162
rect 2773 10104 2778 10160
rect 2834 10104 3238 10160
rect 3294 10104 3299 10160
rect 2773 10102 3299 10104
rect 2773 10099 2839 10102
rect 3233 10099 3299 10102
rect 3601 10162 3667 10165
rect 13813 10162 13879 10165
rect 3601 10160 13879 10162
rect 3601 10104 3606 10160
rect 3662 10104 13818 10160
rect 13874 10104 13879 10160
rect 3601 10102 13879 10104
rect 3601 10099 3667 10102
rect 13813 10099 13879 10102
rect 6821 9890 6887 9893
rect 7373 9890 7439 9893
rect 6821 9888 7439 9890
rect 6821 9832 6826 9888
rect 6882 9832 7378 9888
rect 7434 9832 7439 9888
rect 6821 9830 7439 9832
rect 6821 9827 6887 9830
rect 7373 9827 7439 9830
rect 14000 9888 34000 9920
rect 14000 9832 22190 9888
rect 22246 9832 34000 9888
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9832
rect 5060 9759 5380 9760
rect 3325 9754 3391 9757
rect 3325 9752 3434 9754
rect 3325 9696 3330 9752
rect 3386 9696 3434 9752
rect 3325 9691 3434 9696
rect 3374 9618 3434 9691
rect 4245 9618 4311 9621
rect 3374 9616 4311 9618
rect 3374 9560 4250 9616
rect 4306 9560 4311 9616
rect 3374 9558 4311 9560
rect 4245 9555 4311 9558
rect 1301 9482 1367 9485
rect 4797 9482 4863 9485
rect 1301 9480 4863 9482
rect 1301 9424 1306 9480
rect 1362 9424 4802 9480
rect 4858 9424 4863 9480
rect 1301 9422 4863 9424
rect 1301 9419 1367 9422
rect 4797 9419 4863 9422
rect 14000 9480 34000 9512
rect 14000 9424 22098 9480
rect 22154 9424 34000 9480
rect 14000 9392 34000 9424
rect 5901 9346 5967 9349
rect 6177 9346 6243 9349
rect 6361 9346 6427 9349
rect 5901 9344 6427 9346
rect 5901 9288 5906 9344
rect 5962 9288 6182 9344
rect 6238 9288 6366 9344
rect 6422 9288 6427 9344
rect 5901 9286 6427 9288
rect 5901 9283 5967 9286
rect 6177 9283 6243 9286
rect 6361 9283 6427 9286
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 7560 9280 7880 9281
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9215 7880 9216
rect 3785 9208 3851 9213
rect 3785 9152 3790 9208
rect 3846 9152 3851 9208
rect 3785 9147 3851 9152
rect 3049 9074 3115 9077
rect 3233 9074 3299 9077
rect 3049 9072 3299 9074
rect 3049 9016 3054 9072
rect 3110 9016 3238 9072
rect 3294 9016 3299 9072
rect 3049 9014 3299 9016
rect 3049 9011 3115 9014
rect 3233 9011 3299 9014
rect 2405 8938 2471 8941
rect 3788 8938 3848 9147
rect 13813 9074 13879 9077
rect 14000 9074 34000 9104
rect 13813 9072 34000 9074
rect 13813 9016 13818 9072
rect 13874 9016 34000 9072
rect 13813 9014 34000 9016
rect 13813 9011 13879 9014
rect 14000 8984 34000 9014
rect 2405 8936 3848 8938
rect 2405 8880 2410 8936
rect 2466 8880 3848 8936
rect 2405 8878 3848 8880
rect 2405 8875 2471 8878
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 8671 5380 8672
rect 8109 8666 8175 8669
rect 14000 8666 34000 8696
rect 8109 8664 34000 8666
rect 8109 8608 8114 8664
rect 8170 8608 34000 8664
rect 8109 8606 34000 8608
rect 8109 8603 8175 8606
rect 14000 8576 34000 8606
rect 2037 8530 2103 8533
rect 2037 8528 2652 8530
rect 2037 8472 2042 8528
rect 2098 8472 2652 8528
rect 2037 8470 2652 8472
rect 2037 8467 2103 8470
rect 2592 8394 2652 8470
rect 3141 8394 3207 8397
rect 4613 8394 4679 8397
rect 2592 8334 3066 8394
rect 3006 8258 3066 8334
rect 3141 8392 4679 8394
rect 3141 8336 3146 8392
rect 3202 8336 4618 8392
rect 4674 8336 4679 8392
rect 3141 8334 4679 8336
rect 3141 8331 3207 8334
rect 4613 8331 4679 8334
rect 4613 8258 4679 8261
rect 3006 8256 4679 8258
rect 3006 8200 4618 8256
rect 4674 8200 4679 8256
rect 3006 8198 4679 8200
rect 4613 8195 4679 8198
rect 9673 8258 9739 8261
rect 14000 8258 34000 8288
rect 9673 8256 34000 8258
rect 9673 8200 9678 8256
rect 9734 8200 34000 8256
rect 9673 8198 34000 8200
rect 9673 8195 9739 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 7560 8192 7880 8193
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 14000 8168 34000 8198
rect 7560 8127 7880 8128
rect 2589 7986 2655 7989
rect 4061 7986 4127 7989
rect 2589 7984 4127 7986
rect 2589 7928 2594 7984
rect 2650 7928 4066 7984
rect 4122 7928 4127 7984
rect 2589 7926 4127 7928
rect 2589 7923 2655 7926
rect 4061 7923 4127 7926
rect 13629 7850 13695 7853
rect 14000 7850 34000 7880
rect 13629 7848 34000 7850
rect 13629 7792 13634 7848
rect 13690 7792 34000 7848
rect 13629 7790 34000 7792
rect 13629 7787 13695 7790
rect 14000 7760 34000 7790
rect 6821 7714 6887 7717
rect 13813 7714 13879 7717
rect 6821 7712 13879 7714
rect 6821 7656 6826 7712
rect 6882 7656 13818 7712
rect 13874 7656 13879 7712
rect 6821 7654 13879 7656
rect 6821 7651 6887 7654
rect 13813 7651 13879 7654
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7583 5380 7584
rect 13537 7578 13603 7581
rect 13537 7576 13922 7578
rect 13537 7520 13542 7576
rect 13598 7520 13922 7576
rect 13537 7518 13922 7520
rect 13537 7515 13603 7518
rect 13862 7442 13922 7518
rect 14000 7442 34000 7472
rect 13862 7382 34000 7442
rect 14000 7352 34000 7382
rect 4797 7306 4863 7309
rect 4981 7306 5047 7309
rect 4797 7304 5047 7306
rect 4797 7248 4802 7304
rect 4858 7248 4986 7304
rect 5042 7248 5047 7304
rect 4797 7246 5047 7248
rect 4797 7243 4863 7246
rect 4981 7243 5047 7246
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 7560 7104 7880 7105
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 7039 7880 7040
rect 14000 7034 34000 7064
rect 13862 6974 34000 7034
rect 5901 6898 5967 6901
rect 13862 6898 13922 6974
rect 14000 6944 34000 6974
rect 5901 6896 13922 6898
rect 5901 6840 5906 6896
rect 5962 6840 13922 6896
rect 5901 6838 13922 6840
rect 5901 6835 5967 6838
rect 14000 6624 34000 6656
rect 14000 6568 22282 6624
rect 22338 6568 34000 6624
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6568
rect 5060 6495 5380 6496
rect 1853 6354 1919 6357
rect 5625 6354 5691 6357
rect 1853 6352 5691 6354
rect 1853 6296 1858 6352
rect 1914 6296 5630 6352
rect 5686 6296 5691 6352
rect 1853 6294 5691 6296
rect 1853 6291 1919 6294
rect 5625 6291 5691 6294
rect 2497 6218 2563 6221
rect 3233 6218 3299 6221
rect 3693 6218 3759 6221
rect 2497 6216 3066 6218
rect 2497 6160 2502 6216
rect 2558 6160 3066 6216
rect 2497 6158 3066 6160
rect 2497 6155 2563 6158
rect 3006 6082 3066 6158
rect 3233 6216 3759 6218
rect 3233 6160 3238 6216
rect 3294 6160 3698 6216
rect 3754 6160 3759 6216
rect 3233 6158 3759 6160
rect 3233 6155 3299 6158
rect 3693 6155 3759 6158
rect 4153 6218 4219 6221
rect 4429 6218 4495 6221
rect 4153 6216 4495 6218
rect 4153 6160 4158 6216
rect 4214 6160 4434 6216
rect 4490 6160 4495 6216
rect 4153 6158 4495 6160
rect 4153 6155 4219 6158
rect 4429 6155 4495 6158
rect 10409 6218 10475 6221
rect 14000 6218 34000 6248
rect 10409 6216 34000 6218
rect 10409 6160 10414 6216
rect 10470 6160 34000 6216
rect 10409 6158 34000 6160
rect 10409 6155 10475 6158
rect 14000 6128 34000 6158
rect 4797 6082 4863 6085
rect 3006 6080 4863 6082
rect 3006 6024 4802 6080
rect 4858 6024 4863 6080
rect 3006 6022 4863 6024
rect 4797 6019 4863 6022
rect 5717 6082 5783 6085
rect 6821 6082 6887 6085
rect 5717 6080 6887 6082
rect 5717 6024 5722 6080
rect 5778 6024 6826 6080
rect 6882 6024 6887 6080
rect 5717 6022 6887 6024
rect 5717 6019 5783 6022
rect 6821 6019 6887 6022
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 7560 6016 7880 6017
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 5951 7880 5952
rect 3049 5946 3115 5949
rect 4245 5946 4311 5949
rect 3049 5944 4311 5946
rect 3049 5888 3054 5944
rect 3110 5888 4250 5944
rect 4306 5888 4311 5944
rect 3049 5886 4311 5888
rect 3049 5883 3115 5886
rect 4245 5883 4311 5886
rect 4521 5946 4587 5949
rect 7189 5946 7255 5949
rect 4521 5944 7255 5946
rect 4521 5888 4526 5944
rect 4582 5888 7194 5944
rect 7250 5888 7255 5944
rect 4521 5886 7255 5888
rect 4521 5883 4587 5886
rect 7189 5883 7255 5886
rect 1945 5810 2011 5813
rect 4153 5810 4219 5813
rect 1945 5808 4219 5810
rect 1945 5752 1950 5808
rect 2006 5752 4158 5808
rect 4214 5752 4219 5808
rect 1945 5750 4219 5752
rect 1945 5747 2011 5750
rect 4153 5747 4219 5750
rect 6453 5808 6519 5813
rect 6453 5752 6458 5808
rect 6514 5752 6519 5808
rect 6453 5747 6519 5752
rect 13813 5810 13879 5813
rect 14000 5810 34000 5840
rect 13813 5808 34000 5810
rect 13813 5752 13818 5808
rect 13874 5752 34000 5808
rect 13813 5750 34000 5752
rect 13813 5747 13879 5750
rect 2957 5674 3023 5677
rect 3417 5674 3483 5677
rect 2957 5672 3483 5674
rect 2957 5616 2962 5672
rect 3018 5616 3422 5672
rect 3478 5616 3483 5672
rect 2957 5614 3483 5616
rect 6456 5674 6516 5747
rect 14000 5720 34000 5750
rect 8201 5674 8267 5677
rect 6456 5672 8267 5674
rect 6456 5616 8206 5672
rect 8262 5616 8267 5672
rect 6456 5614 8267 5616
rect 2957 5611 3023 5614
rect 3417 5611 3483 5614
rect 8201 5611 8267 5614
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 5407 5380 5408
rect 6637 5402 6703 5405
rect 14000 5402 34000 5432
rect 6637 5400 34000 5402
rect 6637 5344 6642 5400
rect 6698 5344 34000 5400
rect 6637 5342 34000 5344
rect 6637 5339 6703 5342
rect 14000 5312 34000 5342
rect 4061 5266 4127 5269
rect 5809 5266 5875 5269
rect 4061 5264 5875 5266
rect 4061 5208 4066 5264
rect 4122 5208 5814 5264
rect 5870 5208 5875 5264
rect 4061 5206 5875 5208
rect 4061 5203 4127 5206
rect 5809 5203 5875 5206
rect 9673 4994 9739 4997
rect 14000 4994 34000 5024
rect 9673 4992 34000 4994
rect 9673 4936 9678 4992
rect 9734 4936 34000 4992
rect 9673 4934 34000 4936
rect 9673 4931 9739 4934
rect 7560 4928 7880 4929
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 14000 4904 34000 4934
rect 7560 4863 7880 4864
rect 13629 4586 13695 4589
rect 14000 4586 34000 4616
rect 13629 4584 34000 4586
rect 13629 4528 13634 4584
rect 13690 4528 34000 4584
rect 13629 4526 34000 4528
rect 13629 4523 13695 4526
rect 14000 4496 34000 4526
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 4319 5380 4320
rect 4429 4314 4495 4317
rect 4248 4312 4495 4314
rect 4248 4256 4434 4312
rect 4490 4256 4495 4312
rect 4248 4254 4495 4256
rect 4248 4181 4308 4254
rect 4429 4251 4495 4254
rect 4245 4176 4311 4181
rect 4245 4120 4250 4176
rect 4306 4120 4311 4176
rect 4245 4115 4311 4120
rect 7373 4178 7439 4181
rect 13813 4178 13879 4181
rect 14000 4178 34000 4208
rect 7373 4176 8218 4178
rect 7373 4120 7378 4176
rect 7434 4120 8218 4176
rect 7373 4118 8218 4120
rect 7373 4115 7439 4118
rect 7741 4042 7807 4045
rect 2454 4040 7807 4042
rect 2454 3984 7746 4040
rect 7802 3984 7807 4040
rect 2454 3982 7807 3984
rect 2454 3332 2514 3982
rect 7741 3979 7807 3982
rect 7560 3840 7880 3841
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 3775 7880 3776
rect 4705 3770 4771 3773
rect 5441 3770 5507 3773
rect 4705 3768 5507 3770
rect 4705 3712 4710 3768
rect 4766 3712 5446 3768
rect 5502 3712 5507 3768
rect 4705 3710 5507 3712
rect 4705 3707 4771 3710
rect 5441 3707 5507 3710
rect 6453 3770 6519 3773
rect 6729 3770 6795 3773
rect 6453 3768 6795 3770
rect 6453 3712 6458 3768
rect 6514 3712 6734 3768
rect 6790 3712 6795 3768
rect 6453 3710 6795 3712
rect 6453 3707 6519 3710
rect 6729 3707 6795 3710
rect 8158 3637 8218 4118
rect 13813 4176 34000 4178
rect 13813 4120 13818 4176
rect 13874 4120 34000 4176
rect 13813 4118 34000 4120
rect 13813 4115 13879 4118
rect 14000 4088 34000 4118
rect 8753 3770 8819 3773
rect 9213 3770 9279 3773
rect 8753 3768 9279 3770
rect 8753 3712 8758 3768
rect 8814 3712 9218 3768
rect 9274 3712 9279 3768
rect 8753 3710 9279 3712
rect 8753 3707 8819 3710
rect 9213 3707 9279 3710
rect 13813 3770 13879 3773
rect 14000 3770 34000 3800
rect 13813 3768 34000 3770
rect 13813 3712 13818 3768
rect 13874 3712 34000 3768
rect 13813 3710 34000 3712
rect 13813 3707 13879 3710
rect 14000 3680 34000 3710
rect 4981 3634 5047 3637
rect 4524 3632 5047 3634
rect 4524 3576 4986 3632
rect 5042 3576 5047 3632
rect 4524 3574 5047 3576
rect 4524 3365 4584 3574
rect 4981 3571 5047 3574
rect 5441 3634 5507 3637
rect 7833 3634 7899 3637
rect 5441 3632 7899 3634
rect 5441 3576 5446 3632
rect 5502 3576 7838 3632
rect 7894 3576 7899 3632
rect 5441 3574 7899 3576
rect 8158 3632 8267 3637
rect 9673 3634 9739 3637
rect 8158 3576 8206 3632
rect 8262 3576 8267 3632
rect 8158 3574 8267 3576
rect 5441 3571 5507 3574
rect 7833 3571 7899 3574
rect 8201 3571 8267 3574
rect 9630 3632 9739 3634
rect 9630 3576 9678 3632
rect 9734 3576 9739 3632
rect 9630 3571 9739 3576
rect 5165 3498 5231 3501
rect 5165 3496 8770 3498
rect 5165 3440 5170 3496
rect 5226 3440 8770 3496
rect 5165 3438 8770 3440
rect 5165 3435 5231 3438
rect 4521 3360 4587 3365
rect 4521 3304 4526 3360
rect 4582 3304 4587 3360
rect 4521 3299 4587 3304
rect 5717 3362 5783 3365
rect 8109 3362 8175 3365
rect 5717 3360 8175 3362
rect 5717 3304 5722 3360
rect 5778 3304 8114 3360
rect 8170 3304 8175 3360
rect 5717 3302 8175 3304
rect 8710 3362 8770 3438
rect 9213 3362 9279 3365
rect 8710 3360 9279 3362
rect 8710 3304 9218 3360
rect 9274 3304 9279 3360
rect 8710 3302 9279 3304
rect 5717 3299 5783 3302
rect 8109 3299 8175 3302
rect 9213 3299 9279 3302
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 3231 5380 3232
rect 4613 3226 4679 3229
rect 4889 3226 4955 3229
rect 4613 3224 4955 3226
rect 4613 3168 4618 3224
rect 4674 3168 4894 3224
rect 4950 3168 4955 3224
rect 4613 3166 4955 3168
rect 4613 3163 4679 3166
rect 4889 3163 4955 3166
rect 7833 3226 7899 3229
rect 9630 3226 9690 3571
rect 13813 3362 13879 3365
rect 14000 3362 34000 3392
rect 13813 3360 34000 3362
rect 13813 3304 13818 3360
rect 13874 3304 34000 3360
rect 13813 3302 34000 3304
rect 13813 3299 13879 3302
rect 14000 3272 34000 3302
rect 7833 3224 9690 3226
rect 7833 3168 7838 3224
rect 7894 3168 9690 3224
rect 7833 3166 9690 3168
rect 7833 3163 7899 3166
rect 3785 3090 3851 3093
rect 5901 3090 5967 3093
rect 3785 3088 5967 3090
rect 3785 3032 3790 3088
rect 3846 3032 5906 3088
rect 5962 3032 5967 3088
rect 3785 3030 5967 3032
rect 3785 3027 3851 3030
rect 5901 3027 5967 3030
rect 5257 2954 5323 2957
rect 9857 2954 9923 2957
rect 5257 2952 9923 2954
rect 5257 2896 5262 2952
rect 5318 2896 9862 2952
rect 9918 2896 9923 2952
rect 5257 2894 9923 2896
rect 5257 2891 5323 2894
rect 9857 2891 9923 2894
rect 13813 2954 13879 2957
rect 14000 2954 34000 2984
rect 13813 2952 34000 2954
rect 13813 2896 13818 2952
rect 13874 2896 34000 2952
rect 13813 2894 34000 2896
rect 13813 2891 13879 2894
rect 14000 2864 34000 2894
rect 4613 2818 4679 2821
rect 6361 2818 6427 2821
rect 4613 2816 6427 2818
rect 4613 2760 4618 2816
rect 4674 2760 6366 2816
rect 6422 2760 6427 2816
rect 4613 2758 6427 2760
rect 4613 2755 4679 2758
rect 6361 2755 6427 2758
rect 7560 2752 7880 2753
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 2687 7880 2688
rect 4521 2682 4587 2685
rect 5257 2682 5323 2685
rect 4521 2680 5323 2682
rect 4521 2624 4526 2680
rect 4582 2624 5262 2680
rect 5318 2624 5323 2680
rect 4521 2622 5323 2624
rect 4521 2619 4587 2622
rect 5257 2619 5323 2622
rect 4061 2546 4127 2549
rect 5717 2546 5783 2549
rect 4061 2544 5783 2546
rect 4061 2488 4066 2544
rect 4122 2488 5722 2544
rect 5778 2488 5783 2544
rect 4061 2486 5783 2488
rect 4061 2483 4127 2486
rect 5717 2483 5783 2486
rect 8661 2546 8727 2549
rect 8845 2546 8911 2549
rect 8661 2544 8911 2546
rect 8661 2488 8666 2544
rect 8722 2488 8850 2544
rect 8906 2488 8911 2544
rect 8661 2486 8911 2488
rect 8661 2483 8727 2486
rect 8845 2483 8911 2486
rect 14000 2544 34000 2576
rect 14000 2488 16670 2544
rect 16726 2488 34000 2544
rect 14000 2456 34000 2488
rect 3141 2410 3207 2413
rect 7833 2410 7899 2413
rect 3141 2408 7899 2410
rect 3141 2352 3146 2408
rect 3202 2352 7838 2408
rect 7894 2352 7899 2408
rect 3141 2350 7899 2352
rect 3141 2347 3207 2350
rect 7833 2347 7899 2350
rect 8017 2410 8083 2413
rect 13813 2410 13879 2413
rect 8017 2408 13879 2410
rect 8017 2352 8022 2408
rect 8078 2352 13818 2408
rect 13874 2352 13879 2408
rect 8017 2350 13879 2352
rect 8017 2347 8083 2350
rect 13813 2347 13879 2350
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 2143 5380 2144
rect 14000 2136 34000 2168
rect 14000 2080 16578 2136
rect 16634 2080 34000 2136
rect 14000 2048 34000 2080
rect 14000 1728 34000 1760
rect 14000 1672 16578 1728
rect 16634 1672 34000 1728
rect 7560 1664 7880 1665
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 14000 1640 34000 1672
rect 7560 1599 7880 1600
rect 8937 1322 9003 1325
rect 14000 1322 34000 1352
rect 8937 1320 34000 1322
rect 8937 1264 8942 1320
rect 8998 1264 34000 1320
rect 8937 1262 34000 1264
rect 8937 1259 9003 1262
rect 14000 1232 34000 1262
rect 5060 1120 5380 1121
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 5060 1055 5380 1056
rect 9305 914 9371 917
rect 14000 914 34000 944
rect 9305 912 34000 914
rect 9305 856 9310 912
rect 9366 856 34000 912
rect 9305 854 34000 856
rect 9305 851 9371 854
rect 14000 824 34000 854
rect 9121 506 9187 509
rect 14000 506 34000 536
rect 9121 504 34000 506
rect 9121 448 9126 504
rect 9182 448 34000 504
rect 9121 446 34000 448
rect 9121 443 9187 446
rect 14000 416 34000 446
rect 3325 234 3391 237
rect 22093 234 22159 237
rect 3325 232 22159 234
rect 3325 176 3330 232
rect 3386 176 22098 232
rect 22154 176 22159 232
rect 3325 174 22159 176
rect 3325 171 3391 174
rect 22093 171 22159 174
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 5068 1116 5132 1120
rect 5068 1060 5072 1116
rect 5072 1060 5128 1116
rect 5128 1060 5132 1116
rect 5068 1056 5132 1060
rect 5148 1116 5212 1120
rect 5148 1060 5152 1116
rect 5152 1060 5208 1116
rect 5208 1060 5212 1116
rect 5148 1056 5212 1060
rect 5228 1116 5292 1120
rect 5228 1060 5232 1116
rect 5232 1060 5288 1116
rect 5288 1060 5292 1116
rect 5228 1056 5292 1060
rect 5308 1116 5372 1120
rect 5308 1060 5312 1116
rect 5312 1060 5368 1116
rect 5368 1060 5372 1116
rect 5308 1056 5372 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 5060 10912 5380 11472
rect 7560 11456 7880 11472
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 9908 5380 10848
rect 5060 9824 5102 9908
rect 5338 9824 5380 9908
rect 5060 9760 5068 9824
rect 5372 9760 5380 9824
rect 5060 9672 5102 9760
rect 5338 9672 5380 9760
rect 5060 8736 5380 9672
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 6560 5380 7584
rect 5060 6496 5068 6560
rect 5132 6528 5148 6560
rect 5212 6528 5228 6560
rect 5292 6528 5308 6560
rect 5372 6496 5380 6560
rect 5060 6292 5102 6496
rect 5338 6292 5380 6496
rect 5060 5472 5380 6292
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3296 5380 4320
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 3148 5380 3232
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2208 5380 2912
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1120 5380 2144
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 6060 10956 6380 11424
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 1088 6380 3960
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 8218 7880 9216
rect 7560 8192 7602 8218
rect 7838 8192 7880 8218
rect 7560 8128 7568 8192
rect 7872 8128 7880 8192
rect 7560 7982 7602 8128
rect 7838 7982 7880 8128
rect 7560 7104 7880 7982
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 4928 7880 5952
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 4838 7880 4864
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 3840 7880 4602
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1458 7880 1600
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 5060 1040 5380 1056
rect 7560 1040 7880 1222
rect 8560 9266 8880 11424
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 1088 8880 2270
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 5102 9824 5338 9908
rect 5102 9760 5132 9824
rect 5132 9760 5148 9824
rect 5148 9760 5212 9824
rect 5212 9760 5228 9824
rect 5228 9760 5292 9824
rect 5292 9760 5308 9824
rect 5308 9760 5338 9824
rect 5102 9672 5338 9760
rect 5102 6496 5132 6528
rect 5132 6496 5148 6528
rect 5148 6496 5212 6528
rect 5212 6496 5228 6528
rect 5228 6496 5292 6528
rect 5292 6496 5308 6528
rect 5308 6496 5338 6528
rect 5102 6292 5338 6496
rect 5102 2912 5338 3148
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 8192 7838 8218
rect 7602 8128 7632 8192
rect 7632 8128 7648 8192
rect 7648 8128 7712 8192
rect 7712 8128 7728 8192
rect 7728 8128 7792 8192
rect 7792 8128 7808 8192
rect 7808 8128 7838 8192
rect 7602 7982 7838 8128
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 6102 10956
rect 6338 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 5102 9908
rect 5338 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 6102 7576
rect 6338 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 5102 6528
rect 5338 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 5102 3148
rect 5338 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__clkbuf_1  output36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1637331468
transform 1 0 3312 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1637331468
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1637331468
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_26
timestamp 1637331468
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1637331468
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1637331468
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 3312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1637331468
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1637331468
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1637331468
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use gpio_logic_high  gpio_logic_high
timestamp 1637551221
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 3588 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1637331468
transform 1 0 4416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1637331468
transform 1 0 4140 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1637331468
transform 1 0 3864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1637331468
transform 1 0 3588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 5428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_47
timestamp 1637331468
transform 1 0 5244 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_52
timestamp 1637331468
transform 1 0 5704 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 4692 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1637331468
transform 1 0 4968 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1637331468
transform 1 0 4692 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform -1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_31
timestamp 1637331468
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1637331468
transform 1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1637331468
transform 1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1637331468
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1637331468
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1637331468
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1637331468
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1637331468
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50
timestamp 1637331468
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _124_
timestamp 1637331468
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1637331468
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1637331468
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1637331468
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1637331468
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 4324 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1637331468
transform 1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1637331468
transform 1 0 3864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1637331468
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1637331468
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1637331468
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1637331468
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1637331468
transform 1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1637331468
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1637331468
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _208_
timestamp 1637331468
transform 1 0 3588 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__decap_6  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 6348 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 1637331468
transform 1 0 7268 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_65
timestamp 1637331468
transform 1 0 6900 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64
timestamp 1637331468
transform 1 0 6808 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1637331468
transform 1 0 7452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 6992 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1637331468
transform 1 0 7636 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1637331468
transform 1 0 7728 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1637331468
transform 1 0 7636 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72
timestamp 1637331468
transform 1 0 7544 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1637331468
transform 1 0 7912 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76
timestamp 1637331468
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1637331468
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1637331468
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1637331468
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_80
timestamp 1637331468
transform 1 0 8280 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _131_
timestamp 1637331468
transform 1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _130_
timestamp 1637331468
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 7544 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1637331468
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1637331468
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1637331468
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1637331468
transform -1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1637331468
transform 1 0 6532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1637331468
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 6808 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1637331468
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 7544 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 1637331468
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1637331468
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1637331468
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfbbn_1  _205_
timestamp 1637331468
transform 1 0 6532 0 1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__einvp_2  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 7544 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1637331468
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1637331468
transform 1 0 6072 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1637331468
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1637331468
transform 1 0 5980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1637331468
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1637331468
transform 1 0 8648 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1637331468
transform 1 0 8372 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1637331468
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1637331468
transform 1 0 9200 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1637331468
transform 1 0 8740 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90
timestamp 1637331468
transform 1 0 9200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_83
timestamp 1637331468
transform 1 0 8556 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1637331468
transform 1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1637331468
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1637331468
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _183_
timestamp 1637331468
transform 1 0 8740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1637331468
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1637331468
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1637331468
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 8648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1637331468
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1637331468
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _179_
timestamp 1637331468
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1637331468
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1637331468
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1637331468
transform 1 0 8648 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1637331468
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1637331468
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_26
timestamp 1637331468
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1637331468
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 3312 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1637331468
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1637331468
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1637331468
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1637331468
transform 1 0 1196 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1637331468
transform 1 0 1472 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1637331468
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _147_
timestamp 1637331468
transform 1 0 2576 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _128_
timestamp 1637331468
transform 1 0 3036 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1637331468
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _188_
timestamp 1637331468
transform 1 0 1288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _149_
timestamp 1637331468
transform 1 0 1564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _118_
timestamp 1637331468
transform 1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__5
timestamp 1637331468
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 1637331468
transform 1 0 2392 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1637331468
transform 1 0 1196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1637331468
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1637331468
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _215_
timestamp 1637331468
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1637331468
transform 1 0 1196 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1637331468
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _113_
timestamp 1637331468
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _114_
timestamp 1637331468
transform 1 0 3680 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _108_
timestamp 1637331468
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1637331468
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1637331468
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1637331468
transform 1 0 4232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1637331468
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _116_
timestamp 1637331468
transform 1 0 5336 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_7_46
timestamp 1637331468
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _206_
timestamp 1637331468
transform 1 0 5796 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _145_
timestamp 1637331468
transform 1 0 3588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1637331468
transform 1 0 4232 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1637331468
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1637331468
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1637331468
transform 1 0 4968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1637331468
transform 1 0 4232 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1637331468
transform 1 0 5704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1637331468
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _203_
timestamp 1637331468
transform 1 0 3588 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1637331468
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1637331468
transform 1 0 6256 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1637331468
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1637331468
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1637331468
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _120_
timestamp 1637331468
transform 1 0 6164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1637331468
transform 1 0 6808 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp 1637331468
transform 1 0 6716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1637331468
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1637331468
transform 1 0 6164 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1637331468
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _207_
timestamp 1637331468
transform 1 0 6900 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _102_
timestamp 1637331468
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1637331468
transform 1 0 6532 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1637331468
transform 1 0 8832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1637331468
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 8648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1637331468
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1637331468
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1
timestamp 1637331468
transform 1 0 8740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1637331468
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1637331468
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1637331468
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1637331468
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1637331468
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1637331468
transform 1 0 8740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1637331468
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1637331468
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1637331468
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1637331468
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 1288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1637331468
transform 1 0 1196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1637331468
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1637331468
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _202_
timestamp 1637331468
transform 1 0 2576 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__inv_2  _106__4
timestamp 1637331468
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1637331468
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1637331468
transform 1 0 1196 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1637331468
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1637331468
transform 1 0 1288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1637331468
transform 1 0 1564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1637331468
transform 1 0 2300 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1637331468
transform 1 0 1196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1637331468
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__3
timestamp 1637331468
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1637331468
transform 1 0 1288 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1637331468
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1637331468
transform 1 0 1196 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1637331468
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1637331468
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1637331468
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp 1637331468
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1637331468
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1637331468
transform 1 0 1656 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1637331468
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1637331468
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__2
timestamp 1637331468
transform 1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _137_
timestamp 1637331468
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp 1637331468
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _204_
timestamp 1637331468
transform 1 0 2668 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1637331468
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1637331468
transform 1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _107_
timestamp 1637331468
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _151_
timestamp 1637331468
transform 1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1637331468
transform 1 0 3588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1637331468
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _210_
timestamp 1637331468
transform 1 0 5152 0 1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1637331468
transform 1 0 4140 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1637331468
transform 1 0 4140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1637331468
transform 1 0 5336 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1637331468
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1637331468
transform 1 0 5152 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 1637331468
transform 1 0 4876 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 1637331468
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1637331468
transform 1 0 5060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1637331468
transform 1 0 3588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1637331468
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _126_
timestamp 1637331468
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 6164 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1637331468
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1637331468
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1637331468
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1637331468
transform 1 0 6164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1637331468
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1637331468
transform 1 0 5980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1637331468
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _201_
timestamp 1637331468
transform 1 0 7176 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_12  input17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 7176 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1637331468
transform 1 0 6164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _106__1
timestamp 1637331468
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1637331468
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _200_
timestamp 1637331468
transform 1 0 7176 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1637331468
transform 1 0 8648 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1637331468
transform 1 0 8556 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1637331468
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1637331468
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1637331468
transform 1 0 8740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1637331468
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1637331468
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1637331468
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1637331468
transform 1 0 8740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1637331468
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1637331468
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1637331468
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1637331468
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1637331468
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _189_
timestamp 1637331468
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1637331468
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1637331468
transform 1 0 1196 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1637331468
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp 1637331468
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _139_
timestamp 1637331468
transform 1 0 3128 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1637331468
transform 1 0 2392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1637331468
transform 1 0 1288 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1637331468
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1637331468
transform 1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1637331468
transform 1 0 1196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1637331468
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1637331468
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1637331468
transform 1 0 1196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1637331468
transform 1 0 1288 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _174_
timestamp 1637331468
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1637331468
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1637331468
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1637331468
transform 1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1637331468
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp 1637331468
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1637331468
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1637331468
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1637331468
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _199_
timestamp 1637331468
transform 1 0 3680 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1637331468
transform 1 0 3772 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1637331468
transform 1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1637331468
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1637331468
transform 1 0 5612 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1637331468
transform 1 0 4324 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1637331468
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_45
timestamp 1637331468
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1637331468
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 1637331468
transform 1 0 3588 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_18_34
timestamp 1637331468
transform 1 0 4048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1637331468
transform 1 0 4140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1637331468
transform 1 0 4416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_41
timestamp 1637331468
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1637331468
transform 1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1637331468
transform 1 0 5336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1637331468
transform 1 0 5060 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1637331468
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _157_
timestamp 1637331468
transform 1 0 7912 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1637331468
transform 1 0 6072 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1637331468
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _198_
timestamp 1637331468
transform 1 0 6164 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 1637331468
transform 1 0 6164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _163_
timestamp 1637331468
transform 1 0 7636 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1637331468
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1637331468
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1637331468
transform 1 0 8280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1637331468
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_68
timestamp 1637331468
transform 1 0 7176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_63
timestamp 1637331468
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1637331468
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1637331468
transform 1 0 8740 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1637331468
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1637331468
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1637331468
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1637331468
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _181_
timestamp 1637331468
transform 1 0 9016 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1637331468
transform 1 0 8740 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _192_
timestamp 1637331468
transform 1 0 9016 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1637331468
transform 1 0 8556 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1637331468
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1637331468
transform 1 0 9476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_92
timestamp 1637331468
transform 1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1637331468
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1637331468
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 7560 1040 7880 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 8560 1088 8880 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 5060 1040 5380 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 6060 1088 6380 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
