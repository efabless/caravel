magic
tech sky130A
magscale 1 2
timestamp 1666443267
<< checkpaint >>
rect -55820 -1312 -53299 1209
rect -1260 -1260 718860 1038860
<< metal1 >>
rect 676030 897104 676036 897116
rect 663766 897076 676036 897104
rect 652018 896996 652024 897048
rect 652076 897036 652082 897048
rect 663766 897036 663794 897076
rect 676030 897064 676036 897076
rect 676088 897064 676094 897116
rect 652076 897008 663794 897036
rect 652076 896996 652082 897008
rect 654778 895772 654784 895824
rect 654836 895812 654842 895824
rect 675846 895812 675852 895824
rect 654836 895784 675852 895812
rect 654836 895772 654842 895784
rect 675846 895772 675852 895784
rect 675904 895772 675910 895824
rect 672718 895636 672724 895688
rect 672776 895676 672782 895688
rect 676030 895676 676036 895688
rect 672776 895648 676036 895676
rect 672776 895636 672782 895648
rect 676030 895636 676036 895648
rect 676088 895636 676094 895688
rect 672534 894412 672540 894464
rect 672592 894452 672598 894464
rect 675846 894452 675852 894464
rect 672592 894424 675852 894452
rect 672592 894412 672598 894424
rect 675846 894412 675852 894424
rect 675904 894412 675910 894464
rect 673362 894276 673368 894328
rect 673420 894316 673426 894328
rect 676030 894316 676036 894328
rect 673420 894288 676036 894316
rect 673420 894276 673426 894288
rect 676030 894276 676036 894288
rect 676088 894276 676094 894328
rect 671982 892984 671988 893036
rect 672040 893024 672046 893036
rect 676030 893024 676036 893036
rect 672040 892996 676036 893024
rect 672040 892984 672046 892996
rect 676030 892984 676036 892996
rect 676088 892984 676094 893036
rect 670878 892848 670884 892900
rect 670936 892888 670942 892900
rect 675846 892888 675852 892900
rect 670936 892860 675852 892888
rect 670936 892848 670942 892860
rect 675846 892848 675852 892860
rect 675904 892848 675910 892900
rect 674926 890332 674932 890384
rect 674984 890372 674990 890384
rect 676030 890372 676036 890384
rect 674984 890344 676036 890372
rect 674984 890332 674990 890344
rect 676030 890332 676036 890344
rect 676088 890332 676094 890384
rect 676214 890128 676220 890180
rect 676272 890168 676278 890180
rect 676858 890168 676864 890180
rect 676272 890140 676864 890168
rect 676272 890128 676278 890140
rect 676858 890128 676864 890140
rect 676916 890128 676922 890180
rect 674466 888904 674472 888956
rect 674524 888944 674530 888956
rect 676030 888944 676036 888956
rect 674524 888916 676036 888944
rect 674524 888904 674530 888916
rect 676030 888904 676036 888916
rect 676088 888904 676094 888956
rect 676214 888700 676220 888752
rect 676272 888740 676278 888752
rect 677042 888740 677048 888752
rect 676272 888712 677048 888740
rect 676272 888700 676278 888712
rect 677042 888700 677048 888712
rect 677100 888700 677106 888752
rect 674282 887272 674288 887324
rect 674340 887312 674346 887324
rect 676030 887312 676036 887324
rect 674340 887284 676036 887312
rect 674340 887272 674346 887284
rect 676030 887272 676036 887284
rect 676088 887272 676094 887324
rect 673178 886864 673184 886916
rect 673236 886904 673242 886916
rect 676030 886904 676036 886916
rect 673236 886876 676036 886904
rect 673236 886864 673242 886876
rect 676030 886864 676036 886876
rect 676088 886864 676094 886916
rect 671798 885640 671804 885692
rect 671856 885680 671862 885692
rect 676030 885680 676036 885692
rect 671856 885652 676036 885680
rect 671856 885640 671862 885652
rect 676030 885640 676036 885652
rect 676088 885640 676094 885692
rect 653398 880472 653404 880524
rect 653456 880512 653462 880524
rect 675570 880512 675576 880524
rect 653456 880484 675576 880512
rect 653456 880472 653462 880484
rect 675570 880472 675576 880484
rect 675628 880472 675634 880524
rect 675938 880404 675944 880456
rect 675996 880444 676002 880456
rect 679618 880444 679624 880456
rect 675996 880416 679624 880444
rect 675996 880404 676002 880416
rect 679618 880404 679624 880416
rect 679676 880404 679682 880456
rect 675386 879316 675392 879368
rect 675444 879356 675450 879368
rect 676858 879356 676864 879368
rect 675444 879328 676864 879356
rect 675444 879316 675450 879328
rect 676858 879316 676864 879328
rect 676916 879316 676922 879368
rect 675754 879180 675760 879232
rect 675812 879220 675818 879232
rect 678238 879220 678244 879232
rect 675812 879192 678244 879220
rect 675812 879180 675818 879192
rect 678238 879180 678244 879192
rect 678296 879180 678302 879232
rect 675202 879044 675208 879096
rect 675260 879084 675266 879096
rect 676398 879084 676404 879096
rect 675260 879056 676404 879084
rect 675260 879044 675266 879056
rect 676398 879044 676404 879056
rect 676456 879044 676462 879096
rect 674788 878636 674794 878688
rect 674846 878676 674852 878688
rect 677042 878676 677048 878688
rect 674846 878648 677048 878676
rect 674846 878636 674852 878648
rect 677042 878636 677048 878648
rect 677100 878636 677106 878688
rect 675938 878432 675944 878484
rect 675996 878432 676002 878484
rect 675956 878200 675984 878432
rect 675496 878172 675984 878200
rect 675496 877804 675524 878172
rect 675478 877752 675484 877804
rect 675536 877752 675542 877804
rect 675202 874284 675208 874336
rect 675260 874284 675266 874336
rect 675220 874200 675248 874284
rect 675202 874148 675208 874200
rect 675260 874148 675266 874200
rect 675018 874012 675024 874064
rect 675076 874052 675082 874064
rect 675386 874052 675392 874064
rect 675076 874024 675392 874052
rect 675076 874012 675082 874024
rect 675386 874012 675392 874024
rect 675444 874012 675450 874064
rect 674834 873672 674840 873724
rect 674892 873712 674898 873724
rect 675386 873712 675392 873724
rect 674892 873684 675392 873712
rect 674892 873672 674898 873684
rect 675386 873672 675392 873684
rect 675444 873672 675450 873724
rect 657538 869388 657544 869440
rect 657596 869428 657602 869440
rect 675018 869428 675024 869440
rect 657596 869400 675024 869428
rect 657596 869388 657602 869400
rect 675018 869388 675024 869400
rect 675076 869388 675082 869440
rect 674834 869252 674840 869304
rect 674892 869292 674898 869304
rect 675294 869292 675300 869304
rect 674892 869264 675300 869292
rect 674892 869252 674898 869264
rect 675294 869252 675300 869264
rect 675352 869252 675358 869304
rect 651466 868844 651472 868896
rect 651524 868884 651530 868896
rect 654778 868884 654784 868896
rect 651524 868856 654784 868884
rect 651524 868844 651530 868856
rect 654778 868844 654784 868856
rect 654836 868844 654842 868896
rect 654134 868028 654140 868080
rect 654192 868068 654198 868080
rect 675018 868068 675024 868080
rect 654192 868040 675024 868068
rect 654192 868028 654198 868040
rect 675018 868028 675024 868040
rect 675076 868028 675082 868080
rect 674834 867552 674840 867604
rect 674892 867592 674898 867604
rect 675202 867592 675208 867604
rect 674892 867564 675208 867592
rect 674892 867552 674898 867564
rect 675202 867552 675208 867564
rect 675260 867552 675266 867604
rect 651466 866600 651472 866652
rect 651524 866640 651530 866652
rect 672718 866640 672724 866652
rect 651524 866612 672724 866640
rect 651524 866600 651530 866612
rect 672718 866600 672724 866612
rect 672776 866600 672782 866652
rect 651374 865172 651380 865224
rect 651432 865212 651438 865224
rect 653398 865212 653404 865224
rect 651432 865184 653404 865212
rect 651432 865172 651438 865184
rect 653398 865172 653404 865184
rect 653456 865172 653462 865224
rect 651466 863812 651472 863864
rect 651524 863852 651530 863864
rect 657538 863852 657544 863864
rect 651524 863824 657544 863852
rect 651524 863812 651530 863824
rect 657538 863812 657544 863824
rect 657596 863812 657602 863864
rect 651466 862452 651472 862504
rect 651524 862492 651530 862504
rect 654134 862492 654140 862504
rect 651524 862464 654140 862492
rect 651524 862452 651530 862464
rect 654134 862452 654140 862464
rect 654192 862452 654198 862504
rect 35618 817096 35624 817148
rect 35676 817096 35682 817148
rect 35802 817096 35808 817148
rect 35860 817136 35866 817148
rect 46198 817136 46204 817148
rect 35860 817108 46204 817136
rect 35860 817096 35866 817108
rect 46198 817096 46204 817108
rect 46256 817096 46262 817148
rect 35636 817000 35664 817096
rect 61378 817000 61384 817012
rect 35636 816972 61384 817000
rect 61378 816960 61384 816972
rect 61436 816960 61442 817012
rect 35618 815736 35624 815788
rect 35676 815776 35682 815788
rect 44818 815776 44824 815788
rect 35676 815748 44824 815776
rect 35676 815736 35682 815748
rect 44818 815736 44824 815748
rect 44876 815736 44882 815788
rect 35802 815600 35808 815652
rect 35860 815640 35866 815652
rect 45002 815640 45008 815652
rect 35860 815612 45008 815640
rect 35860 815600 35866 815612
rect 45002 815600 45008 815612
rect 45060 815600 45066 815652
rect 35618 814376 35624 814428
rect 35676 814416 35682 814428
rect 44266 814416 44272 814428
rect 35676 814388 44272 814416
rect 35676 814376 35682 814388
rect 44266 814376 44272 814388
rect 44324 814376 44330 814428
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 44542 814280 44548 814292
rect 35860 814252 44548 814280
rect 35860 814240 35866 814252
rect 44542 814240 44548 814252
rect 44600 814240 44606 814292
rect 41322 812812 41328 812864
rect 41380 812852 41386 812864
rect 43254 812852 43260 812864
rect 41380 812824 43260 812852
rect 41380 812812 41386 812824
rect 43254 812812 43260 812824
rect 43312 812812 43318 812864
rect 41138 810704 41144 810756
rect 41196 810744 41202 810756
rect 42518 810744 42524 810756
rect 41196 810716 42524 810744
rect 41196 810704 41202 810716
rect 42518 810704 42524 810716
rect 42576 810704 42582 810756
rect 41138 807440 41144 807492
rect 41196 807480 41202 807492
rect 43070 807480 43076 807492
rect 41196 807452 43076 807480
rect 41196 807440 41202 807452
rect 43070 807440 43076 807452
rect 43128 807440 43134 807492
rect 40954 807304 40960 807356
rect 41012 807344 41018 807356
rect 45186 807344 45192 807356
rect 41012 807316 45192 807344
rect 41012 807304 41018 807316
rect 45186 807304 45192 807316
rect 45244 807304 45250 807356
rect 31754 806624 31760 806676
rect 31812 806664 31818 806676
rect 35618 806664 35624 806676
rect 31812 806636 35624 806664
rect 31812 806624 31818 806636
rect 35618 806624 35624 806636
rect 35676 806624 35682 806676
rect 44818 806556 44824 806608
rect 44876 806596 44882 806608
rect 62758 806596 62764 806608
rect 44876 806568 62764 806596
rect 44876 806556 44882 806568
rect 62758 806556 62764 806568
rect 62816 806556 62822 806608
rect 41322 805944 41328 805996
rect 41380 805984 41386 805996
rect 43806 805984 43812 805996
rect 41380 805956 43812 805984
rect 41380 805944 41386 805956
rect 43806 805944 43812 805956
rect 43864 805944 43870 805996
rect 35618 802544 35624 802596
rect 35676 802584 35682 802596
rect 35676 802556 42380 802584
rect 35676 802544 35682 802556
rect 42352 802460 42380 802556
rect 33042 802408 33048 802460
rect 33100 802448 33106 802460
rect 42150 802448 42156 802460
rect 33100 802420 42156 802448
rect 33100 802408 33106 802420
rect 42150 802408 42156 802420
rect 42208 802408 42214 802460
rect 42334 802408 42340 802460
rect 42392 802408 42398 802460
rect 33778 801184 33784 801236
rect 33836 801224 33842 801236
rect 40126 801224 40132 801236
rect 33836 801196 40132 801224
rect 33836 801184 33842 801196
rect 40126 801184 40132 801196
rect 40184 801184 40190 801236
rect 31018 801048 31024 801100
rect 31076 801088 31082 801100
rect 43622 801088 43628 801100
rect 31076 801060 43628 801088
rect 31076 801048 31082 801060
rect 43622 801048 43628 801060
rect 43680 801048 43686 801100
rect 39298 800844 39304 800896
rect 39356 800884 39362 800896
rect 41966 800884 41972 800896
rect 39356 800856 41972 800884
rect 39356 800844 39362 800856
rect 41966 800844 41972 800856
rect 42024 800844 42030 800896
rect 43438 799008 43444 799060
rect 43496 799048 43502 799060
rect 53098 799048 53104 799060
rect 43496 799020 53104 799048
rect 43496 799008 43502 799020
rect 53098 799008 53104 799020
rect 53156 799008 53162 799060
rect 42518 797648 42524 797700
rect 42576 797688 42582 797700
rect 57238 797688 57244 797700
rect 42576 797660 57244 797688
rect 42576 797648 42582 797660
rect 57238 797648 57244 797660
rect 57296 797648 57302 797700
rect 42886 796492 42892 796544
rect 42944 796532 42950 796544
rect 43622 796532 43628 796544
rect 42944 796504 43628 796532
rect 42944 796492 42950 796504
rect 43622 796492 43628 796504
rect 43680 796492 43686 796544
rect 42426 794996 42432 795048
rect 42484 795036 42490 795048
rect 43070 795036 43076 795048
rect 42484 795008 43076 795036
rect 42484 794996 42490 795008
rect 43070 794996 43076 795008
rect 43128 794996 43134 795048
rect 43070 794860 43076 794912
rect 43128 794900 43134 794912
rect 45186 794900 45192 794912
rect 43128 794872 45192 794900
rect 43128 794860 43134 794872
rect 45186 794860 45192 794872
rect 45244 794860 45250 794912
rect 42426 794044 42432 794096
rect 42484 794084 42490 794096
rect 43070 794084 43076 794096
rect 42484 794056 43076 794084
rect 42484 794044 42490 794056
rect 43070 794044 43076 794056
rect 43128 794044 43134 794096
rect 669222 790916 669228 790968
rect 669280 790956 669286 790968
rect 675202 790956 675208 790968
rect 669280 790928 675208 790956
rect 669280 790916 669286 790928
rect 675202 790916 675208 790928
rect 675260 790916 675266 790968
rect 653398 790780 653404 790832
rect 653456 790820 653462 790832
rect 675386 790820 675392 790832
rect 653456 790792 675392 790820
rect 653456 790780 653462 790792
rect 675386 790780 675392 790792
rect 675444 790780 675450 790832
rect 53098 790712 53104 790764
rect 53156 790752 53162 790764
rect 62206 790752 62212 790764
rect 53156 790724 62212 790752
rect 53156 790712 53162 790724
rect 62206 790712 62212 790724
rect 62264 790712 62270 790764
rect 42242 789692 42248 789744
rect 42300 789692 42306 789744
rect 42260 789540 42288 789692
rect 42242 789488 42248 789540
rect 42300 789488 42306 789540
rect 670602 789352 670608 789404
rect 670660 789392 670666 789404
rect 675110 789392 675116 789404
rect 670660 789364 675116 789392
rect 670660 789352 670666 789364
rect 675110 789352 675116 789364
rect 675168 789352 675174 789404
rect 57238 789148 57244 789200
rect 57296 789188 57302 789200
rect 62114 789188 62120 789200
rect 57296 789160 62120 789188
rect 57296 789148 57302 789160
rect 62114 789148 62120 789160
rect 62172 789148 62178 789200
rect 42610 786632 42616 786684
rect 42668 786672 42674 786684
rect 62114 786672 62120 786684
rect 42668 786644 62120 786672
rect 42668 786632 42674 786644
rect 62114 786632 62120 786644
rect 62172 786632 62178 786684
rect 46198 785136 46204 785188
rect 46256 785176 46262 785188
rect 62114 785176 62120 785188
rect 46256 785148 62120 785176
rect 46256 785136 46262 785148
rect 62114 785136 62120 785148
rect 62172 785136 62178 785188
rect 672994 783844 673000 783896
rect 673052 783884 673058 783896
rect 675110 783884 675116 783896
rect 673052 783856 675116 783884
rect 673052 783844 673058 783856
rect 675110 783844 675116 783856
rect 675168 783844 675174 783896
rect 670418 782484 670424 782536
rect 670476 782524 670482 782536
rect 675294 782524 675300 782536
rect 670476 782496 675300 782524
rect 670476 782484 670482 782496
rect 675294 782484 675300 782496
rect 675352 782484 675358 782536
rect 655514 781056 655520 781108
rect 655572 781096 655578 781108
rect 675018 781096 675024 781108
rect 655572 781068 675024 781096
rect 655572 781056 655578 781068
rect 675018 781056 675024 781068
rect 675076 781056 675082 781108
rect 673546 779968 673552 780020
rect 673604 780008 673610 780020
rect 675110 780008 675116 780020
rect 673604 779980 675116 780008
rect 673604 779968 673610 779980
rect 675110 779968 675116 779980
rect 675168 779968 675174 780020
rect 655146 778472 655152 778524
rect 655204 778512 655210 778524
rect 675018 778512 675024 778524
rect 655204 778484 675024 778512
rect 655204 778472 655210 778484
rect 675018 778472 675024 778484
rect 675076 778472 675082 778524
rect 651466 777588 651472 777640
rect 651524 777628 651530 777640
rect 660298 777628 660304 777640
rect 651524 777600 660304 777628
rect 651524 777588 651530 777600
rect 660298 777588 660304 777600
rect 660356 777588 660362 777640
rect 670234 776976 670240 777028
rect 670292 777016 670298 777028
rect 675018 777016 675024 777028
rect 670292 776988 675024 777016
rect 670292 776976 670298 776988
rect 675018 776976 675024 776988
rect 675076 776976 675082 777028
rect 651466 775684 651472 775736
rect 651524 775724 651530 775736
rect 669958 775724 669964 775736
rect 651524 775696 669964 775724
rect 651524 775684 651530 775696
rect 669958 775684 669964 775696
rect 670016 775684 670022 775736
rect 668394 775548 668400 775600
rect 668452 775588 668458 775600
rect 675018 775588 675024 775600
rect 668452 775560 675024 775588
rect 668452 775548 668458 775560
rect 675018 775548 675024 775560
rect 675076 775548 675082 775600
rect 651374 775276 651380 775328
rect 651432 775316 651438 775328
rect 653398 775316 653404 775328
rect 651432 775288 653404 775316
rect 651432 775276 651438 775288
rect 653398 775276 653404 775288
rect 653456 775276 653462 775328
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 41690 774228 41696 774240
rect 35860 774200 41696 774228
rect 35860 774188 35866 774200
rect 41690 774188 41696 774200
rect 41748 774188 41754 774240
rect 42058 774188 42064 774240
rect 42116 774228 42122 774240
rect 59998 774228 60004 774240
rect 42116 774200 60004 774228
rect 42116 774188 42122 774200
rect 59998 774188 60004 774200
rect 60056 774188 60062 774240
rect 651466 774120 651472 774172
rect 651524 774160 651530 774172
rect 655514 774160 655520 774172
rect 651524 774132 655520 774160
rect 651524 774120 651530 774132
rect 655514 774120 655520 774132
rect 655572 774120 655578 774172
rect 651466 773780 651472 773832
rect 651524 773820 651530 773832
rect 655146 773820 655152 773832
rect 651524 773792 655152 773820
rect 651524 773780 651530 773792
rect 655146 773780 655152 773792
rect 655204 773780 655210 773832
rect 35802 773372 35808 773424
rect 35860 773412 35866 773424
rect 40494 773412 40500 773424
rect 35860 773384 40500 773412
rect 35860 773372 35866 773384
rect 40494 773372 40500 773384
rect 40552 773372 40558 773424
rect 36004 773180 38654 773208
rect 35526 773100 35532 773152
rect 35584 773140 35590 773152
rect 36004 773140 36032 773180
rect 35584 773112 36032 773140
rect 38626 773140 38654 773180
rect 40494 773140 40500 773152
rect 38626 773112 40500 773140
rect 35584 773100 35590 773112
rect 40494 773100 40500 773112
rect 40552 773100 40558 773152
rect 40696 773044 41414 773072
rect 35342 772964 35348 773016
rect 35400 773004 35406 773016
rect 40696 773004 40724 773044
rect 35400 772976 40724 773004
rect 41386 773004 41414 773044
rect 41690 773004 41696 773016
rect 41386 772976 41696 773004
rect 35400 772964 35406 772976
rect 41690 772964 41696 772976
rect 41748 772964 41754 773016
rect 42058 772964 42064 773016
rect 42116 773004 42122 773016
rect 46198 773004 46204 773016
rect 42116 772976 46204 773004
rect 42116 772964 42122 772976
rect 46198 772964 46204 772976
rect 46256 772964 46262 773016
rect 35158 772828 35164 772880
rect 35216 772868 35222 772880
rect 61378 772868 61384 772880
rect 35216 772840 41736 772868
rect 35216 772828 35222 772840
rect 41708 772744 41736 772840
rect 42076 772840 61384 772868
rect 42076 772744 42104 772840
rect 61378 772828 61384 772840
rect 61436 772828 61442 772880
rect 41690 772692 41696 772744
rect 41748 772692 41754 772744
rect 42058 772692 42064 772744
rect 42116 772692 42122 772744
rect 35802 771808 35808 771860
rect 35860 771848 35866 771860
rect 39574 771848 39580 771860
rect 35860 771820 39580 771848
rect 35860 771808 35866 771820
rect 39574 771808 39580 771820
rect 39632 771808 39638 771860
rect 41322 771644 41328 771656
rect 36004 771616 41328 771644
rect 35618 771536 35624 771588
rect 35676 771576 35682 771588
rect 36004 771576 36032 771616
rect 41322 771604 41328 771616
rect 41380 771604 41386 771656
rect 35676 771548 36032 771576
rect 35676 771536 35682 771548
rect 42058 771468 42064 771520
rect 42116 771508 42122 771520
rect 44542 771508 44548 771520
rect 42116 771480 44548 771508
rect 42116 771468 42122 771480
rect 44542 771468 44548 771480
rect 44600 771468 44606 771520
rect 35802 771400 35808 771452
rect 35860 771440 35866 771452
rect 41690 771440 41696 771452
rect 35860 771412 41696 771440
rect 35860 771400 35866 771412
rect 41690 771400 41696 771412
rect 41748 771400 41754 771452
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 40034 770488 40040 770500
rect 35860 770460 40040 770488
rect 35860 770448 35866 770460
rect 40034 770448 40040 770460
rect 40092 770448 40098 770500
rect 35618 770176 35624 770228
rect 35676 770216 35682 770228
rect 40310 770216 40316 770228
rect 35676 770188 40316 770216
rect 35676 770176 35682 770188
rect 40310 770176 40316 770188
rect 40368 770176 40374 770228
rect 35802 770040 35808 770092
rect 35860 770080 35866 770092
rect 41690 770080 41696 770092
rect 35860 770052 41696 770080
rect 35860 770040 35866 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 42058 770040 42064 770092
rect 42116 770080 42122 770092
rect 44266 770080 44272 770092
rect 42116 770052 44272 770080
rect 42116 770040 42122 770052
rect 44266 770040 44272 770052
rect 44324 770040 44330 770092
rect 35802 768952 35808 769004
rect 35860 768992 35866 769004
rect 39758 768992 39764 769004
rect 35860 768964 39764 768992
rect 35860 768952 35866 768964
rect 39758 768952 39764 768964
rect 39816 768952 39822 769004
rect 35526 768816 35532 768868
rect 35584 768856 35590 768868
rect 40678 768856 40684 768868
rect 35584 768828 40684 768856
rect 35584 768816 35590 768828
rect 40678 768816 40684 768828
rect 40736 768816 40742 768868
rect 35342 768680 35348 768732
rect 35400 768720 35406 768732
rect 41690 768720 41696 768732
rect 35400 768692 41696 768720
rect 35400 768680 35406 768692
rect 41690 768680 41696 768692
rect 41748 768680 41754 768732
rect 35802 767456 35808 767508
rect 35860 767496 35866 767508
rect 36538 767496 36544 767508
rect 35860 767468 36544 767496
rect 35860 767456 35866 767468
rect 36538 767456 36544 767468
rect 36596 767456 36602 767508
rect 39040 767400 40080 767428
rect 35618 767320 35624 767372
rect 35676 767360 35682 767372
rect 39040 767360 39068 767400
rect 35676 767332 39068 767360
rect 35676 767320 35682 767332
rect 40052 767292 40080 767400
rect 41690 767292 41696 767304
rect 40052 767264 41696 767292
rect 41690 767252 41696 767264
rect 41748 767252 41754 767304
rect 35802 766028 35808 766080
rect 35860 766068 35866 766080
rect 39298 766068 39304 766080
rect 35860 766040 39304 766068
rect 35860 766028 35866 766040
rect 39298 766028 39304 766040
rect 39356 766028 39362 766080
rect 35802 764804 35808 764856
rect 35860 764844 35866 764856
rect 40402 764844 40408 764856
rect 35860 764816 40408 764844
rect 35860 764804 35866 764816
rect 40402 764804 40408 764816
rect 40460 764804 40466 764856
rect 35802 764532 35808 764584
rect 35860 764572 35866 764584
rect 41690 764572 41696 764584
rect 35860 764544 41696 764572
rect 35860 764532 35866 764544
rect 41690 764532 41696 764544
rect 41748 764532 41754 764584
rect 37090 763648 37096 763700
rect 37148 763688 37154 763700
rect 39298 763688 39304 763700
rect 37148 763660 39304 763688
rect 37148 763648 37154 763660
rect 39298 763648 39304 763660
rect 39356 763648 39362 763700
rect 35802 763240 35808 763292
rect 35860 763280 35866 763292
rect 41690 763280 41696 763292
rect 35860 763252 41696 763280
rect 35860 763240 35866 763252
rect 41690 763240 41696 763252
rect 41748 763240 41754 763292
rect 35802 761880 35808 761932
rect 35860 761920 35866 761932
rect 39942 761920 39948 761932
rect 35860 761892 39948 761920
rect 35860 761880 35866 761892
rect 39942 761880 39948 761892
rect 40000 761880 40006 761932
rect 33042 760996 33048 761048
rect 33100 761036 33106 761048
rect 41506 761036 41512 761048
rect 33100 761008 41512 761036
rect 33100 760996 33106 761008
rect 41506 760996 41512 761008
rect 41564 760996 41570 761048
rect 35158 759568 35164 759620
rect 35216 759608 35222 759620
rect 35216 759580 38654 759608
rect 35216 759568 35222 759580
rect 38626 759540 38654 759580
rect 40494 759540 40500 759552
rect 38626 759512 40500 759540
rect 40494 759500 40500 759512
rect 40552 759500 40558 759552
rect 39298 757732 39304 757784
rect 39356 757772 39362 757784
rect 41598 757772 41604 757784
rect 39356 757744 41604 757772
rect 39356 757732 39362 757744
rect 41598 757732 41604 757744
rect 41656 757732 41662 757784
rect 44726 755488 44732 755540
rect 44784 755528 44790 755540
rect 62758 755528 62764 755540
rect 44784 755500 62764 755528
rect 44784 755488 44790 755500
rect 62758 755488 62764 755500
rect 62816 755488 62822 755540
rect 43438 754876 43444 754928
rect 43496 754916 43502 754928
rect 45094 754916 45100 754928
rect 43496 754888 45100 754916
rect 43496 754876 43502 754888
rect 45094 754876 45100 754888
rect 45152 754876 45158 754928
rect 42334 753924 42340 753976
rect 42392 753964 42398 753976
rect 43622 753964 43628 753976
rect 42392 753936 43628 753964
rect 42392 753924 42398 753936
rect 43622 753924 43628 753936
rect 43680 753924 43686 753976
rect 42242 753516 42248 753568
rect 42300 753556 42306 753568
rect 45278 753556 45284 753568
rect 42300 753528 45284 753556
rect 42300 753516 42306 753528
rect 45278 753516 45284 753528
rect 45336 753516 45342 753568
rect 61378 746988 61384 747040
rect 61436 747028 61442 747040
rect 62390 747028 62396 747040
rect 61436 747000 62396 747028
rect 61436 746988 61442 747000
rect 62390 746988 62396 747000
rect 62448 746988 62454 747040
rect 45094 746512 45100 746564
rect 45152 746552 45158 746564
rect 62114 746552 62120 746564
rect 45152 746524 62120 746552
rect 45152 746512 45158 746524
rect 62114 746512 62120 746524
rect 62172 746512 62178 746564
rect 671062 745220 671068 745272
rect 671120 745260 671126 745272
rect 675110 745260 675116 745272
rect 671120 745232 675116 745260
rect 671120 745220 671126 745232
rect 675110 745220 675116 745232
rect 675168 745220 675174 745272
rect 42518 743996 42524 744048
rect 42576 744036 42582 744048
rect 42576 744008 45554 744036
rect 42576 743996 42582 744008
rect 45526 743900 45554 744008
rect 62114 743900 62120 743912
rect 45526 743872 62120 743900
rect 62114 743860 62120 743872
rect 62172 743860 62178 743912
rect 46198 743724 46204 743776
rect 46256 743764 46262 743776
rect 62114 743764 62120 743776
rect 46256 743736 62120 743764
rect 46256 743724 46262 743736
rect 62114 743724 62120 743736
rect 62172 743724 62178 743776
rect 671338 743724 671344 743776
rect 671396 743764 671402 743776
rect 675478 743764 675484 743776
rect 671396 743736 675484 743764
rect 671396 743724 671402 743736
rect 675478 743724 675484 743736
rect 675536 743724 675542 743776
rect 672350 742432 672356 742484
rect 672408 742472 672414 742484
rect 675386 742472 675392 742484
rect 672408 742444 675392 742472
rect 672408 742432 672414 742444
rect 675386 742432 675392 742444
rect 675444 742432 675450 742484
rect 59998 742364 60004 742416
rect 60056 742404 60062 742416
rect 62114 742404 62120 742416
rect 60056 742376 62120 742404
rect 60056 742364 60062 742376
rect 62114 742364 62120 742376
rect 62172 742364 62178 742416
rect 668762 741072 668768 741124
rect 668820 741112 668826 741124
rect 675294 741112 675300 741124
rect 668820 741084 675300 741112
rect 668820 741072 668826 741084
rect 675294 741072 675300 741084
rect 675352 741072 675358 741124
rect 669774 739916 669780 739968
rect 669832 739956 669838 739968
rect 675386 739956 675392 739968
rect 669832 739928 675392 739956
rect 669832 739916 669838 739928
rect 675386 739916 675392 739928
rect 675444 739916 675450 739968
rect 652018 736176 652024 736228
rect 652076 736216 652082 736228
rect 653398 736216 653404 736228
rect 652076 736188 653404 736216
rect 652076 736176 652082 736188
rect 653398 736176 653404 736188
rect 653456 736176 653462 736228
rect 672166 735740 672172 735752
rect 663766 735712 672172 735740
rect 657538 735564 657544 735616
rect 657596 735604 657602 735616
rect 663766 735604 663794 735712
rect 672166 735700 672172 735712
rect 672224 735700 672230 735752
rect 657596 735576 663794 735604
rect 657596 735564 657602 735576
rect 672166 734544 672172 734596
rect 672224 734584 672230 734596
rect 675294 734584 675300 734596
rect 672224 734556 675300 734584
rect 672224 734544 672230 734556
rect 675294 734544 675300 734556
rect 675352 734544 675358 734596
rect 669590 734408 669596 734460
rect 669648 734448 669654 734460
rect 675110 734448 675116 734460
rect 669648 734420 675116 734448
rect 669648 734408 669654 734420
rect 675110 734408 675116 734420
rect 675168 734408 675174 734460
rect 675110 734312 675116 734324
rect 663766 734284 675116 734312
rect 654778 734136 654784 734188
rect 654836 734176 654842 734188
rect 663766 734176 663794 734284
rect 675110 734272 675116 734284
rect 675168 734272 675174 734324
rect 654836 734148 663794 734176
rect 654836 734136 654842 734148
rect 651466 733388 651472 733440
rect 651524 733428 651530 733440
rect 668578 733428 668584 733440
rect 651524 733400 668584 733428
rect 651524 733388 651530 733400
rect 668578 733388 668584 733400
rect 668636 733388 668642 733440
rect 651466 732776 651472 732828
rect 651524 732816 651530 732828
rect 661678 732816 661684 732828
rect 651524 732788 661684 732816
rect 651524 732776 651530 732788
rect 661678 732776 661684 732788
rect 661736 732776 661742 732828
rect 674466 731824 674472 731876
rect 674524 731864 674530 731876
rect 675294 731864 675300 731876
rect 674524 731836 675300 731864
rect 674524 731824 674530 731836
rect 675294 731824 675300 731836
rect 675352 731824 675358 731876
rect 651466 731416 651472 731468
rect 651524 731456 651530 731468
rect 658918 731456 658924 731468
rect 651524 731428 658924 731456
rect 651524 731416 651530 731428
rect 658918 731416 658924 731428
rect 658976 731416 658982 731468
rect 651466 731280 651472 731332
rect 651524 731320 651530 731332
rect 671338 731320 671344 731332
rect 651524 731292 671344 731320
rect 651524 731280 651530 731292
rect 671338 731280 671344 731292
rect 671396 731280 671402 731332
rect 42058 731144 42064 731196
rect 42116 731184 42122 731196
rect 61378 731184 61384 731196
rect 42116 731156 61384 731184
rect 42116 731144 42122 731156
rect 61378 731144 61384 731156
rect 61436 731144 61442 731196
rect 35802 731076 35808 731128
rect 35860 731116 35866 731128
rect 41690 731116 41696 731128
rect 35860 731088 41696 731116
rect 35860 731076 35866 731088
rect 41690 731076 41696 731088
rect 41748 731076 41754 731128
rect 674834 731076 674840 731128
rect 674892 731076 674898 731128
rect 674852 730912 674880 731076
rect 675202 730912 675208 730924
rect 674852 730884 675208 730912
rect 675202 730872 675208 730884
rect 675260 730872 675266 730924
rect 35802 730532 35808 730584
rect 35860 730572 35866 730584
rect 39942 730572 39948 730584
rect 35860 730544 39948 730572
rect 35860 730532 35866 730544
rect 39942 730532 39948 730544
rect 40000 730532 40006 730584
rect 674834 730464 674840 730516
rect 674892 730504 674898 730516
rect 675294 730504 675300 730516
rect 674892 730476 675300 730504
rect 674892 730464 674898 730476
rect 675294 730464 675300 730476
rect 675352 730464 675358 730516
rect 35618 730260 35624 730312
rect 35676 730300 35682 730312
rect 41690 730300 41696 730312
rect 35676 730272 41696 730300
rect 35676 730260 35682 730272
rect 41690 730260 41696 730272
rect 41748 730260 41754 730312
rect 671246 730056 671252 730108
rect 671304 730096 671310 730108
rect 675294 730096 675300 730108
rect 671304 730068 675300 730096
rect 671304 730056 671310 730068
rect 675294 730056 675300 730068
rect 675352 730056 675358 730108
rect 651466 729988 651472 730040
rect 651524 730028 651530 730040
rect 657538 730028 657544 730040
rect 651524 730000 657544 730028
rect 651524 729988 651530 730000
rect 657538 729988 657544 730000
rect 657596 729988 657602 730040
rect 35434 729376 35440 729428
rect 35492 729416 35498 729428
rect 41690 729416 41696 729428
rect 35492 729388 41696 729416
rect 35492 729376 35498 729388
rect 41690 729376 41696 729388
rect 41748 729376 41754 729428
rect 42058 729308 42064 729360
rect 42116 729348 42122 729360
rect 62758 729348 62764 729360
rect 42116 729320 62764 729348
rect 42116 729308 42122 729320
rect 62758 729308 62764 729320
rect 62816 729308 62822 729360
rect 35802 729036 35808 729088
rect 35860 729076 35866 729088
rect 41690 729076 41696 729088
rect 35860 729048 41696 729076
rect 35860 729036 35866 729048
rect 41690 729036 41696 729048
rect 41748 729036 41754 729088
rect 35618 728764 35624 728816
rect 35676 728804 35682 728816
rect 39574 728804 39580 728816
rect 35676 728776 39580 728804
rect 35676 728764 35682 728776
rect 39574 728764 39580 728776
rect 39632 728764 39638 728816
rect 35250 728628 35256 728680
rect 35308 728668 35314 728680
rect 41690 728668 41696 728680
rect 35308 728640 41696 728668
rect 35308 728628 35314 728640
rect 41690 728628 41696 728640
rect 41748 728628 41754 728680
rect 42058 728628 42064 728680
rect 42116 728668 42122 728680
rect 43070 728668 43076 728680
rect 42116 728640 43076 728668
rect 42116 728628 42122 728640
rect 43070 728628 43076 728640
rect 43128 728628 43134 728680
rect 672718 728628 672724 728680
rect 672776 728668 672782 728680
rect 675294 728668 675300 728680
rect 672776 728640 675300 728668
rect 672776 728628 672782 728640
rect 675294 728628 675300 728640
rect 675352 728628 675358 728680
rect 651466 728492 651472 728544
rect 651524 728532 651530 728544
rect 654778 728532 654784 728544
rect 651524 728504 654784 728532
rect 651524 728492 651530 728504
rect 654778 728492 654784 728504
rect 654836 728492 654842 728544
rect 671798 728288 671804 728340
rect 671856 728328 671862 728340
rect 671856 728300 674176 728328
rect 671856 728288 671862 728300
rect 673178 728084 673184 728136
rect 673236 728124 673242 728136
rect 673236 728096 674058 728124
rect 673236 728084 673242 728096
rect 42058 727880 42064 727932
rect 42116 727920 42122 727932
rect 44266 727920 44272 727932
rect 42116 727892 44272 727920
rect 42116 727880 42122 727892
rect 44266 727880 44272 727892
rect 44324 727880 44330 727932
rect 675846 727880 675852 727932
rect 675904 727920 675910 727932
rect 683298 727920 683304 727932
rect 675904 727892 683304 727920
rect 675904 727880 675910 727892
rect 683298 727880 683304 727892
rect 683356 727880 683362 727932
rect 35802 727812 35808 727864
rect 35860 727852 35866 727864
rect 41506 727852 41512 727864
rect 35860 727824 41512 727852
rect 35860 727812 35866 727824
rect 41506 727812 41512 727824
rect 41564 727812 41570 727864
rect 35618 727540 35624 727592
rect 35676 727580 35682 727592
rect 40402 727580 40408 727592
rect 35676 727552 40408 727580
rect 35676 727540 35682 727552
rect 40402 727540 40408 727552
rect 40460 727540 40466 727592
rect 35802 727404 35808 727456
rect 35860 727444 35866 727456
rect 41690 727444 41696 727456
rect 35860 727416 41696 727444
rect 35860 727404 35866 727416
rect 41690 727404 41696 727416
rect 41748 727404 41754 727456
rect 35802 727268 35808 727320
rect 35860 727308 35866 727320
rect 41690 727308 41696 727320
rect 35860 727280 41696 727308
rect 35860 727268 35866 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 45002 727308 45008 727320
rect 42116 727280 45008 727308
rect 42116 727268 42122 727280
rect 45002 727268 45008 727280
rect 45060 727268 45066 727320
rect 676030 726520 676036 726572
rect 676088 726560 676094 726572
rect 683482 726560 683488 726572
rect 676088 726532 683488 726560
rect 676088 726520 676094 726532
rect 683482 726520 683488 726532
rect 683540 726520 683546 726572
rect 41322 726180 41328 726232
rect 41380 726220 41386 726232
rect 41690 726220 41696 726232
rect 41380 726192 41696 726220
rect 41380 726180 41386 726192
rect 41690 726180 41696 726192
rect 41748 726180 41754 726232
rect 41138 725908 41144 725960
rect 41196 725948 41202 725960
rect 41598 725948 41604 725960
rect 41196 725920 41604 725948
rect 41196 725908 41202 725920
rect 41598 725908 41604 725920
rect 41656 725908 41662 725960
rect 674374 721692 674380 721744
rect 674432 721692 674438 721744
rect 675110 721692 675116 721744
rect 675168 721692 675174 721744
rect 674392 721268 674420 721692
rect 675128 721268 675156 721692
rect 674374 721216 674380 721268
rect 674432 721216 674438 721268
rect 675110 721216 675116 721268
rect 675168 721216 675174 721268
rect 674374 720808 674380 720860
rect 674432 720808 674438 720860
rect 675110 720808 675116 720860
rect 675168 720808 675174 720860
rect 674392 720520 674420 720808
rect 674374 720468 674380 720520
rect 674432 720468 674438 720520
rect 675128 720508 675156 720808
rect 675386 720508 675392 720520
rect 675128 720480 675392 720508
rect 675386 720468 675392 720480
rect 675444 720468 675450 720520
rect 653398 716252 653404 716304
rect 653456 716292 653462 716304
rect 674006 716292 674012 716304
rect 653456 716264 674012 716292
rect 653456 716252 653462 716264
rect 674006 716252 674012 716264
rect 674064 716252 674070 716304
rect 35158 715776 35164 715828
rect 35216 715816 35222 715828
rect 41690 715816 41696 715828
rect 35216 715788 41696 715816
rect 35216 715776 35222 715788
rect 41690 715776 41696 715788
rect 41748 715776 41754 715828
rect 669958 715708 669964 715760
rect 670016 715748 670022 715760
rect 673270 715748 673276 715760
rect 670016 715720 673276 715748
rect 670016 715708 670022 715720
rect 673270 715708 673276 715720
rect 673328 715708 673334 715760
rect 33778 715640 33784 715692
rect 33836 715680 33842 715692
rect 37734 715680 37740 715692
rect 33836 715652 37740 715680
rect 33836 715640 33842 715652
rect 37734 715640 37740 715652
rect 37792 715640 37798 715692
rect 33042 715504 33048 715556
rect 33100 715544 33106 715556
rect 39850 715544 39856 715556
rect 33100 715516 39856 715544
rect 33100 715504 33106 715516
rect 39850 715504 39856 715516
rect 39908 715504 39914 715556
rect 674006 714932 674012 714944
rect 663766 714904 674012 714932
rect 660298 714824 660304 714876
rect 660356 714864 660362 714876
rect 663766 714864 663794 714904
rect 674006 714892 674012 714904
rect 674064 714892 674070 714944
rect 660356 714836 663794 714864
rect 660356 714824 660362 714836
rect 670878 713668 670884 713720
rect 670936 713708 670942 713720
rect 674006 713708 674012 713720
rect 670936 713680 674012 713708
rect 670936 713668 670942 713680
rect 674006 713668 674012 713680
rect 674064 713668 674070 713720
rect 671338 713192 671344 713244
rect 671396 713232 671402 713244
rect 674006 713232 674012 713244
rect 671396 713204 674012 713232
rect 671396 713192 671402 713204
rect 674006 713192 674012 713204
rect 674064 713192 674070 713244
rect 671982 712376 671988 712428
rect 672040 712416 672046 712428
rect 674006 712416 674012 712428
rect 672040 712388 674012 712416
rect 672040 712376 672046 712388
rect 674006 712376 674012 712388
rect 674064 712376 674070 712428
rect 43622 712104 43628 712156
rect 43680 712144 43686 712156
rect 50338 712144 50344 712156
rect 43680 712116 50344 712144
rect 43680 712104 43686 712116
rect 50338 712104 50344 712116
rect 50396 712104 50402 712156
rect 42242 711696 42248 711748
rect 42300 711696 42306 711748
rect 42260 711136 42288 711696
rect 42242 711084 42248 711136
rect 42300 711084 42306 711136
rect 669222 710676 669228 710728
rect 669280 710716 669286 710728
rect 674006 710716 674012 710728
rect 669280 710688 674012 710716
rect 669280 710676 669286 710688
rect 674006 710676 674012 710688
rect 674064 710676 674070 710728
rect 670418 710404 670424 710456
rect 670476 710444 670482 710456
rect 674006 710444 674012 710456
rect 670476 710416 674012 710444
rect 670476 710404 670482 710416
rect 674006 710404 674012 710416
rect 674064 710404 674070 710456
rect 668394 709996 668400 710048
rect 668452 710036 668458 710048
rect 674006 710036 674012 710048
rect 668452 710008 674012 710036
rect 668452 709996 668458 710008
rect 674006 709996 674012 710008
rect 674064 709996 674070 710048
rect 670602 709588 670608 709640
rect 670660 709628 670666 709640
rect 674006 709628 674012 709640
rect 670660 709600 674012 709628
rect 670660 709588 670666 709600
rect 674006 709588 674012 709600
rect 674064 709588 674070 709640
rect 43622 709316 43628 709368
rect 43680 709356 43686 709368
rect 44450 709356 44456 709368
rect 43680 709328 44456 709356
rect 43680 709316 43686 709328
rect 44450 709316 44456 709328
rect 44508 709316 44514 709368
rect 42242 709180 42248 709232
rect 42300 709220 42306 709232
rect 44634 709220 44640 709232
rect 42300 709192 44640 709220
rect 42300 709180 42306 709192
rect 44634 709180 44640 709192
rect 44692 709180 44698 709232
rect 671614 707956 671620 708008
rect 671672 707996 671678 708008
rect 674006 707996 674012 708008
rect 671672 707968 674012 707996
rect 671672 707956 671678 707968
rect 674006 707956 674012 707968
rect 674064 707956 674070 708008
rect 42610 707412 42616 707464
rect 42668 707412 42674 707464
rect 42426 707072 42432 707124
rect 42484 707072 42490 707124
rect 42444 706648 42472 707072
rect 42628 706716 42656 707412
rect 42610 706664 42616 706716
rect 42668 706664 42674 706716
rect 42426 706596 42432 706648
rect 42484 706596 42490 706648
rect 670234 705304 670240 705356
rect 670292 705344 670298 705356
rect 674006 705344 674012 705356
rect 670292 705316 674012 705344
rect 670292 705304 670298 705316
rect 674006 705304 674012 705316
rect 674064 705304 674070 705356
rect 675846 705168 675852 705220
rect 675904 705208 675910 705220
rect 683114 705208 683120 705220
rect 675904 705180 683120 705208
rect 675904 705168 675910 705180
rect 683114 705168 683120 705180
rect 683172 705168 683178 705220
rect 50338 705100 50344 705152
rect 50396 705140 50402 705152
rect 62114 705140 62120 705152
rect 50396 705112 62120 705140
rect 50396 705100 50402 705112
rect 62114 705100 62120 705112
rect 62172 705100 62178 705152
rect 670602 703808 670608 703860
rect 670660 703848 670666 703860
rect 674006 703848 674012 703860
rect 670660 703820 674012 703848
rect 670660 703808 670666 703820
rect 674006 703808 674012 703820
rect 674064 703808 674070 703860
rect 44450 703740 44456 703792
rect 44508 703780 44514 703792
rect 62114 703780 62120 703792
rect 44508 703752 62120 703780
rect 44508 703740 44514 703752
rect 62114 703740 62120 703752
rect 62172 703740 62178 703792
rect 42702 701020 42708 701072
rect 42760 701060 42766 701072
rect 62206 701060 62212 701072
rect 42760 701032 62212 701060
rect 42760 701020 42766 701032
rect 62206 701020 62212 701032
rect 62264 701020 62270 701072
rect 654778 701020 654784 701072
rect 654836 701060 654842 701072
rect 673546 701060 673552 701072
rect 654836 701032 673552 701060
rect 654836 701020 654842 701032
rect 673546 701020 673552 701032
rect 673604 701020 673610 701072
rect 46198 698164 46204 698216
rect 46256 698204 46262 698216
rect 62114 698204 62120 698216
rect 46256 698176 62120 698204
rect 46256 698164 46262 698176
rect 62114 698164 62120 698176
rect 62172 698164 62178 698216
rect 666462 697076 666468 697128
rect 666520 697116 666526 697128
rect 673546 697116 673552 697128
rect 666520 697088 673552 697116
rect 666520 697076 666526 697088
rect 673546 697076 673552 697088
rect 673604 697076 673610 697128
rect 656802 690004 656808 690056
rect 656860 690044 656866 690056
rect 673546 690044 673552 690056
rect 656860 690016 673552 690044
rect 656860 690004 656866 690016
rect 673546 690004 673552 690016
rect 673604 690004 673610 690056
rect 674282 690004 674288 690056
rect 674340 690044 674346 690056
rect 675110 690044 675116 690056
rect 674340 690016 675116 690044
rect 674340 690004 674346 690016
rect 675110 690004 675116 690016
rect 675168 690004 675174 690056
rect 652754 688780 652760 688832
rect 652812 688820 652818 688832
rect 673546 688820 673552 688832
rect 652812 688792 673552 688820
rect 652812 688780 652818 688792
rect 673546 688780 673552 688792
rect 673604 688780 673610 688832
rect 651650 688644 651656 688696
rect 651708 688684 651714 688696
rect 660298 688684 660304 688696
rect 651708 688656 660304 688684
rect 651708 688644 651714 688656
rect 660298 688644 660304 688656
rect 660356 688644 660362 688696
rect 651466 687896 651472 687948
rect 651524 687936 651530 687948
rect 667198 687936 667204 687948
rect 651524 687908 667204 687936
rect 651524 687896 651530 687908
rect 667198 687896 667204 687908
rect 667256 687896 667262 687948
rect 42702 687284 42708 687336
rect 42760 687324 42766 687336
rect 42760 687296 51074 687324
rect 42760 687284 42766 687296
rect 51046 687256 51074 687296
rect 61378 687256 61384 687268
rect 51046 687228 61384 687256
rect 61378 687216 61384 687228
rect 61436 687216 61442 687268
rect 674466 687216 674472 687268
rect 674524 687256 674530 687268
rect 675110 687256 675116 687268
rect 674524 687228 675116 687256
rect 674524 687216 674530 687228
rect 675110 687216 675116 687228
rect 675168 687216 675174 687268
rect 651466 687148 651472 687200
rect 651524 687188 651530 687200
rect 654778 687188 654784 687200
rect 651524 687160 654784 687188
rect 651524 687148 651530 687160
rect 654778 687148 654784 687160
rect 654836 687148 654842 687200
rect 43438 686468 43444 686520
rect 43496 686508 43502 686520
rect 62758 686508 62764 686520
rect 43496 686480 62764 686508
rect 43496 686468 43502 686480
rect 62758 686468 62764 686480
rect 62816 686468 62822 686520
rect 41138 685992 41144 686044
rect 41196 686032 41202 686044
rect 41690 686032 41696 686044
rect 41196 686004 41696 686032
rect 41196 685992 41202 686004
rect 41690 685992 41696 686004
rect 41748 685992 41754 686044
rect 42058 685992 42064 686044
rect 42116 686032 42122 686044
rect 44634 686032 44640 686044
rect 42116 686004 44640 686032
rect 42116 685992 42122 686004
rect 44634 685992 44640 686004
rect 44692 685992 44698 686044
rect 670234 685924 670240 685976
rect 670292 685964 670298 685976
rect 673178 685964 673184 685976
rect 670292 685936 673184 685964
rect 670292 685924 670298 685936
rect 673178 685924 673184 685936
rect 673236 685924 673242 685976
rect 40862 685856 40868 685908
rect 40920 685896 40926 685908
rect 41690 685896 41696 685908
rect 40920 685868 41696 685896
rect 40920 685856 40926 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 45186 685896 45192 685908
rect 42116 685868 45192 685896
rect 42116 685856 42122 685868
rect 45186 685856 45192 685868
rect 45244 685856 45250 685908
rect 651466 685516 651472 685568
rect 651524 685556 651530 685568
rect 656802 685556 656808 685568
rect 651524 685528 656808 685556
rect 651524 685516 651530 685528
rect 656802 685516 656808 685528
rect 656860 685516 656866 685568
rect 41046 684700 41052 684752
rect 41104 684740 41110 684752
rect 41690 684740 41696 684752
rect 41104 684712 41696 684740
rect 41104 684700 41110 684712
rect 41690 684700 41696 684712
rect 41748 684700 41754 684752
rect 40862 684564 40868 684616
rect 40920 684604 40926 684616
rect 40920 684576 41414 684604
rect 40920 684564 40926 684576
rect 41386 684536 41414 684576
rect 41690 684536 41696 684548
rect 41386 684508 41696 684536
rect 41690 684496 41696 684508
rect 41748 684496 41754 684548
rect 42058 684496 42064 684548
rect 42116 684536 42122 684548
rect 45186 684536 45192 684548
rect 42116 684508 45192 684536
rect 42116 684496 42122 684508
rect 45186 684496 45192 684508
rect 45244 684496 45250 684548
rect 41322 683408 41328 683460
rect 41380 683448 41386 683460
rect 41690 683448 41696 683460
rect 41380 683420 41696 683448
rect 41380 683408 41386 683420
rect 41690 683408 41696 683420
rect 41748 683408 41754 683460
rect 675846 682524 675852 682576
rect 675904 682564 675910 682576
rect 683206 682564 683212 682576
rect 675904 682536 683212 682564
rect 675904 682524 675910 682536
rect 683206 682524 683212 682536
rect 683264 682524 683270 682576
rect 683390 682428 683396 682440
rect 675864 682400 683396 682428
rect 675864 682304 675892 682400
rect 683390 682388 683396 682400
rect 683448 682388 683454 682440
rect 675846 682252 675852 682304
rect 675904 682252 675910 682304
rect 40954 679124 40960 679176
rect 41012 679164 41018 679176
rect 41322 679164 41328 679176
rect 41012 679136 41328 679164
rect 41012 679124 41018 679136
rect 41322 679124 41328 679136
rect 41380 679124 41386 679176
rect 41138 678988 41144 679040
rect 41196 679028 41202 679040
rect 41690 679028 41696 679040
rect 41196 679000 41696 679028
rect 41196 678988 41202 679000
rect 41690 678988 41696 679000
rect 41748 678988 41754 679040
rect 42058 678988 42064 679040
rect 42116 679028 42122 679040
rect 45002 679028 45008 679040
rect 42116 679000 45008 679028
rect 42116 678988 42122 679000
rect 45002 678988 45008 679000
rect 45060 678988 45066 679040
rect 40954 677696 40960 677748
rect 41012 677736 41018 677748
rect 41598 677736 41604 677748
rect 41012 677708 41604 677736
rect 41012 677696 41018 677708
rect 41598 677696 41604 677708
rect 41656 677696 41662 677748
rect 35158 672868 35164 672920
rect 35216 672908 35222 672920
rect 38930 672908 38936 672920
rect 35216 672880 38936 672908
rect 35216 672868 35222 672880
rect 38930 672868 38936 672880
rect 38988 672868 38994 672920
rect 33778 672732 33784 672784
rect 33836 672772 33842 672784
rect 38194 672772 38200 672784
rect 33836 672744 38200 672772
rect 33836 672732 33842 672744
rect 38194 672732 38200 672744
rect 38252 672732 38258 672784
rect 668578 671100 668584 671152
rect 668636 671140 668642 671152
rect 674006 671140 674012 671152
rect 668636 671112 674012 671140
rect 668636 671100 668642 671112
rect 674006 671100 674012 671112
rect 674064 671100 674070 671152
rect 661678 670692 661684 670744
rect 661736 670732 661742 670744
rect 673638 670732 673644 670744
rect 661736 670704 673644 670732
rect 661736 670692 661742 670704
rect 673638 670692 673644 670704
rect 673696 670692 673702 670744
rect 671798 670080 671804 670132
rect 671856 670120 671862 670132
rect 674006 670120 674012 670132
rect 671856 670092 674012 670120
rect 671856 670080 671862 670092
rect 674006 670080 674012 670092
rect 674064 670080 674070 670132
rect 658918 669468 658924 669520
rect 658976 669508 658982 669520
rect 673638 669508 673644 669520
rect 658976 669480 673644 669508
rect 658976 669468 658982 669480
rect 673638 669468 673644 669480
rect 673696 669468 673702 669520
rect 45370 669332 45376 669384
rect 45428 669372 45434 669384
rect 53098 669372 53104 669384
rect 45428 669344 53104 669372
rect 45428 669332 45434 669344
rect 53098 669332 53104 669344
rect 53156 669332 53162 669384
rect 670418 669332 670424 669384
rect 670476 669372 670482 669384
rect 674006 669372 674012 669384
rect 670476 669344 674012 669372
rect 670476 669332 670482 669344
rect 674006 669332 674012 669344
rect 674064 669332 674070 669384
rect 670970 669196 670976 669248
rect 671028 669236 671034 669248
rect 671798 669236 671804 669248
rect 671028 669208 671804 669236
rect 671028 669196 671034 669208
rect 671798 669196 671804 669208
rect 671856 669196 671862 669248
rect 671338 668516 671344 668568
rect 671396 668556 671402 668568
rect 674006 668556 674012 668568
rect 671396 668528 674012 668556
rect 671396 668516 671402 668528
rect 674006 668516 674012 668528
rect 674064 668516 674070 668568
rect 671614 668176 671620 668228
rect 671672 668216 671678 668228
rect 673638 668216 673644 668228
rect 671672 668188 673644 668216
rect 671672 668176 671678 668188
rect 673638 668176 673644 668188
rect 673696 668176 673702 668228
rect 45738 667904 45744 667956
rect 45796 667944 45802 667956
rect 57238 667944 57244 667956
rect 45796 667916 57244 667944
rect 45796 667904 45802 667916
rect 57238 667904 57244 667916
rect 57296 667904 57302 667956
rect 671338 667904 671344 667956
rect 671396 667944 671402 667956
rect 674006 667944 674012 667956
rect 671396 667916 674012 667944
rect 671396 667904 671402 667916
rect 674006 667904 674012 667916
rect 674064 667904 674070 667956
rect 42242 667428 42248 667480
rect 42300 667468 42306 667480
rect 45370 667468 45376 667480
rect 42300 667440 45376 667468
rect 42300 667428 42306 667440
rect 45370 667428 45376 667440
rect 45428 667428 45434 667480
rect 671982 666884 671988 666936
rect 672040 666924 672046 666936
rect 674006 666924 674012 666936
rect 672040 666896 674012 666924
rect 672040 666884 672046 666896
rect 674006 666884 674012 666896
rect 674064 666884 674070 666936
rect 670970 666544 670976 666596
rect 671028 666584 671034 666596
rect 673638 666584 673644 666596
rect 671028 666556 673644 666584
rect 671028 666544 671034 666556
rect 673638 666544 673644 666556
rect 673696 666544 673702 666596
rect 669774 665592 669780 665644
rect 669832 665632 669838 665644
rect 674006 665632 674012 665644
rect 669832 665604 674012 665632
rect 669832 665592 669838 665604
rect 674006 665592 674012 665604
rect 674064 665592 674070 665644
rect 671798 665252 671804 665304
rect 671856 665292 671862 665304
rect 673638 665292 673644 665304
rect 671856 665264 673644 665292
rect 671856 665252 671862 665264
rect 673638 665252 673644 665264
rect 673696 665252 673702 665304
rect 672350 665116 672356 665168
rect 672408 665156 672414 665168
rect 673362 665156 673368 665168
rect 672408 665128 673368 665156
rect 672408 665116 672414 665128
rect 673362 665116 673368 665128
rect 673420 665116 673426 665168
rect 42242 664844 42248 664896
rect 42300 664884 42306 664896
rect 43990 664884 43996 664896
rect 42300 664856 43996 664884
rect 42300 664844 42306 664856
rect 43990 664844 43996 664856
rect 44048 664844 44054 664896
rect 42242 664164 42248 664216
rect 42300 664204 42306 664216
rect 42702 664204 42708 664216
rect 42300 664176 42708 664204
rect 42300 664164 42306 664176
rect 42702 664164 42708 664176
rect 42760 664164 42766 664216
rect 42242 663008 42248 663060
rect 42300 663048 42306 663060
rect 43622 663048 43628 663060
rect 42300 663020 43628 663048
rect 42300 663008 42306 663020
rect 43622 663008 43628 663020
rect 43680 663008 43686 663060
rect 668762 662940 668768 662992
rect 668820 662980 668826 662992
rect 674006 662980 674012 662992
rect 668820 662952 674012 662980
rect 668820 662940 668826 662952
rect 674006 662940 674012 662952
rect 674064 662940 674070 662992
rect 669590 662532 669596 662584
rect 669648 662572 669654 662584
rect 674006 662572 674012 662584
rect 669648 662544 674012 662572
rect 669648 662532 669654 662544
rect 674006 662532 674012 662544
rect 674064 662532 674070 662584
rect 669038 661580 669044 661632
rect 669096 661620 669102 661632
rect 674006 661620 674012 661632
rect 669096 661592 674012 661620
rect 669096 661580 669102 661592
rect 674006 661580 674012 661592
rect 674064 661580 674070 661632
rect 667842 661104 667848 661156
rect 667900 661144 667906 661156
rect 674006 661144 674012 661156
rect 667900 661116 674012 661144
rect 667900 661104 667906 661116
rect 674006 661104 674012 661116
rect 674064 661104 674070 661156
rect 53098 660900 53104 660952
rect 53156 660940 53162 660952
rect 62114 660940 62120 660952
rect 53156 660912 62120 660940
rect 53156 660900 53162 660912
rect 62114 660900 62120 660912
rect 62172 660900 62178 660952
rect 671154 660084 671160 660136
rect 671212 660124 671218 660136
rect 674006 660124 674012 660136
rect 671212 660096 674012 660124
rect 671212 660084 671218 660096
rect 674006 660084 674012 660096
rect 674064 660084 674070 660136
rect 675846 659812 675852 659864
rect 675904 659852 675910 659864
rect 683114 659852 683120 659864
rect 675904 659824 683120 659852
rect 675904 659812 675910 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 57238 659540 57244 659592
rect 57296 659580 57302 659592
rect 62114 659580 62120 659592
rect 57296 659552 62120 659580
rect 57296 659540 57302 659552
rect 62114 659540 62120 659552
rect 62172 659540 62178 659592
rect 42518 657500 42524 657552
rect 42576 657540 42582 657552
rect 62114 657540 62120 657552
rect 42576 657512 62120 657540
rect 42576 657500 42582 657512
rect 62114 657500 62120 657512
rect 62172 657500 62178 657552
rect 42058 657364 42064 657416
rect 42116 657404 42122 657416
rect 42702 657404 42708 657416
rect 42116 657376 42708 657404
rect 42116 657364 42122 657376
rect 42702 657364 42708 657376
rect 42760 657364 42766 657416
rect 653398 655528 653404 655580
rect 653456 655568 653462 655580
rect 674006 655568 674012 655580
rect 653456 655540 674012 655568
rect 653456 655528 653462 655540
rect 674006 655528 674012 655540
rect 674064 655528 674070 655580
rect 44818 655460 44824 655512
rect 44876 655500 44882 655512
rect 62114 655500 62120 655512
rect 44876 655472 62120 655500
rect 44876 655460 44882 655472
rect 62114 655460 62120 655472
rect 62172 655460 62178 655512
rect 668210 654100 668216 654152
rect 668268 654140 668274 654152
rect 674006 654140 674012 654152
rect 668268 654112 674012 654140
rect 668268 654100 668274 654112
rect 674006 654100 674012 654112
rect 674064 654100 674070 654152
rect 667382 647232 667388 647284
rect 667440 647272 667446 647284
rect 674006 647272 674012 647284
rect 667440 647244 674012 647272
rect 667440 647232 667446 647244
rect 674006 647232 674012 647244
rect 674064 647232 674070 647284
rect 655514 645872 655520 645924
rect 655572 645912 655578 645924
rect 671154 645912 671160 645924
rect 655572 645884 671160 645912
rect 655572 645872 655578 645884
rect 671154 645872 671160 645884
rect 671212 645872 671218 645924
rect 674926 645192 674932 645244
rect 674984 645232 674990 645244
rect 675294 645232 675300 645244
rect 674984 645204 675300 645232
rect 674984 645192 674990 645204
rect 675294 645192 675300 645204
rect 675352 645192 675358 645244
rect 652018 645124 652024 645176
rect 652076 645164 652082 645176
rect 668578 645164 668584 645176
rect 652076 645136 668584 645164
rect 652076 645124 652082 645136
rect 668578 645124 668584 645136
rect 668636 645124 668642 645176
rect 35802 644444 35808 644496
rect 35860 644484 35866 644496
rect 41690 644484 41696 644496
rect 35860 644456 41696 644484
rect 35860 644444 35866 644456
rect 41690 644444 41696 644456
rect 41748 644444 41754 644496
rect 42058 644444 42064 644496
rect 42116 644484 42122 644496
rect 59998 644484 60004 644496
rect 42116 644456 60004 644484
rect 42116 644444 42122 644456
rect 59998 644444 60004 644456
rect 60056 644444 60062 644496
rect 674558 643628 674564 643680
rect 674616 643628 674622 643680
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 39942 643532 39948 643544
rect 35860 643504 39948 643532
rect 35860 643492 35866 643504
rect 39942 643492 39948 643504
rect 40000 643492 40006 643544
rect 674576 643340 674604 643628
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 44634 643328 44640 643340
rect 42116 643300 44640 643328
rect 42116 643288 42122 643300
rect 44634 643288 44640 643300
rect 44692 643288 44698 643340
rect 674558 643288 674564 643340
rect 674616 643288 674622 643340
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 675110 643220 675116 643272
rect 675168 643220 675174 643272
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 61378 643124 61384 643136
rect 42116 643096 61384 643124
rect 42116 643084 42122 643096
rect 61378 643084 61384 643096
rect 61436 643084 61442 643136
rect 655330 643084 655336 643136
rect 655388 643124 655394 643136
rect 674006 643124 674012 643136
rect 655388 643096 674012 643124
rect 655388 643084 655394 643096
rect 674006 643084 674012 643096
rect 674064 643084 674070 643136
rect 674466 643084 674472 643136
rect 674524 643124 674530 643136
rect 675128 643124 675156 643220
rect 674524 643096 675156 643124
rect 674524 643084 674530 643096
rect 38562 642472 38568 642524
rect 38620 642512 38626 642524
rect 41690 642512 41696 642524
rect 38620 642484 41696 642512
rect 38620 642472 38626 642484
rect 41690 642472 41696 642484
rect 41748 642472 41754 642524
rect 42058 642336 42064 642388
rect 42116 642376 42122 642388
rect 62758 642376 62764 642388
rect 42116 642348 62764 642376
rect 42116 642336 42122 642348
rect 62758 642336 62764 642348
rect 62816 642336 62822 642388
rect 651466 642336 651472 642388
rect 651524 642376 651530 642388
rect 658918 642376 658924 642388
rect 651524 642348 658924 642376
rect 651524 642336 651530 642348
rect 658918 642336 658924 642348
rect 658976 642336 658982 642388
rect 35618 641996 35624 642048
rect 35676 642036 35682 642048
rect 40126 642036 40132 642048
rect 35676 642008 40132 642036
rect 35676 641996 35682 642008
rect 40126 641996 40132 642008
rect 40184 641996 40190 642048
rect 35802 641724 35808 641776
rect 35860 641764 35866 641776
rect 41690 641764 41696 641776
rect 35860 641736 41696 641764
rect 35860 641724 35866 641736
rect 41690 641724 41696 641736
rect 41748 641724 41754 641776
rect 42058 641724 42064 641776
rect 42116 641764 42122 641776
rect 45186 641764 45192 641776
rect 42116 641736 45192 641764
rect 42116 641724 42122 641736
rect 45186 641724 45192 641736
rect 45244 641724 45250 641776
rect 35802 640704 35808 640756
rect 35860 640744 35866 640756
rect 39758 640744 39764 640756
rect 35860 640716 39764 640744
rect 35860 640704 35866 640716
rect 39758 640704 39764 640716
rect 39816 640704 39822 640756
rect 35434 640432 35440 640484
rect 35492 640472 35498 640484
rect 40034 640472 40040 640484
rect 35492 640444 40040 640472
rect 35492 640432 35498 640444
rect 40034 640432 40040 640444
rect 40092 640432 40098 640484
rect 35618 640296 35624 640348
rect 35676 640336 35682 640348
rect 41690 640336 41696 640348
rect 35676 640308 41696 640336
rect 35676 640296 35682 640308
rect 41690 640296 41696 640308
rect 41748 640296 41754 640348
rect 42058 640296 42064 640348
rect 42116 640336 42122 640348
rect 45278 640336 45284 640348
rect 42116 640308 45284 640336
rect 42116 640296 42122 640308
rect 45278 640296 45284 640308
rect 45336 640296 45342 640348
rect 651466 640296 651472 640348
rect 651524 640336 651530 640348
rect 669958 640336 669964 640348
rect 651524 640308 669964 640336
rect 651524 640296 651530 640308
rect 669958 640296 669964 640308
rect 670016 640296 670022 640348
rect 651374 640092 651380 640144
rect 651432 640132 651438 640144
rect 653398 640132 653404 640144
rect 651432 640104 653404 640132
rect 651432 640092 651438 640104
rect 653398 640092 653404 640104
rect 653456 640092 653462 640144
rect 35802 639140 35808 639192
rect 35860 639180 35866 639192
rect 35860 639140 35894 639180
rect 35866 639112 35894 639140
rect 37918 639112 37924 639124
rect 35866 639084 37924 639112
rect 37918 639072 37924 639084
rect 37976 639072 37982 639124
rect 39132 639016 40080 639044
rect 35802 638936 35808 638988
rect 35860 638976 35866 638988
rect 39132 638976 39160 639016
rect 35860 638948 39160 638976
rect 35860 638936 35866 638948
rect 40052 638908 40080 639016
rect 41414 638908 41420 638920
rect 40052 638880 41420 638908
rect 41414 638868 41420 638880
rect 41472 638868 41478 638920
rect 651650 638868 651656 638920
rect 651708 638908 651714 638920
rect 655330 638908 655336 638920
rect 651708 638880 655336 638908
rect 651708 638868 651714 638880
rect 655330 638868 655336 638880
rect 655388 638868 655394 638920
rect 651466 638732 651472 638784
rect 651524 638772 651530 638784
rect 655514 638772 655520 638784
rect 651524 638744 655520 638772
rect 651524 638732 651530 638744
rect 655514 638732 655520 638744
rect 655572 638732 655578 638784
rect 35802 637712 35808 637764
rect 35860 637752 35866 637764
rect 36538 637752 36544 637764
rect 35860 637724 36544 637752
rect 35860 637712 35866 637724
rect 36538 637712 36544 637724
rect 36596 637712 36602 637764
rect 674558 636964 674564 637016
rect 674616 637004 674622 637016
rect 675478 637004 675484 637016
rect 674616 636976 675484 637004
rect 674616 636964 674622 636976
rect 675478 636964 675484 636976
rect 675536 636964 675542 637016
rect 35618 636896 35624 636948
rect 35676 636936 35682 636948
rect 40678 636936 40684 636948
rect 35676 636908 40684 636936
rect 35676 636896 35682 636908
rect 40678 636896 40684 636908
rect 40736 636896 40742 636948
rect 675846 636828 675852 636880
rect 675904 636868 675910 636880
rect 683390 636868 683396 636880
rect 675904 636840 683396 636868
rect 675904 636828 675910 636840
rect 683390 636828 683396 636840
rect 683448 636828 683454 636880
rect 35526 636488 35532 636540
rect 35584 636528 35590 636540
rect 35584 636500 36032 636528
rect 35584 636488 35590 636500
rect 36004 636460 36032 636500
rect 39850 636460 39856 636472
rect 36004 636432 39856 636460
rect 39850 636420 39856 636432
rect 39908 636420 39914 636472
rect 35802 636216 35808 636268
rect 35860 636256 35866 636268
rect 41690 636256 41696 636268
rect 35860 636228 41696 636256
rect 35860 636216 35866 636228
rect 41690 636216 41696 636228
rect 41748 636216 41754 636268
rect 42058 636216 42064 636268
rect 42116 636256 42122 636268
rect 44542 636256 44548 636268
rect 42116 636228 44548 636256
rect 42116 636216 42122 636228
rect 44542 636216 44548 636228
rect 44600 636216 44606 636268
rect 35802 634924 35808 634976
rect 35860 634964 35866 634976
rect 41598 634964 41604 634976
rect 35860 634936 41604 634964
rect 35860 634924 35866 634936
rect 41598 634924 41604 634936
rect 41656 634924 41662 634976
rect 35802 633700 35808 633752
rect 35860 633740 35866 633752
rect 35860 633712 36032 633740
rect 35860 633700 35866 633712
rect 36004 633672 36032 633712
rect 39574 633672 39580 633684
rect 36004 633644 39580 633672
rect 39574 633632 39580 633644
rect 39632 633632 39638 633684
rect 35618 633428 35624 633480
rect 35676 633468 35682 633480
rect 40126 633468 40132 633480
rect 35676 633440 40132 633468
rect 35676 633428 35682 633440
rect 40126 633428 40132 633440
rect 40184 633428 40190 633480
rect 674926 631796 674932 631848
rect 674984 631836 674990 631848
rect 675478 631836 675484 631848
rect 674984 631808 675484 631836
rect 674984 631796 674990 631808
rect 675478 631796 675484 631808
rect 675536 631796 675542 631848
rect 36538 630708 36544 630760
rect 36596 630748 36602 630760
rect 41598 630748 41604 630760
rect 36596 630720 41604 630748
rect 36596 630708 36602 630720
rect 41598 630708 41604 630720
rect 41656 630708 41662 630760
rect 31938 629892 31944 629944
rect 31996 629932 32002 629944
rect 40218 629932 40224 629944
rect 31996 629904 40224 629932
rect 31996 629892 32002 629904
rect 40218 629892 40224 629904
rect 40276 629892 40282 629944
rect 38562 628260 38568 628312
rect 38620 628300 38626 628312
rect 40494 628300 40500 628312
rect 38620 628272 40500 628300
rect 38620 628260 38626 628272
rect 40494 628260 40500 628272
rect 40552 628260 40558 628312
rect 44174 625812 44180 625864
rect 44232 625852 44238 625864
rect 62942 625852 62948 625864
rect 44232 625824 62948 625852
rect 44232 625812 44238 625824
rect 62942 625812 62948 625824
rect 63000 625812 63006 625864
rect 667198 625812 667204 625864
rect 667256 625852 667262 625864
rect 674006 625852 674012 625864
rect 667256 625824 674012 625852
rect 667256 625812 667262 625824
rect 674006 625812 674012 625824
rect 674064 625812 674070 625864
rect 668578 625540 668584 625592
rect 668636 625580 668642 625592
rect 674006 625580 674012 625592
rect 668636 625552 674012 625580
rect 668636 625540 668642 625552
rect 674006 625540 674012 625552
rect 674064 625540 674070 625592
rect 42242 625336 42248 625388
rect 42300 625376 42306 625388
rect 42518 625376 42524 625388
rect 42300 625348 42524 625376
rect 42300 625336 42306 625348
rect 42518 625336 42524 625348
rect 42576 625336 42582 625388
rect 673454 625240 673460 625252
rect 663766 625212 673460 625240
rect 660298 625132 660304 625184
rect 660356 625172 660362 625184
rect 663766 625172 663794 625212
rect 673454 625200 673460 625212
rect 673512 625200 673518 625252
rect 660356 625144 663794 625172
rect 660356 625132 660362 625144
rect 42518 625064 42524 625116
rect 42576 625104 42582 625116
rect 42702 625104 42708 625116
rect 42576 625076 42708 625104
rect 42576 625064 42582 625076
rect 42702 625064 42708 625076
rect 42760 625064 42766 625116
rect 670418 625064 670424 625116
rect 670476 625104 670482 625116
rect 674006 625104 674012 625116
rect 670476 625076 674012 625104
rect 670476 625064 670482 625076
rect 674006 625064 674012 625076
rect 674064 625064 674070 625116
rect 671154 624656 671160 624708
rect 671212 624696 671218 624708
rect 674006 624696 674012 624708
rect 671212 624668 674012 624696
rect 671212 624656 671218 624668
rect 674006 624656 674012 624668
rect 674064 624656 674070 624708
rect 42334 624384 42340 624436
rect 42392 624424 42398 624436
rect 44174 624424 44180 624436
rect 42392 624396 44180 624424
rect 42392 624384 42398 624396
rect 44174 624384 44180 624396
rect 44232 624384 44238 624436
rect 671614 624316 671620 624368
rect 671672 624356 671678 624368
rect 674006 624356 674012 624368
rect 671672 624328 674012 624356
rect 671672 624316 671678 624328
rect 674006 624316 674012 624328
rect 674064 624316 674070 624368
rect 42242 624044 42248 624096
rect 42300 624084 42306 624096
rect 44450 624084 44456 624096
rect 42300 624056 44456 624084
rect 42300 624044 42306 624056
rect 44450 624044 44456 624056
rect 44508 624044 44514 624096
rect 671614 623840 671620 623892
rect 671672 623880 671678 623892
rect 674006 623880 674012 623892
rect 671672 623852 674012 623880
rect 671672 623840 671678 623852
rect 674006 623840 674012 623852
rect 674064 623840 674070 623892
rect 671338 623500 671344 623552
rect 671396 623540 671402 623552
rect 674006 623540 674012 623552
rect 671396 623512 674012 623540
rect 671396 623500 671402 623512
rect 674006 623500 674012 623512
rect 674064 623500 674070 623552
rect 669590 623024 669596 623076
rect 669648 623064 669654 623076
rect 674006 623064 674012 623076
rect 669648 623036 674012 623064
rect 669648 623024 669654 623036
rect 674006 623024 674012 623036
rect 674064 623024 674070 623076
rect 675846 623024 675852 623076
rect 675904 623064 675910 623076
rect 683114 623064 683120 623076
rect 675904 623036 683120 623064
rect 675904 623024 675910 623036
rect 683114 623024 683120 623036
rect 683172 623024 683178 623076
rect 670970 622684 670976 622736
rect 671028 622724 671034 622736
rect 674006 622724 674012 622736
rect 671028 622696 674012 622724
rect 671028 622684 671034 622696
rect 674006 622684 674012 622696
rect 674064 622684 674070 622736
rect 669774 622208 669780 622260
rect 669832 622248 669838 622260
rect 674006 622248 674012 622260
rect 669832 622220 674012 622248
rect 669832 622208 669838 622220
rect 674006 622208 674012 622220
rect 674064 622208 674070 622260
rect 669406 621188 669412 621240
rect 669464 621228 669470 621240
rect 674006 621228 674012 621240
rect 669464 621200 674012 621228
rect 669464 621188 669470 621200
rect 674006 621188 674012 621200
rect 674064 621188 674070 621240
rect 672166 620576 672172 620628
rect 672224 620616 672230 620628
rect 673086 620616 673092 620628
rect 672224 620588 673092 620616
rect 672224 620576 672230 620588
rect 673086 620576 673092 620588
rect 673144 620576 673150 620628
rect 670234 619828 670240 619880
rect 670292 619868 670298 619880
rect 673086 619868 673092 619880
rect 670292 619840 673092 619868
rect 670292 619828 670298 619840
rect 673086 619828 673092 619840
rect 673144 619828 673150 619880
rect 42242 619624 42248 619676
rect 42300 619664 42306 619676
rect 44358 619664 44364 619676
rect 42300 619636 44364 619664
rect 42300 619624 42306 619636
rect 44358 619624 44364 619636
rect 44416 619624 44422 619676
rect 666462 619624 666468 619676
rect 666520 619664 666526 619676
rect 673454 619664 673460 619676
rect 666520 619636 673460 619664
rect 666520 619624 666526 619636
rect 673454 619624 673460 619636
rect 673512 619624 673518 619676
rect 669222 619012 669228 619064
rect 669280 619052 669286 619064
rect 673454 619052 673460 619064
rect 669280 619024 673460 619052
rect 669280 619012 669286 619024
rect 673454 619012 673460 619024
rect 673512 619012 673518 619064
rect 44174 616768 44180 616820
rect 44232 616808 44238 616820
rect 62114 616808 62120 616820
rect 44232 616780 62120 616808
rect 44232 616768 44238 616780
rect 62114 616768 62120 616780
rect 62172 616768 62178 616820
rect 670786 616564 670792 616616
rect 670844 616604 670850 616616
rect 673454 616604 673460 616616
rect 670844 616576 673460 616604
rect 670844 616564 670850 616576
rect 673454 616564 673460 616576
rect 673512 616564 673518 616616
rect 675846 615476 675852 615528
rect 675904 615516 675910 615528
rect 683114 615516 683120 615528
rect 675904 615488 683120 615516
rect 675904 615476 675910 615488
rect 683114 615476 683120 615488
rect 683172 615476 683178 615528
rect 43070 615408 43076 615460
rect 43128 615448 43134 615460
rect 44082 615448 44088 615460
rect 43128 615420 44088 615448
rect 43128 615408 43134 615420
rect 44082 615408 44088 615420
rect 44140 615408 44146 615460
rect 669406 614864 669412 614916
rect 669464 614904 669470 614916
rect 673454 614904 673460 614916
rect 669464 614876 673460 614904
rect 669464 614864 669470 614876
rect 673454 614864 673460 614876
rect 673512 614864 673518 614916
rect 42610 614116 42616 614168
rect 42668 614156 42674 614168
rect 62114 614156 62120 614168
rect 42668 614128 62120 614156
rect 42668 614116 42674 614128
rect 62114 614116 62120 614128
rect 62172 614116 62178 614168
rect 59998 612620 60004 612672
rect 60056 612660 60062 612672
rect 62114 612660 62120 612672
rect 60056 612632 62120 612660
rect 60056 612620 60062 612632
rect 62114 612620 62120 612632
rect 62172 612620 62178 612672
rect 43806 612592 43812 612604
rect 43548 612564 43812 612592
rect 43548 612510 43576 612564
rect 43806 612552 43812 612564
rect 43864 612552 43870 612604
rect 44082 612388 44088 612400
rect 43663 612360 44088 612388
rect 43663 612306 43691 612360
rect 44082 612348 44088 612360
rect 44140 612348 44146 612400
rect 43898 612212 43904 612264
rect 43956 612252 43962 612264
rect 44450 612252 44456 612264
rect 43956 612224 44456 612252
rect 43956 612212 43962 612224
rect 44450 612212 44456 612224
rect 44508 612212 44514 612264
rect 43766 612196 43818 612202
rect 43766 612138 43818 612144
rect 44082 612048 44088 612060
rect 43887 612020 44088 612048
rect 43887 611966 43915 612020
rect 44082 612008 44088 612020
rect 44140 612008 44146 612060
rect 43996 611788 44048 611794
rect 43996 611730 44048 611736
rect 44088 611584 44140 611590
rect 44088 611526 44140 611532
rect 44450 611396 44456 611448
rect 44508 611396 44514 611448
rect 44205 611328 44211 611380
rect 44263 611328 44269 611380
rect 44468 611300 44496 611396
rect 653398 611328 653404 611380
rect 653456 611368 653462 611380
rect 673454 611368 673460 611380
rect 653456 611340 673460 611368
rect 653456 611328 653462 611340
rect 673454 611328 673460 611340
rect 673512 611328 673518 611380
rect 44468 611272 45140 611300
rect 44312 611124 44318 611176
rect 44370 611124 44376 611176
rect 44910 611164 44916 611176
rect 44447 611136 44916 611164
rect 44447 610946 44475 611136
rect 44910 611124 44916 611136
rect 44968 611124 44974 611176
rect 45112 611028 45140 611272
rect 44560 611000 45140 611028
rect 44560 610742 44588 611000
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 36538 601712 36544 601724
rect 35860 601684 36544 601712
rect 35860 601672 35866 601684
rect 36538 601672 36544 601684
rect 36596 601672 36602 601724
rect 657538 600448 657544 600500
rect 657596 600488 657602 600500
rect 673454 600488 673460 600500
rect 657596 600460 673460 600488
rect 657596 600448 657602 600460
rect 673454 600448 673460 600460
rect 673512 600448 673518 600500
rect 654778 598952 654784 599004
rect 654836 598992 654842 599004
rect 673454 598992 673460 599004
rect 654836 598964 673460 598992
rect 654836 598952 654842 598964
rect 673454 598952 673460 598964
rect 673512 598952 673518 599004
rect 651466 597524 651472 597576
rect 651524 597564 651530 597576
rect 668578 597564 668584 597576
rect 651524 597536 668584 597564
rect 651524 597524 651530 597536
rect 668578 597524 668584 597536
rect 668636 597524 668642 597576
rect 42978 597388 42984 597440
rect 43036 597388 43042 597440
rect 42996 597032 43024 597388
rect 42978 596980 42984 597032
rect 43036 596980 43042 597032
rect 651466 596164 651472 596216
rect 651524 596204 651530 596216
rect 667198 596204 667204 596216
rect 651524 596176 667204 596204
rect 651524 596164 651530 596176
rect 667198 596164 667204 596176
rect 667256 596164 667262 596216
rect 39942 595756 39948 595808
rect 40000 595796 40006 595808
rect 41690 595796 41696 595808
rect 40000 595768 41696 595796
rect 40000 595756 40006 595768
rect 41690 595756 41696 595768
rect 41748 595756 41754 595808
rect 651650 595416 651656 595468
rect 651708 595456 651714 595468
rect 653398 595456 653404 595468
rect 651708 595428 653404 595456
rect 651708 595416 651714 595428
rect 653398 595416 653404 595428
rect 653456 595416 653462 595468
rect 651466 594872 651472 594924
rect 651524 594912 651530 594924
rect 656158 594912 656164 594924
rect 651524 594884 656164 594912
rect 651524 594872 651530 594884
rect 656158 594872 656164 594884
rect 656216 594872 656222 594924
rect 651466 594668 651472 594720
rect 651524 594708 651530 594720
rect 657538 594708 657544 594720
rect 651524 594680 657544 594708
rect 651524 594668 651530 594680
rect 657538 594668 657544 594680
rect 657596 594668 657602 594720
rect 38562 594260 38568 594312
rect 38620 594300 38626 594312
rect 41598 594300 41604 594312
rect 38620 594272 41604 594300
rect 38620 594260 38626 594272
rect 41598 594260 41604 594272
rect 41656 594260 41662 594312
rect 651466 593036 651472 593088
rect 651524 593076 651530 593088
rect 654778 593076 654784 593088
rect 651524 593048 654784 593076
rect 651524 593036 651530 593048
rect 654778 593036 654784 593048
rect 654836 593036 654842 593088
rect 36538 592900 36544 592952
rect 36596 592940 36602 592952
rect 41690 592940 41696 592952
rect 36596 592912 41696 592940
rect 36596 592900 36602 592912
rect 41690 592900 41696 592912
rect 41748 592900 41754 592952
rect 675846 592832 675852 592884
rect 675904 592872 675910 592884
rect 678238 592872 678244 592884
rect 675904 592844 678244 592872
rect 675904 592832 675910 592844
rect 678238 592832 678244 592844
rect 678296 592832 678302 592884
rect 675846 591404 675852 591456
rect 675904 591444 675910 591456
rect 683390 591444 683396 591456
rect 675904 591416 683396 591444
rect 675904 591404 675910 591416
rect 683390 591404 683396 591416
rect 683448 591404 683454 591456
rect 675846 591268 675852 591320
rect 675904 591308 675910 591320
rect 684218 591308 684224 591320
rect 675904 591280 684224 591308
rect 675904 591268 675910 591280
rect 684218 591268 684224 591280
rect 684276 591268 684282 591320
rect 675846 589228 675852 589280
rect 675904 589268 675910 589280
rect 680998 589268 681004 589280
rect 675904 589240 681004 589268
rect 675904 589228 675910 589240
rect 680998 589228 681004 589240
rect 681056 589228 681062 589280
rect 35434 587256 35440 587308
rect 35492 587296 35498 587308
rect 40678 587296 40684 587308
rect 35492 587268 40684 587296
rect 35492 587256 35498 587268
rect 40678 587256 40684 587268
rect 40736 587256 40742 587308
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 41506 587160 41512 587172
rect 33100 587132 41512 587160
rect 33100 587120 33106 587132
rect 41506 587120 41512 587132
rect 41564 587120 41570 587172
rect 33778 585896 33784 585948
rect 33836 585936 33842 585948
rect 40126 585936 40132 585948
rect 33836 585908 40132 585936
rect 33836 585896 33842 585908
rect 40126 585896 40132 585908
rect 40184 585896 40190 585948
rect 31018 585760 31024 585812
rect 31076 585800 31082 585812
rect 40586 585800 40592 585812
rect 31076 585772 40592 585800
rect 31076 585760 31082 585772
rect 40586 585760 40592 585772
rect 40644 585760 40650 585812
rect 652018 581000 652024 581052
rect 652076 581040 652082 581052
rect 674006 581040 674012 581052
rect 652076 581012 674012 581040
rect 652076 581000 652082 581012
rect 674006 581000 674012 581012
rect 674064 581000 674070 581052
rect 669958 580252 669964 580304
rect 670016 580292 670022 580304
rect 674006 580292 674012 580304
rect 670016 580264 674012 580292
rect 670016 580252 670022 580264
rect 674006 580252 674012 580264
rect 674064 580252 674070 580304
rect 671154 579980 671160 580032
rect 671212 580020 671218 580032
rect 674006 580020 674012 580032
rect 671212 579992 674012 580020
rect 671212 579980 671218 579992
rect 674006 579980 674012 579992
rect 674064 579980 674070 580032
rect 658918 579640 658924 579692
rect 658976 579680 658982 579692
rect 673638 579680 673644 579692
rect 658976 579652 673644 579680
rect 658976 579640 658982 579652
rect 673638 579640 673644 579652
rect 673696 579640 673702 579692
rect 671614 578756 671620 578808
rect 671672 578796 671678 578808
rect 674006 578796 674012 578808
rect 671672 578768 674012 578796
rect 671672 578756 671678 578768
rect 674006 578756 674012 578768
rect 674064 578756 674070 578808
rect 670142 578348 670148 578400
rect 670200 578388 670206 578400
rect 674006 578388 674012 578400
rect 670200 578360 674012 578388
rect 670200 578348 670206 578360
rect 674006 578348 674012 578360
rect 674064 578348 674070 578400
rect 669958 578212 669964 578264
rect 670016 578252 670022 578264
rect 673454 578252 673460 578264
rect 670016 578224 673460 578252
rect 670016 578212 670022 578224
rect 673454 578212 673460 578224
rect 673512 578212 673518 578264
rect 42242 577804 42248 577856
rect 42300 577844 42306 577856
rect 42702 577844 42708 577856
rect 42300 577816 42708 577844
rect 42300 577804 42306 577816
rect 42702 577804 42708 577816
rect 42760 577804 42766 577856
rect 669774 577396 669780 577448
rect 669832 577436 669838 577448
rect 674006 577436 674012 577448
rect 669832 577408 674012 577436
rect 669832 577396 669838 577408
rect 674006 577396 674012 577408
rect 674064 577396 674070 577448
rect 669590 577124 669596 577176
rect 669648 577164 669654 577176
rect 673638 577164 673644 577176
rect 669648 577136 673644 577164
rect 669648 577124 669654 577136
rect 673638 577124 673644 577136
rect 673696 577124 673702 577176
rect 670234 576988 670240 577040
rect 670292 577028 670298 577040
rect 673408 577028 673414 577040
rect 670292 577000 673414 577028
rect 670292 576988 670298 577000
rect 673408 576988 673414 577000
rect 673466 576988 673472 577040
rect 674006 576960 674012 576972
rect 673564 576932 674012 576960
rect 671154 576852 671160 576904
rect 671212 576892 671218 576904
rect 673564 576892 673592 576932
rect 674006 576920 674012 576932
rect 674064 576920 674070 576972
rect 671212 576864 673592 576892
rect 671212 576852 671218 576864
rect 671982 575900 671988 575952
rect 672040 575940 672046 575952
rect 674006 575940 674012 575952
rect 672040 575912 674012 575940
rect 672040 575900 672046 575912
rect 674006 575900 674012 575912
rect 674064 575900 674070 575952
rect 44634 575424 44640 575476
rect 44692 575464 44698 575476
rect 62114 575464 62120 575476
rect 44692 575436 62120 575464
rect 44692 575424 44698 575436
rect 62114 575424 62120 575436
rect 62172 575424 62178 575476
rect 668210 574404 668216 574456
rect 668268 574444 668274 574456
rect 674006 574444 674012 574456
rect 668268 574416 674012 574444
rect 668268 574404 668274 574416
rect 674006 574404 674012 574416
rect 674064 574404 674070 574456
rect 668854 574132 668860 574184
rect 668912 574172 668918 574184
rect 673638 574172 673644 574184
rect 668912 574144 673644 574172
rect 668912 574132 668918 574144
rect 673638 574132 673644 574144
rect 673696 574132 673702 574184
rect 45554 573996 45560 574048
rect 45612 574036 45618 574048
rect 62114 574036 62120 574048
rect 45612 574008 62120 574036
rect 45612 573996 45618 574008
rect 62114 573996 62120 574008
rect 62172 573996 62178 574048
rect 42150 573452 42156 573504
rect 42208 573492 42214 573504
rect 42610 573492 42616 573504
rect 42208 573464 42616 573492
rect 42208 573452 42214 573464
rect 42610 573452 42616 573464
rect 42668 573452 42674 573504
rect 671798 572840 671804 572892
rect 671856 572880 671862 572892
rect 674006 572880 674012 572892
rect 671856 572852 674012 572880
rect 671856 572840 671862 572852
rect 674006 572840 674012 572852
rect 674064 572840 674070 572892
rect 667382 571684 667388 571736
rect 667440 571724 667446 571736
rect 673638 571724 673644 571736
rect 667440 571696 673644 571724
rect 667440 571684 667446 571696
rect 673638 571684 673644 571696
rect 673696 571684 673702 571736
rect 669038 571412 669044 571464
rect 669096 571452 669102 571464
rect 674006 571452 674012 571464
rect 669096 571424 674012 571452
rect 669096 571412 669102 571424
rect 674006 571412 674012 571424
rect 674064 571412 674070 571464
rect 680998 571276 681004 571328
rect 681056 571316 681062 571328
rect 683114 571316 683120 571328
rect 681056 571288 683120 571316
rect 681056 571276 681062 571288
rect 683114 571276 683120 571288
rect 683172 571276 683178 571328
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 42610 570976 42616 570988
rect 42116 570948 42616 570976
rect 42116 570936 42122 570948
rect 42610 570936 42616 570948
rect 42668 570936 42674 570988
rect 653398 565836 653404 565888
rect 653456 565876 653462 565888
rect 674006 565876 674012 565888
rect 653456 565848 674012 565876
rect 653456 565836 653462 565848
rect 674006 565836 674012 565848
rect 674064 565836 674070 565888
rect 672718 557812 672724 557864
rect 672776 557852 672782 557864
rect 673270 557852 673276 557864
rect 672776 557824 673276 557852
rect 672776 557812 672782 557824
rect 673270 557812 673276 557824
rect 673328 557812 673334 557864
rect 673822 556588 673828 556640
rect 673880 556628 673886 556640
rect 674006 556628 674012 556640
rect 673880 556600 674012 556628
rect 673880 556588 673886 556600
rect 674006 556588 674012 556600
rect 674064 556588 674070 556640
rect 672718 555432 672724 555484
rect 672776 555472 672782 555484
rect 673270 555472 673276 555484
rect 672776 555444 673276 555472
rect 672776 555432 672782 555444
rect 673270 555432 673276 555444
rect 673328 555432 673334 555484
rect 674650 554888 674656 554940
rect 674708 554928 674714 554940
rect 675110 554928 675116 554940
rect 674708 554900 675116 554928
rect 674708 554888 674714 554900
rect 675110 554888 675116 554900
rect 675168 554888 675174 554940
rect 674006 554860 674012 554872
rect 669286 554832 674012 554860
rect 657814 554752 657820 554804
rect 657872 554792 657878 554804
rect 669286 554792 669314 554832
rect 674006 554820 674012 554832
rect 674064 554820 674070 554872
rect 657872 554764 669314 554792
rect 657872 554752 657878 554764
rect 655146 553392 655152 553444
rect 655204 553432 655210 553444
rect 674006 553432 674012 553444
rect 655204 553404 674012 553432
rect 655204 553392 655210 553404
rect 674006 553392 674012 553404
rect 674064 553392 674070 553444
rect 651466 552644 651472 552696
rect 651524 552684 651530 552696
rect 665818 552684 665824 552696
rect 651524 552656 665824 552684
rect 651524 552644 651530 552656
rect 665818 552644 665824 552656
rect 665876 552644 665882 552696
rect 651466 552032 651472 552084
rect 651524 552072 651530 552084
rect 660298 552072 660304 552084
rect 651524 552044 660304 552072
rect 651524 552032 651530 552044
rect 660298 552032 660304 552044
rect 660356 552032 660362 552084
rect 40034 550944 40040 550996
rect 40092 550984 40098 550996
rect 41690 550984 41696 550996
rect 40092 550956 41696 550984
rect 40092 550944 40098 550956
rect 41690 550944 41696 550956
rect 41748 550944 41754 550996
rect 668854 550604 668860 550656
rect 668912 550644 668918 550656
rect 673454 550644 673460 550656
rect 668912 550616 673460 550644
rect 668912 550604 668918 550616
rect 673454 550604 673460 550616
rect 673512 550604 673518 550656
rect 651374 550332 651380 550384
rect 651432 550372 651438 550384
rect 653398 550372 653404 550384
rect 651432 550344 653404 550372
rect 651432 550332 651438 550344
rect 653398 550332 653404 550344
rect 653456 550332 653462 550384
rect 651466 549040 651472 549092
rect 651524 549080 651530 549092
rect 657814 549080 657820 549092
rect 651524 549052 657820 549080
rect 651524 549040 651530 549052
rect 657814 549040 657820 549052
rect 657872 549040 657878 549092
rect 673178 548904 673184 548956
rect 673236 548904 673242 548956
rect 651466 548768 651472 548820
rect 651524 548808 651530 548820
rect 655146 548808 655152 548820
rect 651524 548780 655152 548808
rect 651524 548768 651530 548780
rect 655146 548768 655152 548780
rect 655204 548768 655210 548820
rect 672994 548496 673000 548548
rect 673052 548536 673058 548548
rect 673196 548536 673224 548904
rect 673052 548508 673224 548536
rect 673052 548496 673058 548508
rect 675478 547584 675484 547596
rect 674806 547556 675484 547584
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 41690 547448 41696 547460
rect 31812 547420 41696 547448
rect 31812 547408 31818 547420
rect 41690 547408 41696 547420
rect 41748 547408 41754 547460
rect 674282 547408 674288 547460
rect 674340 547448 674346 547460
rect 674806 547448 674834 547556
rect 675478 547544 675484 547556
rect 675536 547544 675542 547596
rect 675846 547544 675852 547596
rect 675904 547584 675910 547596
rect 684218 547584 684224 547596
rect 675904 547556 684224 547584
rect 675904 547544 675910 547556
rect 684218 547544 684224 547556
rect 684276 547544 684282 547596
rect 674340 547420 674834 547448
rect 674340 547408 674346 547420
rect 676030 547408 676036 547460
rect 676088 547448 676094 547460
rect 683390 547448 683396 547460
rect 676088 547420 683396 547448
rect 676088 547408 676094 547420
rect 683390 547408 683396 547420
rect 683448 547408 683454 547460
rect 675478 547312 675484 547324
rect 674806 547284 675484 547312
rect 674282 547136 674288 547188
rect 674340 547176 674346 547188
rect 674806 547176 674834 547284
rect 675478 547272 675484 547284
rect 675536 547272 675542 547324
rect 675846 547272 675852 547324
rect 675904 547312 675910 547324
rect 683206 547312 683212 547324
rect 675904 547284 683212 547312
rect 675904 547272 675910 547284
rect 683206 547272 683212 547284
rect 683264 547272 683270 547324
rect 674340 547148 674834 547176
rect 674340 547136 674346 547148
rect 674282 547000 674288 547052
rect 674340 547040 674346 547052
rect 675478 547040 675484 547052
rect 674340 547012 675484 547040
rect 674340 547000 674346 547012
rect 675478 547000 675484 547012
rect 675536 547000 675542 547052
rect 34422 544348 34428 544400
rect 34480 544388 34486 544400
rect 41322 544388 41328 544400
rect 34480 544360 41328 544388
rect 34480 544348 34486 544360
rect 41322 544348 41328 544360
rect 41380 544348 41386 544400
rect 42978 538160 42984 538212
rect 43036 538160 43042 538212
rect 42794 537888 42800 537940
rect 42852 537928 42858 537940
rect 42996 537928 43024 538160
rect 42852 537900 43024 537928
rect 42852 537888 42858 537900
rect 668578 535644 668584 535696
rect 668636 535684 668642 535696
rect 674006 535684 674012 535696
rect 668636 535656 674012 535684
rect 668636 535644 668642 535656
rect 674006 535644 674012 535656
rect 674064 535644 674070 535696
rect 667198 535440 667204 535492
rect 667256 535480 667262 535492
rect 673822 535480 673828 535492
rect 667256 535452 673828 535480
rect 667256 535440 667262 535452
rect 673822 535440 673828 535452
rect 673880 535440 673886 535492
rect 669958 534488 669964 534540
rect 670016 534528 670022 534540
rect 674006 534528 674012 534540
rect 670016 534500 674012 534528
rect 670016 534488 670022 534500
rect 674006 534488 674012 534500
rect 674064 534488 674070 534540
rect 670142 534352 670148 534404
rect 670200 534392 670206 534404
rect 674006 534392 674012 534404
rect 670200 534364 674012 534392
rect 670200 534352 670206 534364
rect 674006 534352 674012 534364
rect 674064 534352 674070 534404
rect 656158 534216 656164 534268
rect 656216 534256 656222 534268
rect 673454 534256 673460 534268
rect 656216 534228 673460 534256
rect 656216 534216 656222 534228
rect 673454 534216 673460 534228
rect 673512 534216 673518 534268
rect 670786 534080 670792 534132
rect 670844 534120 670850 534132
rect 673822 534120 673828 534132
rect 670844 534092 673828 534120
rect 670844 534080 670850 534092
rect 673822 534080 673828 534092
rect 673880 534080 673886 534132
rect 671614 533536 671620 533588
rect 671672 533576 671678 533588
rect 674006 533576 674012 533588
rect 671672 533548 674012 533576
rect 671672 533536 671678 533548
rect 674006 533536 674012 533548
rect 674064 533536 674070 533588
rect 670234 533332 670240 533384
rect 670292 533372 670298 533384
rect 674006 533372 674012 533384
rect 670292 533344 674012 533372
rect 670292 533332 670298 533344
rect 674006 533332 674012 533344
rect 674064 533332 674070 533384
rect 675846 533332 675852 533384
rect 675904 533372 675910 533384
rect 683574 533372 683580 533384
rect 675904 533344 683580 533372
rect 675904 533332 675910 533344
rect 683574 533332 683580 533344
rect 683632 533332 683638 533384
rect 42426 532720 42432 532772
rect 42484 532760 42490 532772
rect 43162 532760 43168 532772
rect 42484 532732 43168 532760
rect 42484 532720 42490 532732
rect 43162 532720 43168 532732
rect 43220 532720 43226 532772
rect 671798 532720 671804 532772
rect 671856 532760 671862 532772
rect 674006 532760 674012 532772
rect 671856 532732 674012 532760
rect 671856 532720 671862 532732
rect 674006 532720 674012 532732
rect 674064 532720 674070 532772
rect 671154 532516 671160 532568
rect 671212 532556 671218 532568
rect 674006 532556 674012 532568
rect 671212 532528 674012 532556
rect 671212 532516 671218 532528
rect 674006 532516 674012 532528
rect 674064 532516 674070 532568
rect 672442 531904 672448 531956
rect 672500 531944 672506 531956
rect 674006 531944 674012 531956
rect 672500 531916 674012 531944
rect 672500 531904 672506 531916
rect 674006 531904 674012 531916
rect 674064 531904 674070 531956
rect 672626 531700 672632 531752
rect 672684 531740 672690 531752
rect 674006 531740 674012 531752
rect 672684 531712 674012 531740
rect 672684 531700 672690 531712
rect 674006 531700 674012 531712
rect 674064 531700 674070 531752
rect 59998 531224 60004 531276
rect 60056 531264 60062 531276
rect 62114 531264 62120 531276
rect 60056 531236 62120 531264
rect 60056 531224 60062 531236
rect 62114 531224 62120 531236
rect 62172 531224 62178 531276
rect 44726 531088 44732 531140
rect 44784 531128 44790 531140
rect 62114 531128 62120 531140
rect 44784 531100 62120 531128
rect 44784 531088 44790 531100
rect 62114 531088 62120 531100
rect 62172 531088 62178 531140
rect 672718 530204 672724 530256
rect 672776 530244 672782 530256
rect 673454 530244 673460 530256
rect 672776 530216 673460 530244
rect 672776 530204 672782 530216
rect 673454 530204 673460 530216
rect 673512 530204 673518 530256
rect 42150 530068 42156 530120
rect 42208 530108 42214 530120
rect 42978 530108 42984 530120
rect 42208 530080 42984 530108
rect 42208 530068 42214 530080
rect 42978 530068 42984 530080
rect 43036 530068 43042 530120
rect 670418 530068 670424 530120
rect 670476 530108 670482 530120
rect 673822 530108 673828 530120
rect 670476 530080 673828 530108
rect 670476 530068 670482 530080
rect 673822 530068 673828 530080
rect 673880 530068 673886 530120
rect 667566 529932 667572 529984
rect 667624 529972 667630 529984
rect 674006 529972 674012 529984
rect 667624 529944 674012 529972
rect 667624 529932 667630 529944
rect 674006 529932 674012 529944
rect 674064 529932 674070 529984
rect 670970 529660 670976 529712
rect 671028 529700 671034 529712
rect 674006 529700 674012 529712
rect 671028 529672 674012 529700
rect 671028 529660 671034 529672
rect 674006 529660 674012 529672
rect 674064 529660 674070 529712
rect 45094 528572 45100 528624
rect 45152 528612 45158 528624
rect 62114 528612 62120 528624
rect 45152 528584 62120 528612
rect 45152 528572 45158 528584
rect 62114 528572 62120 528584
rect 62172 528572 62178 528624
rect 669222 528572 669228 528624
rect 669280 528612 669286 528624
rect 674006 528612 674012 528624
rect 669280 528584 674012 528612
rect 669280 528572 669286 528584
rect 674006 528572 674012 528584
rect 674064 528572 674070 528624
rect 672258 528436 672264 528488
rect 672316 528476 672322 528488
rect 674006 528476 674012 528488
rect 672316 528448 674012 528476
rect 672316 528436 672322 528448
rect 674006 528436 674012 528448
rect 674064 528436 674070 528488
rect 42058 527756 42064 527808
rect 42116 527796 42122 527808
rect 42610 527796 42616 527808
rect 42116 527768 42616 527796
rect 42116 527756 42122 527768
rect 42610 527756 42616 527768
rect 42668 527756 42674 527808
rect 672718 526464 672724 526516
rect 672776 526504 672782 526516
rect 673270 526504 673276 526516
rect 672776 526476 673276 526504
rect 672776 526464 672782 526476
rect 673270 526464 673276 526476
rect 673328 526464 673334 526516
rect 671338 524628 671344 524680
rect 671396 524668 671402 524680
rect 674006 524668 674012 524680
rect 671396 524640 674012 524668
rect 671396 524628 671402 524640
rect 674006 524628 674012 524640
rect 674064 524628 674070 524680
rect 675846 524560 675852 524612
rect 675904 524600 675910 524612
rect 683114 524600 683120 524612
rect 675904 524572 683120 524600
rect 675904 524560 675910 524572
rect 683114 524560 683120 524572
rect 683172 524560 683178 524612
rect 675846 518848 675852 518900
rect 675904 518888 675910 518900
rect 677686 518888 677692 518900
rect 675904 518860 677692 518888
rect 675904 518848 675910 518860
rect 677686 518848 677692 518860
rect 677744 518848 677750 518900
rect 677870 518780 677876 518832
rect 677928 518780 677934 518832
rect 676030 518644 676036 518696
rect 676088 518684 676094 518696
rect 677888 518684 677916 518780
rect 676088 518656 677916 518684
rect 676088 518644 676094 518656
rect 675294 503888 675300 503940
rect 675352 503888 675358 503940
rect 675478 503888 675484 503940
rect 675536 503888 675542 503940
rect 675312 503668 675340 503888
rect 675496 503668 675524 503888
rect 676122 503752 676128 503804
rect 676180 503792 676186 503804
rect 678238 503792 678244 503804
rect 676180 503764 678244 503792
rect 676180 503752 676186 503764
rect 678238 503752 678244 503764
rect 678296 503752 678302 503804
rect 675294 503616 675300 503668
rect 675352 503616 675358 503668
rect 675478 503616 675484 503668
rect 675536 503616 675542 503668
rect 677410 503616 677416 503668
rect 677468 503656 677474 503668
rect 683390 503656 683396 503668
rect 677468 503628 683396 503656
rect 677468 503616 677474 503628
rect 683390 503616 683396 503628
rect 683448 503616 683454 503668
rect 675846 500760 675852 500812
rect 675904 500800 675910 500812
rect 680998 500800 681004 500812
rect 675904 500772 681004 500800
rect 675904 500760 675910 500772
rect 680998 500760 681004 500772
rect 681056 500760 681062 500812
rect 652018 493280 652024 493332
rect 652076 493320 652082 493332
rect 672902 493320 672908 493332
rect 652076 493292 672908 493320
rect 652076 493280 652082 493292
rect 672902 493280 672908 493292
rect 672960 493280 672966 493332
rect 665818 491444 665824 491496
rect 665876 491484 665882 491496
rect 674006 491484 674012 491496
rect 665876 491456 674012 491484
rect 665876 491444 665882 491456
rect 674006 491444 674012 491456
rect 674064 491444 674070 491496
rect 660298 491308 660304 491360
rect 660356 491348 660362 491360
rect 673822 491348 673828 491360
rect 660356 491320 673828 491348
rect 660356 491308 660362 491320
rect 673822 491308 673828 491320
rect 673880 491308 673886 491360
rect 670786 490900 670792 490952
rect 670844 490940 670850 490952
rect 674006 490940 674012 490952
rect 670844 490912 674012 490940
rect 670844 490900 670850 490912
rect 674006 490900 674012 490912
rect 674064 490900 674070 490952
rect 671614 490084 671620 490136
rect 671672 490124 671678 490136
rect 674006 490124 674012 490136
rect 671672 490096 674012 490124
rect 671672 490084 671678 490096
rect 674006 490084 674012 490096
rect 674064 490084 674070 490136
rect 676030 490016 676036 490068
rect 676088 490056 676094 490068
rect 676582 490056 676588 490068
rect 676088 490028 676588 490056
rect 676088 490016 676094 490028
rect 676582 490016 676588 490028
rect 676640 490016 676646 490068
rect 672626 489608 672632 489660
rect 672684 489648 672690 489660
rect 674006 489648 674012 489660
rect 672684 489620 674012 489648
rect 672684 489608 672690 489620
rect 674006 489608 674012 489620
rect 674064 489608 674070 489660
rect 671798 489268 671804 489320
rect 671856 489308 671862 489320
rect 674006 489308 674012 489320
rect 671856 489280 674012 489308
rect 671856 489268 671862 489280
rect 674006 489268 674012 489280
rect 674064 489268 674070 489320
rect 672442 488452 672448 488504
rect 672500 488492 672506 488504
rect 674006 488492 674012 488504
rect 672500 488464 674012 488492
rect 672500 488452 672506 488464
rect 674006 488452 674012 488464
rect 674064 488452 674070 488504
rect 676214 487160 676220 487212
rect 676272 487200 676278 487212
rect 677502 487200 677508 487212
rect 676272 487172 677508 487200
rect 676272 487160 676278 487172
rect 677502 487160 677508 487172
rect 677560 487160 677566 487212
rect 668394 485800 668400 485852
rect 668452 485840 668458 485852
rect 674006 485840 674012 485852
rect 668452 485812 674012 485840
rect 668452 485800 668458 485812
rect 674006 485800 674012 485812
rect 674064 485800 674070 485852
rect 669038 484508 669044 484560
rect 669096 484548 669102 484560
rect 674006 484548 674012 484560
rect 669096 484520 674012 484548
rect 669096 484508 669102 484520
rect 674006 484508 674012 484520
rect 674064 484508 674070 484560
rect 668854 484372 668860 484424
rect 668912 484412 668918 484424
rect 673822 484412 673828 484424
rect 668912 484384 673828 484412
rect 668912 484372 668918 484384
rect 673822 484372 673828 484384
rect 673880 484372 673886 484424
rect 671982 482332 671988 482384
rect 672040 482372 672046 482384
rect 674006 482372 674012 482384
rect 672040 482344 674012 482372
rect 672040 482332 672046 482344
rect 674006 482332 674012 482344
rect 674064 482332 674070 482384
rect 676122 480360 676128 480412
rect 676180 480400 676186 480412
rect 683114 480400 683120 480412
rect 676180 480372 683120 480400
rect 676180 480360 676186 480372
rect 683114 480360 683120 480372
rect 683172 480360 683178 480412
rect 670602 456356 670608 456408
rect 670660 456396 670666 456408
rect 670660 456368 673988 456396
rect 670660 456356 670666 456368
rect 673960 456246 673988 456368
rect 676214 456192 676220 456204
rect 676048 456164 676220 456192
rect 676048 455988 676076 456164
rect 676214 456152 676220 456164
rect 676272 456152 676278 456204
rect 676168 455988 676174 456000
rect 676048 455960 676174 455988
rect 676168 455948 676174 455960
rect 676226 455948 676232 456000
rect 673828 455864 673880 455870
rect 673270 455812 673276 455864
rect 673328 455852 673334 455864
rect 673328 455824 673762 455852
rect 673328 455812 673334 455824
rect 673828 455806 673880 455812
rect 667842 455608 667848 455660
rect 667900 455648 667906 455660
rect 667900 455620 673624 455648
rect 667900 455608 667906 455620
rect 673270 455336 673276 455388
rect 673328 455376 673334 455388
rect 673328 455348 673532 455376
rect 673328 455336 673334 455348
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 673276 455048 673328 455054
rect 673276 454990 673328 454996
rect 672074 454792 672080 454844
rect 672132 454832 672138 454844
rect 672132 454804 673190 454832
rect 672132 454792 672138 454804
rect 673046 454640 673098 454646
rect 673046 454582 673098 454588
rect 672954 454368 673006 454374
rect 674282 454316 674288 454368
rect 674340 454356 674346 454368
rect 675478 454356 675484 454368
rect 674340 454328 675484 454356
rect 674340 454316 674346 454328
rect 675478 454316 675484 454328
rect 675536 454316 675542 454368
rect 672954 454310 673006 454316
rect 672816 454096 672868 454102
rect 672816 454038 672868 454044
rect 672442 453908 672448 453960
rect 672500 453948 672506 453960
rect 672500 453920 672750 453948
rect 672500 453908 672506 453920
rect 35802 429156 35808 429208
rect 35860 429196 35866 429208
rect 41690 429196 41696 429208
rect 35860 429168 41696 429196
rect 35860 429156 35866 429168
rect 41690 429156 41696 429168
rect 41748 429156 41754 429208
rect 41322 425076 41328 425128
rect 41380 425116 41386 425128
rect 41690 425116 41696 425128
rect 41380 425088 41696 425116
rect 41380 425076 41386 425088
rect 41690 425076 41696 425088
rect 41748 425076 41754 425128
rect 40954 424260 40960 424312
rect 41012 424300 41018 424312
rect 41506 424300 41512 424312
rect 41012 424272 41512 424300
rect 41012 424260 41018 424272
rect 41506 424260 41512 424272
rect 41564 424260 41570 424312
rect 32030 416168 32036 416220
rect 32088 416208 32094 416220
rect 41690 416208 41696 416220
rect 32088 416180 41696 416208
rect 32088 416168 32094 416180
rect 41690 416168 41696 416180
rect 41748 416168 41754 416220
rect 53834 404268 53840 404320
rect 53892 404308 53898 404320
rect 62114 404308 62120 404320
rect 53892 404280 62120 404308
rect 53892 404268 53898 404280
rect 62114 404268 62120 404280
rect 62172 404268 62178 404320
rect 44818 402908 44824 402960
rect 44876 402948 44882 402960
rect 62114 402948 62120 402960
rect 44876 402920 62120 402948
rect 44876 402908 44882 402920
rect 62114 402908 62120 402920
rect 62172 402908 62178 402960
rect 51074 400188 51080 400240
rect 51132 400228 51138 400240
rect 62114 400228 62120 400240
rect 51132 400200 62120 400228
rect 51132 400188 51138 400200
rect 62114 400188 62120 400200
rect 62172 400188 62178 400240
rect 59998 400052 60004 400104
rect 60056 400092 60062 400104
rect 62114 400092 62120 400104
rect 60056 400064 62120 400092
rect 60056 400052 60062 400064
rect 62114 400052 62120 400064
rect 62172 400052 62178 400104
rect 674834 385568 674840 385620
rect 674892 385608 674898 385620
rect 675294 385608 675300 385620
rect 674892 385580 675300 385608
rect 674892 385568 674898 385580
rect 675294 385568 675300 385580
rect 675352 385568 675358 385620
rect 41322 382236 41328 382288
rect 41380 382276 41386 382288
rect 41690 382276 41696 382288
rect 41380 382248 41696 382276
rect 41380 382236 41386 382248
rect 41690 382236 41696 382248
rect 41748 382236 41754 382288
rect 674466 382168 674472 382220
rect 674524 382208 674530 382220
rect 675386 382208 675392 382220
rect 674524 382180 675392 382208
rect 674524 382168 674530 382180
rect 675386 382168 675392 382180
rect 675444 382168 675450 382220
rect 35802 379652 35808 379704
rect 35860 379692 35866 379704
rect 40586 379692 40592 379704
rect 35860 379664 40592 379692
rect 35860 379652 35866 379664
rect 40586 379652 40592 379664
rect 40644 379652 40650 379704
rect 674374 378088 674380 378140
rect 674432 378128 674438 378140
rect 675110 378128 675116 378140
rect 674432 378100 675116 378128
rect 674432 378088 674438 378100
rect 675110 378088 675116 378100
rect 675168 378088 675174 378140
rect 40218 378020 40224 378072
rect 40276 378060 40282 378072
rect 41690 378060 41696 378072
rect 40276 378032 41696 378060
rect 40276 378020 40282 378032
rect 41690 378020 41696 378032
rect 41748 378020 41754 378072
rect 42058 377952 42064 378004
rect 42116 377992 42122 378004
rect 42702 377992 42708 378004
rect 42116 377964 42708 377992
rect 42116 377952 42122 377964
rect 42702 377952 42708 377964
rect 42760 377952 42766 378004
rect 651466 373940 651472 373992
rect 651524 373980 651530 373992
rect 657538 373980 657544 373992
rect 651524 373952 657544 373980
rect 651524 373940 651530 373952
rect 657538 373940 657544 373952
rect 657596 373940 657602 373992
rect 35158 371832 35164 371884
rect 35216 371872 35222 371884
rect 41690 371872 41696 371884
rect 35216 371844 41696 371872
rect 35216 371832 35222 371844
rect 41690 371832 41696 371844
rect 41748 371832 41754 371884
rect 651466 370948 651472 371000
rect 651524 370988 651530 371000
rect 654778 370988 654784 371000
rect 651524 370960 654784 370988
rect 651524 370948 651530 370960
rect 654778 370948 654784 370960
rect 654836 370948 654842 371000
rect 42242 365236 42248 365288
rect 42300 365236 42306 365288
rect 42260 364948 42288 365236
rect 42242 364896 42248 364948
rect 42300 364896 42306 364948
rect 42242 364284 42248 364336
rect 42300 364284 42306 364336
rect 42260 364188 42288 364284
rect 42702 364188 42708 364200
rect 42260 364160 42708 364188
rect 42702 364148 42708 364160
rect 42760 364148 42766 364200
rect 46566 361496 46572 361548
rect 46624 361536 46630 361548
rect 62114 361536 62120 361548
rect 46624 361508 62120 361536
rect 46624 361496 46630 361508
rect 62114 361496 62120 361508
rect 62172 361496 62178 361548
rect 45370 360136 45376 360188
rect 45428 360176 45434 360188
rect 62114 360176 62120 360188
rect 45428 360148 62120 360176
rect 45428 360136 45434 360148
rect 62114 360136 62120 360148
rect 62172 360136 62178 360188
rect 44634 359592 44640 359644
rect 44692 359632 44698 359644
rect 45370 359632 45376 359644
rect 44692 359604 45376 359632
rect 44692 359592 44698 359604
rect 45370 359592 45376 359604
rect 45428 359592 45434 359644
rect 44818 359456 44824 359508
rect 44876 359496 44882 359508
rect 45462 359496 45468 359508
rect 44876 359468 45468 359496
rect 44876 359456 44882 359468
rect 45462 359456 45468 359468
rect 45520 359456 45526 359508
rect 51718 357416 51724 357468
rect 51776 357456 51782 357468
rect 62114 357456 62120 357468
rect 51776 357428 62120 357456
rect 51776 357416 51782 357428
rect 62114 357416 62120 357428
rect 62172 357416 62178 357468
rect 44640 354748 44692 354754
rect 44818 354696 44824 354748
rect 44876 354696 44882 354748
rect 44640 354690 44692 354696
rect 44836 354600 44864 354696
rect 44836 354572 45002 354600
rect 44732 354476 44784 354482
rect 44849 354424 44855 354476
rect 44907 354424 44913 354476
rect 44732 354418 44784 354424
rect 44867 354314 44895 354424
rect 44974 354110 45002 354572
rect 45830 353920 45836 353932
rect 45105 353892 45836 353920
rect 45830 353880 45836 353892
rect 45888 353880 45894 353932
rect 45830 353716 45836 353728
rect 45218 353688 45836 353716
rect 45830 353676 45836 353688
rect 45888 353676 45894 353728
rect 45303 353524 45355 353530
rect 45303 353466 45355 353472
rect 45422 353252 45474 353258
rect 45422 353194 45474 353200
rect 676030 347420 676036 347472
rect 676088 347460 676094 347472
rect 676490 347460 676496 347472
rect 676088 347432 676496 347460
rect 676088 347420 676094 347432
rect 676490 347420 676496 347432
rect 676548 347420 676554 347472
rect 35802 344564 35808 344616
rect 35860 344604 35866 344616
rect 39850 344604 39856 344616
rect 35860 344576 39856 344604
rect 35860 344564 35866 344576
rect 39850 344564 39856 344576
rect 39908 344564 39914 344616
rect 35618 343612 35624 343664
rect 35676 343652 35682 343664
rect 40034 343652 40040 343664
rect 35676 343624 40040 343652
rect 35676 343612 35682 343624
rect 40034 343612 40040 343624
rect 40092 343612 40098 343664
rect 35802 342184 35808 342236
rect 35860 342224 35866 342236
rect 40218 342224 40224 342236
rect 35860 342196 40224 342224
rect 35860 342184 35866 342196
rect 40218 342184 40224 342196
rect 40276 342184 40282 342236
rect 45462 342184 45468 342236
rect 45520 342224 45526 342236
rect 63126 342224 63132 342236
rect 45520 342196 63132 342224
rect 45520 342184 45526 342196
rect 63126 342184 63132 342196
rect 63184 342184 63190 342236
rect 35802 341504 35808 341556
rect 35860 341544 35866 341556
rect 40218 341544 40224 341556
rect 35860 341516 40224 341544
rect 35860 341504 35866 341516
rect 40218 341504 40224 341516
rect 40276 341504 40282 341556
rect 35802 341028 35808 341080
rect 35860 341068 35866 341080
rect 40126 341068 40132 341080
rect 35860 341040 40132 341068
rect 35860 341028 35866 341040
rect 40126 341028 40132 341040
rect 40184 341028 40190 341080
rect 35526 339600 35532 339652
rect 35584 339640 35590 339652
rect 37090 339640 37096 339652
rect 35584 339612 37096 339640
rect 35584 339600 35590 339612
rect 37090 339600 37096 339612
rect 37148 339600 37154 339652
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 38838 339504 38844 339516
rect 35860 339476 38844 339504
rect 35860 339464 35866 339476
rect 38838 339464 38844 339476
rect 38896 339464 38902 339516
rect 674834 339328 674840 339380
rect 674892 339368 674898 339380
rect 675478 339368 675484 339380
rect 674892 339340 675484 339368
rect 674892 339328 674898 339340
rect 675478 339328 675484 339340
rect 675536 339328 675542 339380
rect 674374 336540 674380 336592
rect 674432 336580 674438 336592
rect 675386 336580 675392 336592
rect 674432 336552 675392 336580
rect 674432 336540 674438 336552
rect 675386 336540 675392 336552
rect 675444 336540 675450 336592
rect 35802 335316 35808 335368
rect 35860 335356 35866 335368
rect 39850 335356 39856 335368
rect 35860 335328 39856 335356
rect 35860 335316 35866 335328
rect 39850 335316 39856 335328
rect 39908 335316 39914 335368
rect 35802 334092 35808 334144
rect 35860 334132 35866 334144
rect 40310 334132 40316 334144
rect 35860 334104 40316 334132
rect 35860 334092 35866 334104
rect 40310 334092 40316 334104
rect 40368 334092 40374 334144
rect 651374 328244 651380 328296
rect 651432 328284 651438 328296
rect 654778 328284 654784 328296
rect 651432 328256 654784 328284
rect 651432 328244 651438 328256
rect 654778 328244 654784 328256
rect 654836 328244 654842 328296
rect 651374 325592 651380 325644
rect 651432 325632 651438 325644
rect 653398 325632 653404 325644
rect 651432 325604 653404 325632
rect 651432 325592 651438 325604
rect 653398 325592 653404 325604
rect 653456 325592 653462 325644
rect 53834 317364 53840 317416
rect 53892 317404 53898 317416
rect 62114 317404 62120 317416
rect 53892 317376 62120 317404
rect 53892 317364 53898 317376
rect 62114 317364 62120 317376
rect 62172 317364 62178 317416
rect 53098 315936 53104 315988
rect 53156 315976 53162 315988
rect 62114 315976 62120 315988
rect 53156 315948 62120 315976
rect 53156 315936 53162 315948
rect 62114 315936 62120 315948
rect 62172 315936 62178 315988
rect 59906 314712 59912 314764
rect 59964 314752 59970 314764
rect 62114 314752 62120 314764
rect 59964 314724 62120 314752
rect 59964 314712 59970 314724
rect 62114 314712 62120 314724
rect 62172 314712 62178 314764
rect 676214 307776 676220 307828
rect 676272 307816 676278 307828
rect 676858 307816 676864 307828
rect 676272 307788 676864 307816
rect 676272 307776 676278 307788
rect 676858 307776 676864 307788
rect 676916 307776 676922 307828
rect 675846 304104 675852 304156
rect 675904 304144 675910 304156
rect 676214 304144 676220 304156
rect 675904 304116 676220 304144
rect 675904 304104 675910 304116
rect 676214 304104 676220 304116
rect 676272 304104 676278 304156
rect 651374 303492 651380 303544
rect 651432 303532 651438 303544
rect 653398 303532 653404 303544
rect 651432 303504 653404 303532
rect 651432 303492 651438 303504
rect 653398 303492 653404 303504
rect 653456 303492 653462 303544
rect 651466 300772 651472 300824
rect 651524 300812 651530 300824
rect 664438 300812 664444 300824
rect 651524 300784 664444 300812
rect 651524 300772 651530 300784
rect 664438 300772 664444 300784
rect 664496 300772 664502 300824
rect 35618 298732 35624 298784
rect 35676 298772 35682 298784
rect 41598 298772 41604 298784
rect 35676 298744 41604 298772
rect 35676 298732 35682 298744
rect 41598 298732 41604 298744
rect 41656 298732 41662 298784
rect 35802 298256 35808 298308
rect 35860 298296 35866 298308
rect 41598 298296 41604 298308
rect 35860 298268 41604 298296
rect 35860 298256 35866 298268
rect 41598 298256 41604 298268
rect 41656 298256 41662 298308
rect 651466 298120 651472 298172
rect 651524 298160 651530 298172
rect 662414 298160 662420 298172
rect 651524 298132 662420 298160
rect 651524 298120 651530 298132
rect 662414 298120 662420 298132
rect 662472 298120 662478 298172
rect 675846 298052 675852 298104
rect 675904 298092 675910 298104
rect 676858 298092 676864 298104
rect 675904 298064 676864 298092
rect 675904 298052 675910 298064
rect 676858 298052 676864 298064
rect 676916 298052 676922 298104
rect 676122 297916 676128 297968
rect 676180 297956 676186 297968
rect 679618 297956 679624 297968
rect 676180 297928 679624 297956
rect 676180 297916 676186 297928
rect 679618 297916 679624 297928
rect 679676 297916 679682 297968
rect 675938 297440 675944 297492
rect 675996 297480 676002 297492
rect 677594 297480 677600 297492
rect 675996 297452 677600 297480
rect 675996 297440 676002 297452
rect 677594 297440 677600 297452
rect 677652 297440 677658 297492
rect 651466 297032 651472 297084
rect 651524 297072 651530 297084
rect 656158 297072 656164 297084
rect 651524 297044 656164 297072
rect 651524 297032 651530 297044
rect 656158 297032 656164 297044
rect 656216 297032 656222 297084
rect 675478 296352 675484 296404
rect 675536 296352 675542 296404
rect 652662 295944 652668 295996
rect 652720 295984 652726 295996
rect 665818 295984 665824 295996
rect 652720 295956 665824 295984
rect 652720 295944 652726 295956
rect 665818 295944 665824 295956
rect 665876 295944 665882 295996
rect 675496 295792 675524 296352
rect 675478 295740 675484 295792
rect 675536 295740 675542 295792
rect 35802 295604 35808 295656
rect 35860 295644 35866 295656
rect 40678 295644 40684 295656
rect 35860 295616 40684 295644
rect 35860 295604 35866 295616
rect 40678 295604 40684 295616
rect 40736 295604 40742 295656
rect 35434 295468 35440 295520
rect 35492 295508 35498 295520
rect 41322 295508 41328 295520
rect 35492 295480 41328 295508
rect 35492 295468 35498 295480
rect 41322 295468 41328 295480
rect 41380 295468 41386 295520
rect 58618 295400 58624 295452
rect 58676 295440 58682 295452
rect 62114 295440 62120 295452
rect 58676 295412 62120 295440
rect 58676 295400 58682 295412
rect 62114 295400 62120 295412
rect 62172 295400 62178 295452
rect 35618 295332 35624 295384
rect 35676 295372 35682 295384
rect 41598 295372 41604 295384
rect 35676 295344 41604 295372
rect 35676 295332 35682 295344
rect 41598 295332 41604 295344
rect 41656 295332 41662 295384
rect 35802 294108 35808 294160
rect 35860 294148 35866 294160
rect 41690 294148 41696 294160
rect 35860 294120 41696 294148
rect 35860 294108 35866 294120
rect 41690 294108 41696 294120
rect 41748 294108 41754 294160
rect 57238 294040 57244 294092
rect 57296 294080 57302 294092
rect 62114 294080 62120 294092
rect 57296 294052 62120 294080
rect 57296 294040 57302 294052
rect 62114 294040 62120 294052
rect 62172 294040 62178 294092
rect 651466 293972 651472 294024
rect 651524 294012 651530 294024
rect 664438 294012 664444 294024
rect 651524 293984 664444 294012
rect 651524 293972 651530 293984
rect 664438 293972 664444 293984
rect 664496 293972 664502 294024
rect 35802 292884 35808 292936
rect 35860 292924 35866 292936
rect 35860 292884 35894 292924
rect 35866 292856 35894 292884
rect 41506 292856 41512 292868
rect 35866 292828 41512 292856
rect 41506 292816 41512 292828
rect 41564 292816 41570 292868
rect 35802 292544 35808 292596
rect 35860 292584 35866 292596
rect 35860 292556 38654 292584
rect 35860 292544 35866 292556
rect 38626 292244 38654 292556
rect 54478 292544 54484 292596
rect 54536 292584 54542 292596
rect 62298 292584 62304 292596
rect 54536 292556 62304 292584
rect 54536 292544 54542 292556
rect 62298 292544 62304 292556
rect 62356 292544 62362 292596
rect 651466 292544 651472 292596
rect 651524 292584 651530 292596
rect 663058 292584 663064 292596
rect 651524 292556 663064 292584
rect 651524 292544 651530 292556
rect 663058 292544 663064 292556
rect 663116 292544 663122 292596
rect 42058 292408 42064 292460
rect 42116 292448 42122 292460
rect 42978 292448 42984 292460
rect 42116 292420 42984 292448
rect 42116 292408 42122 292420
rect 42978 292408 42984 292420
rect 43036 292408 43042 292460
rect 46198 292408 46204 292460
rect 46256 292448 46262 292460
rect 62114 292448 62120 292460
rect 46256 292420 62120 292448
rect 46256 292408 46262 292420
rect 62114 292408 62120 292420
rect 62172 292408 62178 292460
rect 41598 292244 41604 292256
rect 38626 292216 41604 292244
rect 41598 292204 41604 292216
rect 41656 292204 41662 292256
rect 53098 291116 53104 291168
rect 53156 291156 53162 291168
rect 62114 291156 62120 291168
rect 53156 291128 62120 291156
rect 53156 291116 53162 291128
rect 62114 291116 62120 291128
rect 62172 291116 62178 291168
rect 41690 290136 41696 290148
rect 38626 290108 41696 290136
rect 35802 289892 35808 289944
rect 35860 289932 35866 289944
rect 38626 289932 38654 290108
rect 41690 290096 41696 290108
rect 41748 290096 41754 290148
rect 35860 289904 38654 289932
rect 35860 289892 35866 289904
rect 651466 289824 651472 289876
rect 651524 289864 651530 289876
rect 660298 289864 660304 289876
rect 651524 289836 660304 289864
rect 651524 289824 651530 289836
rect 660298 289824 660304 289836
rect 660356 289824 660362 289876
rect 35618 289076 35624 289128
rect 35676 289116 35682 289128
rect 35676 289088 41414 289116
rect 35676 289076 35682 289088
rect 41386 289048 41414 289088
rect 41690 289048 41696 289060
rect 41386 289020 41696 289048
rect 41690 289008 41696 289020
rect 41748 289008 41754 289060
rect 55858 288464 55864 288516
rect 55916 288504 55922 288516
rect 62114 288504 62120 288516
rect 55916 288476 62120 288504
rect 55916 288464 55922 288476
rect 62114 288464 62120 288476
rect 62172 288464 62178 288516
rect 651466 288396 651472 288448
rect 651524 288436 651530 288448
rect 661678 288436 661684 288448
rect 651524 288408 661684 288436
rect 651524 288396 651530 288408
rect 661678 288396 661684 288408
rect 661736 288396 661742 288448
rect 651466 287036 651472 287088
rect 651524 287076 651530 287088
rect 672258 287076 672264 287088
rect 651524 287048 672264 287076
rect 651524 287036 651530 287048
rect 672258 287036 672264 287048
rect 672316 287036 672322 287088
rect 674374 286968 674380 287020
rect 674432 287008 674438 287020
rect 675110 287008 675116 287020
rect 674432 286980 675116 287008
rect 674432 286968 674438 286980
rect 675110 286968 675116 286980
rect 675168 286968 675174 287020
rect 33778 286288 33784 286340
rect 33836 286328 33842 286340
rect 41690 286328 41696 286340
rect 33836 286300 41696 286328
rect 33836 286288 33842 286300
rect 41690 286288 41696 286300
rect 41748 286288 41754 286340
rect 46198 285676 46204 285728
rect 46256 285716 46262 285728
rect 62114 285716 62120 285728
rect 46256 285688 62120 285716
rect 46256 285676 46262 285688
rect 62114 285676 62120 285688
rect 62172 285676 62178 285728
rect 651466 285676 651472 285728
rect 651524 285716 651530 285728
rect 668118 285716 668124 285728
rect 651524 285688 668124 285716
rect 651524 285676 651530 285688
rect 668118 285676 668124 285688
rect 668176 285676 668182 285728
rect 59998 284384 60004 284436
rect 60056 284424 60062 284436
rect 62114 284424 62120 284436
rect 60056 284396 62120 284424
rect 60056 284384 60062 284396
rect 62114 284384 62120 284396
rect 62172 284384 62178 284436
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 672074 284356 672080 284368
rect 651524 284328 672080 284356
rect 651524 284316 651530 284328
rect 672074 284316 672080 284328
rect 672132 284316 672138 284368
rect 47762 280304 47768 280356
rect 47820 280344 47826 280356
rect 62114 280344 62120 280356
rect 47820 280316 62120 280344
rect 47820 280304 47826 280316
rect 62114 280304 62120 280316
rect 62172 280304 62178 280356
rect 651466 280304 651472 280356
rect 651524 280344 651530 280356
rect 667198 280344 667204 280356
rect 651524 280316 667204 280344
rect 651524 280304 651530 280316
rect 667198 280304 667204 280316
rect 667256 280304 667262 280356
rect 651650 280168 651656 280220
rect 651708 280208 651714 280220
rect 667382 280208 667388 280220
rect 651708 280180 667388 280208
rect 651708 280168 651714 280180
rect 667382 280168 667388 280180
rect 667440 280168 667446 280220
rect 42242 280100 42248 280152
rect 42300 280140 42306 280152
rect 42978 280140 42984 280152
rect 42300 280112 42984 280140
rect 42300 280100 42306 280112
rect 42978 280100 42984 280112
rect 43036 280100 43042 280152
rect 482830 277312 482836 277364
rect 482888 277352 482894 277364
rect 557534 277352 557540 277364
rect 482888 277324 557540 277352
rect 482888 277312 482894 277324
rect 557534 277312 557540 277324
rect 557592 277312 557598 277364
rect 485682 277176 485688 277228
rect 485740 277216 485746 277228
rect 562318 277216 562324 277228
rect 485740 277188 562324 277216
rect 485740 277176 485746 277188
rect 562318 277176 562324 277188
rect 562376 277176 562382 277228
rect 495066 277040 495072 277092
rect 495124 277080 495130 277092
rect 576486 277080 576492 277092
rect 495124 277052 576492 277080
rect 495124 277040 495130 277052
rect 576486 277040 576492 277052
rect 576544 277040 576550 277092
rect 511626 276904 511632 276956
rect 511684 276944 511690 276956
rect 600130 276944 600136 276956
rect 511684 276916 600136 276944
rect 511684 276904 511690 276916
rect 600130 276904 600136 276916
rect 600188 276904 600194 276956
rect 514478 276768 514484 276820
rect 514536 276808 514542 276820
rect 603626 276808 603632 276820
rect 514536 276780 603632 276808
rect 514536 276768 514542 276780
rect 603626 276768 603632 276780
rect 603684 276768 603690 276820
rect 518710 276632 518716 276684
rect 518768 276672 518774 276684
rect 609606 276672 609612 276684
rect 518768 276644 609612 276672
rect 518768 276632 518774 276644
rect 609606 276632 609612 276644
rect 609664 276632 609670 276684
rect 477034 276496 477040 276548
rect 477092 276536 477098 276548
rect 550450 276536 550456 276548
rect 477092 276508 550456 276536
rect 477092 276496 477098 276508
rect 550450 276496 550456 276508
rect 550508 276496 550514 276548
rect 478506 276360 478512 276412
rect 478564 276400 478570 276412
rect 551646 276400 551652 276412
rect 478564 276372 551652 276400
rect 478564 276360 478570 276372
rect 551646 276360 551652 276372
rect 551704 276360 551710 276412
rect 471606 276224 471612 276276
rect 471664 276264 471670 276276
rect 543366 276264 543372 276276
rect 471664 276236 543372 276264
rect 471664 276224 471670 276236
rect 543366 276224 543372 276236
rect 543424 276224 543430 276276
rect 543366 276088 543372 276140
rect 543424 276128 543430 276140
rect 549254 276128 549260 276140
rect 543424 276100 549260 276128
rect 543424 276088 543430 276100
rect 549254 276088 549260 276100
rect 549312 276088 549318 276140
rect 107194 275952 107200 276004
rect 107252 275992 107258 276004
rect 162118 275992 162124 276004
rect 107252 275964 162124 275992
rect 107252 275952 107258 275964
rect 162118 275952 162124 275964
rect 162176 275952 162182 276004
rect 185210 275952 185216 276004
rect 185268 275992 185274 276004
rect 221274 275992 221280 276004
rect 185268 275964 221280 275992
rect 185268 275952 185274 275964
rect 221274 275952 221280 275964
rect 221332 275952 221338 276004
rect 454402 275952 454408 276004
rect 454460 275992 454466 276004
rect 454460 275964 454724 275992
rect 454460 275952 454466 275964
rect 100110 275816 100116 275868
rect 100168 275856 100174 275868
rect 161382 275856 161388 275868
rect 100168 275828 161388 275856
rect 100168 275816 100174 275828
rect 161382 275816 161388 275828
rect 161440 275816 161446 275868
rect 161566 275816 161572 275868
rect 161624 275816 161630 275868
rect 161750 275816 161756 275868
rect 161808 275856 161814 275868
rect 166994 275856 167000 275868
rect 161808 275828 167000 275856
rect 161808 275816 161814 275828
rect 166994 275816 167000 275828
rect 167052 275816 167058 275868
rect 178126 275816 178132 275868
rect 178184 275856 178190 275868
rect 216674 275856 216680 275868
rect 178184 275828 216680 275856
rect 178184 275816 178190 275828
rect 216674 275816 216680 275828
rect 216732 275816 216738 275868
rect 217134 275816 217140 275868
rect 217192 275856 217198 275868
rect 224034 275856 224040 275868
rect 217192 275828 224040 275856
rect 217192 275816 217198 275828
rect 224034 275816 224040 275828
rect 224092 275816 224098 275868
rect 232498 275816 232504 275868
rect 232556 275856 232562 275868
rect 239858 275856 239864 275868
rect 232556 275828 239864 275856
rect 232556 275816 232562 275828
rect 239858 275816 239864 275828
rect 239916 275816 239922 275868
rect 284570 275816 284576 275868
rect 284628 275856 284634 275868
rect 290090 275856 290096 275868
rect 284628 275828 290096 275856
rect 284628 275816 284634 275828
rect 290090 275816 290096 275828
rect 290148 275816 290154 275868
rect 445018 275816 445024 275868
rect 445076 275856 445082 275868
rect 454696 275856 454724 275964
rect 457438 275952 457444 276004
rect 457496 275992 457502 276004
rect 509050 275992 509056 276004
rect 457496 275964 509056 275992
rect 457496 275952 457502 275964
rect 509050 275952 509056 275964
rect 509108 275952 509114 276004
rect 517146 275952 517152 276004
rect 517204 275992 517210 276004
rect 608410 275992 608416 276004
rect 517204 275964 608416 275992
rect 517204 275952 517210 275964
rect 608410 275952 608416 275964
rect 608468 275952 608474 276004
rect 475378 275856 475384 275868
rect 445076 275828 454632 275856
rect 454696 275828 475384 275856
rect 445076 275816 445082 275828
rect 93026 275680 93032 275732
rect 93084 275720 93090 275732
rect 155954 275720 155960 275732
rect 93084 275692 155960 275720
rect 93084 275680 93090 275692
rect 155954 275680 155960 275692
rect 156012 275680 156018 275732
rect 161584 275720 161612 275816
rect 163130 275720 163136 275732
rect 161584 275692 163136 275720
rect 163130 275680 163136 275692
rect 163188 275680 163194 275732
rect 164050 275680 164056 275732
rect 164108 275720 164114 275732
rect 164108 275692 166488 275720
rect 164108 275680 164114 275692
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86218 275584 86224 275596
rect 76524 275556 86224 275584
rect 76524 275544 76530 275556
rect 86218 275544 86224 275556
rect 86276 275544 86282 275596
rect 90726 275544 90732 275596
rect 90784 275584 90790 275596
rect 154758 275584 154764 275596
rect 90784 275556 154764 275584
rect 90784 275544 90790 275556
rect 154758 275544 154764 275556
rect 154816 275544 154822 275596
rect 156874 275544 156880 275596
rect 156932 275584 156938 275596
rect 166460 275584 166488 275692
rect 171042 275680 171048 275732
rect 171100 275720 171106 275732
rect 211062 275720 211068 275732
rect 171100 275692 211068 275720
rect 171100 275680 171106 275692
rect 211062 275680 211068 275692
rect 211120 275680 211126 275732
rect 224218 275680 224224 275732
rect 224276 275720 224282 275732
rect 232774 275720 232780 275732
rect 224276 275692 232780 275720
rect 224276 275680 224282 275692
rect 232774 275680 232780 275692
rect 232832 275680 232838 275732
rect 236086 275680 236092 275732
rect 236144 275720 236150 275732
rect 253382 275720 253388 275732
rect 236144 275692 253388 275720
rect 236144 275680 236150 275692
rect 253382 275680 253388 275692
rect 253440 275680 253446 275732
rect 435634 275680 435640 275732
rect 435692 275720 435698 275732
rect 454402 275720 454408 275732
rect 435692 275692 454408 275720
rect 435692 275680 435698 275692
rect 454402 275680 454408 275692
rect 454460 275680 454466 275732
rect 454604 275720 454632 275828
rect 475378 275816 475384 275828
rect 475436 275816 475442 275868
rect 479518 275816 479524 275868
rect 479576 275856 479582 275868
rect 523310 275856 523316 275868
rect 479576 275828 523316 275856
rect 479576 275816 479582 275828
rect 523310 275816 523316 275828
rect 523368 275816 523374 275868
rect 524138 275816 524144 275868
rect 524196 275856 524202 275868
rect 615494 275856 615500 275868
rect 524196 275828 615500 275856
rect 524196 275816 524202 275828
rect 615494 275816 615500 275828
rect 615552 275816 615558 275868
rect 498470 275720 498476 275732
rect 454604 275692 498476 275720
rect 498470 275680 498476 275692
rect 498528 275680 498534 275732
rect 507854 275680 507860 275732
rect 507912 275720 507918 275732
rect 545758 275720 545764 275732
rect 507912 275692 545764 275720
rect 507912 275680 507918 275692
rect 545758 275680 545764 275692
rect 545816 275680 545822 275732
rect 277486 275612 277492 275664
rect 277544 275652 277550 275664
rect 284294 275652 284300 275664
rect 277544 275624 284300 275652
rect 277544 275612 277550 275624
rect 284294 275612 284300 275624
rect 284352 275612 284358 275664
rect 291654 275612 291660 275664
rect 291712 275652 291718 275664
rect 295334 275652 295340 275664
rect 291712 275624 295340 275652
rect 291712 275612 291718 275624
rect 295334 275612 295340 275624
rect 295392 275612 295398 275664
rect 206370 275584 206376 275596
rect 156932 275556 166304 275584
rect 166460 275556 206376 275584
rect 156932 275544 156938 275556
rect 81250 275408 81256 275460
rect 81308 275448 81314 275460
rect 145558 275448 145564 275460
rect 81308 275420 145564 275448
rect 81308 275408 81314 275420
rect 145558 275408 145564 275420
rect 145616 275408 145622 275460
rect 160462 275408 160468 275460
rect 160520 275448 160526 275460
rect 161842 275448 161848 275460
rect 160520 275420 161848 275448
rect 160520 275408 160526 275420
rect 161842 275408 161848 275420
rect 161900 275408 161906 275460
rect 166276 275448 166304 275556
rect 206370 275544 206376 275556
rect 206428 275544 206434 275596
rect 221918 275544 221924 275596
rect 221976 275584 221982 275596
rect 239398 275584 239404 275596
rect 221976 275556 239404 275584
rect 221976 275544 221982 275556
rect 239398 275544 239404 275556
rect 239456 275544 239462 275596
rect 243170 275544 243176 275596
rect 243228 275584 243234 275596
rect 255314 275584 255320 275596
rect 243228 275556 255320 275584
rect 243228 275544 243234 275556
rect 255314 275544 255320 275556
rect 255372 275544 255378 275596
rect 257338 275544 257344 275596
rect 257396 275584 257402 275596
rect 262858 275584 262864 275596
rect 257396 275556 262864 275584
rect 257396 275544 257402 275556
rect 262858 275544 262864 275556
rect 262916 275544 262922 275596
rect 286870 275544 286876 275596
rect 286928 275584 286934 275596
rect 286928 275556 291424 275584
rect 286928 275544 286934 275556
rect 291396 275516 291424 275556
rect 430206 275544 430212 275596
rect 430264 275584 430270 275596
rect 484302 275584 484308 275596
rect 430264 275556 484308 275584
rect 430264 275544 430270 275556
rect 484302 275544 484308 275556
rect 484360 275544 484366 275596
rect 501598 275544 501604 275596
rect 501656 275584 501662 275596
rect 512638 275584 512644 275596
rect 501656 275556 512644 275584
rect 501656 275544 501662 275556
rect 512638 275544 512644 275556
rect 512696 275544 512702 275596
rect 515398 275544 515404 275596
rect 515456 275584 515462 275596
rect 526806 275584 526812 275596
rect 515456 275556 526812 275584
rect 515456 275544 515462 275556
rect 526806 275544 526812 275556
rect 526864 275544 526870 275596
rect 528186 275544 528192 275596
rect 528244 275584 528250 275596
rect 622578 275584 622584 275596
rect 528244 275556 622584 275584
rect 528244 275544 528250 275556
rect 622578 275544 622584 275556
rect 622636 275544 622642 275596
rect 291746 275516 291752 275528
rect 291396 275488 291752 275516
rect 291746 275476 291752 275488
rect 291804 275476 291810 275528
rect 198734 275448 198740 275460
rect 166276 275420 198740 275448
rect 198734 275408 198740 275420
rect 198792 275408 198798 275460
rect 214834 275408 214840 275460
rect 214892 275448 214898 275460
rect 236638 275448 236644 275460
rect 214892 275420 236644 275448
rect 214892 275408 214898 275420
rect 236638 275408 236644 275420
rect 236696 275408 236702 275460
rect 239582 275408 239588 275460
rect 239640 275448 239646 275460
rect 251910 275448 251916 275460
rect 239640 275420 251916 275448
rect 239640 275408 239646 275420
rect 251910 275408 251916 275420
rect 251968 275408 251974 275460
rect 263226 275408 263232 275460
rect 263284 275448 263290 275460
rect 273254 275448 273260 275460
rect 263284 275420 273260 275448
rect 263284 275408 263290 275420
rect 273254 275408 273260 275420
rect 273312 275408 273318 275460
rect 285674 275408 285680 275460
rect 285732 275448 285738 275460
rect 291194 275448 291200 275460
rect 285732 275420 291200 275448
rect 285732 275408 285738 275420
rect 291194 275408 291200 275420
rect 291252 275408 291258 275460
rect 386046 275408 386052 275460
rect 386104 275448 386110 275460
rect 420454 275448 420460 275460
rect 386104 275420 420460 275448
rect 386104 275408 386110 275420
rect 420454 275408 420460 275420
rect 420512 275408 420518 275460
rect 423398 275408 423404 275460
rect 423456 275448 423462 275460
rect 473354 275448 473360 275460
rect 423456 275420 473360 275448
rect 423456 275408 423462 275420
rect 473354 275408 473360 275420
rect 473412 275408 473418 275460
rect 475378 275408 475384 275460
rect 475436 275448 475442 275460
rect 485038 275448 485044 275460
rect 475436 275420 485044 275448
rect 475436 275408 475442 275420
rect 485038 275408 485044 275420
rect 485096 275408 485102 275460
rect 485222 275408 485228 275460
rect 485280 275448 485286 275460
rect 537478 275448 537484 275460
rect 485280 275420 537484 275448
rect 485280 275408 485286 275420
rect 537478 275408 537484 275420
rect 537536 275408 537542 275460
rect 636746 275448 636752 275460
rect 537772 275420 636752 275448
rect 299934 275340 299940 275392
rect 299992 275380 299998 275392
rect 301222 275380 301228 275392
rect 299992 275352 301228 275380
rect 299992 275340 299998 275352
rect 301222 275340 301228 275352
rect 301280 275340 301286 275392
rect 71774 275272 71780 275324
rect 71832 275312 71838 275324
rect 141050 275312 141056 275324
rect 71832 275284 141056 275312
rect 71832 275272 71838 275284
rect 141050 275272 141056 275284
rect 141108 275272 141114 275324
rect 146202 275272 146208 275324
rect 146260 275312 146266 275324
rect 189074 275312 189080 275324
rect 146260 275284 189080 275312
rect 146260 275272 146266 275284
rect 189074 275272 189080 275284
rect 189132 275272 189138 275324
rect 218330 275272 218336 275324
rect 218388 275312 218394 275324
rect 243078 275312 243084 275324
rect 218388 275284 243084 275312
rect 218388 275272 218394 275284
rect 243078 275272 243084 275284
rect 243136 275272 243142 275324
rect 256142 275272 256148 275324
rect 256200 275312 256206 275324
rect 268838 275312 268844 275324
rect 256200 275284 268844 275312
rect 256200 275272 256206 275284
rect 268838 275272 268844 275284
rect 268896 275272 268902 275324
rect 273898 275272 273904 275324
rect 273956 275312 273962 275324
rect 282914 275312 282920 275324
rect 273956 275284 282920 275312
rect 273956 275272 273962 275284
rect 282914 275272 282920 275284
rect 282972 275272 282978 275324
rect 290458 275272 290464 275324
rect 290516 275312 290522 275324
rect 294138 275312 294144 275324
rect 290516 275284 294144 275312
rect 290516 275272 290522 275284
rect 294138 275272 294144 275284
rect 294196 275272 294202 275324
rect 361206 275272 361212 275324
rect 361264 275312 361270 275324
rect 385034 275312 385040 275324
rect 361264 275284 385040 275312
rect 361264 275272 361270 275284
rect 385034 275272 385040 275284
rect 385092 275272 385098 275324
rect 416406 275272 416412 275324
rect 416464 275312 416470 275324
rect 462958 275312 462964 275324
rect 416464 275284 462964 275312
rect 416464 275272 416470 275284
rect 462958 275272 462964 275284
rect 463016 275272 463022 275324
rect 463142 275272 463148 275324
rect 463200 275312 463206 275324
rect 530394 275312 530400 275324
rect 463200 275284 530400 275312
rect 463200 275272 463206 275284
rect 530394 275272 530400 275284
rect 530452 275272 530458 275324
rect 532326 275272 532332 275324
rect 532384 275312 532390 275324
rect 537294 275312 537300 275324
rect 532384 275284 537300 275312
rect 532384 275272 532390 275284
rect 537294 275272 537300 275284
rect 537352 275272 537358 275324
rect 537570 275272 537576 275324
rect 537628 275312 537634 275324
rect 537772 275312 537800 275420
rect 636746 275408 636752 275420
rect 636804 275408 636810 275460
rect 537628 275284 537800 275312
rect 537628 275272 537634 275284
rect 537938 275272 537944 275324
rect 537996 275312 538002 275324
rect 540974 275312 540980 275324
rect 537996 275284 540980 275312
rect 537996 275272 538002 275284
rect 540974 275272 540980 275284
rect 541032 275272 541038 275324
rect 542998 275272 543004 275324
rect 543056 275312 543062 275324
rect 629662 275312 629668 275324
rect 543056 275284 629668 275312
rect 543056 275272 543062 275284
rect 629662 275272 629668 275284
rect 629720 275272 629726 275324
rect 298738 275204 298744 275256
rect 298796 275244 298802 275256
rect 300026 275244 300032 275256
rect 298796 275216 300032 275244
rect 298796 275204 298802 275216
rect 300026 275204 300032 275216
rect 300084 275204 300090 275256
rect 139118 275136 139124 275188
rect 139176 275176 139182 275188
rect 146938 275176 146944 275188
rect 139176 275148 146944 275176
rect 139176 275136 139182 275148
rect 146938 275136 146944 275148
rect 146996 275136 147002 275188
rect 149790 275136 149796 275188
rect 149848 275176 149854 275188
rect 191742 275176 191748 275188
rect 149848 275148 191748 275176
rect 149848 275136 149854 275148
rect 191742 275136 191748 275148
rect 191800 275136 191806 275188
rect 292850 275136 292856 275188
rect 292908 275176 292914 275188
rect 295794 275176 295800 275188
rect 292908 275148 295800 275176
rect 292908 275136 292914 275148
rect 295794 275136 295800 275148
rect 295852 275136 295858 275188
rect 427078 275136 427084 275188
rect 427136 275176 427142 275188
rect 477218 275176 477224 275188
rect 427136 275148 477224 275176
rect 427136 275136 427142 275148
rect 477218 275136 477224 275148
rect 477276 275136 477282 275188
rect 485038 275136 485044 275188
rect 485096 275176 485102 275188
rect 491386 275176 491392 275188
rect 485096 275148 491392 275176
rect 485096 275136 485102 275148
rect 491386 275136 491392 275148
rect 491444 275136 491450 275188
rect 493318 275136 493324 275188
rect 493376 275176 493382 275188
rect 493376 275148 495112 275176
rect 493376 275136 493382 275148
rect 269206 275068 269212 275120
rect 269264 275108 269270 275120
rect 274910 275108 274916 275120
rect 269264 275080 274916 275108
rect 269264 275068 269270 275080
rect 274910 275068 274916 275080
rect 274968 275068 274974 275120
rect 110782 275000 110788 275052
rect 110840 275040 110846 275052
rect 149698 275040 149704 275052
rect 110840 275012 149704 275040
rect 110840 275000 110846 275012
rect 149698 275000 149704 275012
rect 149756 275000 149762 275052
rect 153378 275000 153384 275052
rect 153436 275040 153442 275052
rect 154482 275040 154488 275052
rect 153436 275012 154488 275040
rect 153436 275000 153442 275012
rect 154482 275000 154488 275012
rect 154540 275000 154546 275052
rect 161658 275040 161664 275052
rect 161446 275012 161664 275040
rect 132034 274864 132040 274916
rect 132092 274904 132098 274916
rect 161446 274904 161474 275012
rect 161658 275000 161664 275012
rect 161716 275000 161722 275052
rect 161842 275000 161848 275052
rect 161900 275040 161906 275052
rect 175918 275040 175924 275052
rect 161900 275012 175924 275040
rect 161900 275000 161906 275012
rect 175918 275000 175924 275012
rect 175976 275000 175982 275052
rect 189994 275000 190000 275052
rect 190052 275040 190058 275052
rect 218698 275040 218704 275052
rect 190052 275012 218704 275040
rect 190052 275000 190058 275012
rect 218698 275000 218704 275012
rect 218756 275000 218762 275052
rect 288066 275000 288072 275052
rect 288124 275040 288130 275052
rect 292666 275040 292672 275052
rect 288124 275012 292672 275040
rect 288124 275000 288130 275012
rect 292666 275000 292672 275012
rect 292724 275000 292730 275052
rect 420638 275000 420644 275052
rect 420696 275040 420702 275052
rect 470134 275040 470140 275052
rect 420696 275012 470140 275040
rect 420696 275000 420702 275012
rect 470134 275000 470140 275012
rect 470192 275000 470198 275052
rect 476114 275000 476120 275052
rect 476172 275040 476178 275052
rect 485222 275040 485228 275052
rect 476172 275012 485228 275040
rect 476172 275000 476178 275012
rect 485222 275000 485228 275012
rect 485280 275000 485286 275052
rect 492398 275000 492404 275052
rect 492456 275040 492462 275052
rect 494882 275040 494888 275052
rect 492456 275012 494888 275040
rect 492456 275000 492462 275012
rect 494882 275000 494888 275012
rect 494940 275000 494946 275052
rect 495084 275040 495112 275148
rect 497458 275136 497464 275188
rect 497516 275176 497522 275188
rect 505554 275176 505560 275188
rect 497516 275148 505560 275176
rect 497516 275136 497522 275148
rect 505554 275136 505560 275148
rect 505612 275136 505618 275188
rect 507486 275136 507492 275188
rect 507544 275176 507550 275188
rect 594242 275176 594248 275188
rect 507544 275148 594248 275176
rect 507544 275136 507550 275148
rect 594242 275136 594248 275148
rect 594300 275136 594306 275188
rect 501966 275040 501972 275052
rect 495084 275012 501972 275040
rect 501966 275000 501972 275012
rect 502024 275000 502030 275052
rect 503438 275000 503444 275052
rect 503496 275040 503502 275052
rect 587066 275040 587072 275052
rect 503496 275012 587072 275040
rect 503496 275000 503502 275012
rect 587066 275000 587072 275012
rect 587124 275000 587130 275052
rect 293954 274932 293960 274984
rect 294012 274972 294018 274984
rect 297174 274972 297180 274984
rect 294012 274944 297180 274972
rect 294012 274932 294018 274944
rect 297174 274932 297180 274944
rect 297232 274932 297238 274984
rect 132092 274876 161474 274904
rect 132092 274864 132098 274876
rect 167546 274864 167552 274916
rect 167604 274904 167610 274916
rect 169018 274904 169024 274916
rect 167604 274876 169024 274904
rect 167604 274864 167610 274876
rect 169018 274864 169024 274876
rect 169076 274864 169082 274916
rect 413462 274864 413468 274916
rect 413520 274904 413526 274916
rect 459462 274904 459468 274916
rect 413520 274876 459468 274904
rect 413520 274864 413526 274876
rect 459462 274864 459468 274876
rect 459520 274864 459526 274916
rect 473354 274864 473360 274916
rect 473412 274904 473418 274916
rect 544562 274904 544568 274916
rect 473412 274876 544568 274904
rect 473412 274864 473418 274876
rect 544562 274864 544568 274876
rect 544620 274864 544626 274916
rect 174630 274796 174636 274848
rect 174688 274836 174694 274848
rect 182726 274836 182732 274848
rect 174688 274808 182732 274836
rect 174688 274796 174694 274808
rect 182726 274796 182732 274808
rect 182784 274796 182790 274848
rect 289262 274796 289268 274848
rect 289320 274836 289326 274848
rect 293402 274836 293408 274848
rect 289320 274808 293408 274836
rect 289320 274796 289326 274808
rect 293402 274796 293408 274808
rect 293460 274796 293466 274848
rect 296346 274796 296352 274848
rect 296404 274836 296410 274848
rect 298370 274836 298376 274848
rect 296404 274808 298376 274836
rect 296404 274796 296410 274808
rect 298370 274796 298376 274808
rect 298428 274796 298434 274848
rect 553366 274808 557534 274836
rect 136818 274728 136824 274780
rect 136876 274768 136882 274780
rect 137646 274768 137652 274780
rect 136876 274740 137652 274768
rect 136876 274728 136882 274740
rect 137646 274728 137652 274740
rect 137704 274728 137710 274780
rect 143902 274728 143908 274780
rect 143960 274768 143966 274780
rect 144362 274768 144368 274780
rect 143960 274740 144368 274768
rect 143960 274728 143966 274740
rect 144362 274728 144368 274740
rect 144420 274728 144426 274780
rect 146938 274728 146944 274780
rect 146996 274768 147002 274780
rect 174446 274768 174452 274780
rect 146996 274740 174452 274768
rect 146996 274728 147002 274740
rect 174446 274728 174452 274740
rect 174504 274728 174510 274780
rect 469858 274728 469864 274780
rect 469916 274768 469922 274780
rect 516226 274768 516232 274780
rect 469916 274740 516232 274768
rect 469916 274728 469922 274740
rect 516226 274728 516232 274740
rect 516284 274728 516290 274780
rect 526438 274728 526444 274780
rect 526496 274768 526502 274780
rect 533890 274768 533896 274780
rect 526496 274740 533896 274768
rect 526496 274728 526502 274740
rect 533890 274728 533896 274740
rect 533948 274728 533954 274780
rect 534718 274728 534724 274780
rect 534776 274768 534782 274780
rect 537938 274768 537944 274780
rect 534776 274740 537944 274768
rect 534776 274728 534782 274740
rect 537938 274728 537944 274740
rect 537996 274728 538002 274780
rect 538122 274728 538128 274780
rect 538180 274768 538186 274780
rect 542998 274768 543004 274780
rect 538180 274740 543004 274768
rect 538180 274728 538186 274740
rect 542998 274728 543004 274740
rect 543056 274728 543062 274780
rect 543182 274728 543188 274780
rect 543240 274768 543246 274780
rect 553366 274768 553394 274808
rect 543240 274740 553394 274768
rect 557506 274768 557534 274808
rect 643830 274768 643836 274780
rect 557506 274740 643836 274768
rect 543240 274728 543246 274740
rect 643830 274728 643836 274740
rect 643888 274728 643894 274780
rect 74166 274660 74172 274712
rect 74224 274700 74230 274712
rect 76742 274700 76748 274712
rect 74224 274672 76748 274700
rect 74224 274660 74230 274672
rect 76742 274660 76748 274672
rect 76800 274660 76806 274712
rect 85942 274660 85948 274712
rect 86000 274700 86006 274712
rect 90358 274700 90364 274712
rect 86000 274672 90364 274700
rect 86000 274660 86006 274672
rect 90358 274660 90364 274672
rect 90416 274660 90422 274712
rect 103698 274660 103704 274712
rect 103756 274700 103762 274712
rect 104802 274700 104808 274712
rect 103756 274672 104808 274700
rect 103756 274660 103762 274672
rect 104802 274660 104808 274672
rect 104860 274660 104866 274712
rect 253842 274660 253848 274712
rect 253900 274700 253906 274712
rect 258350 274700 258356 274712
rect 253900 274672 258356 274700
rect 253900 274660 253906 274672
rect 258350 274660 258356 274672
rect 258408 274660 258414 274712
rect 268010 274660 268016 274712
rect 268068 274700 268074 274712
rect 272426 274700 272432 274712
rect 268068 274672 272432 274700
rect 268068 274660 268074 274672
rect 272426 274660 272432 274672
rect 272484 274660 272490 274712
rect 283374 274660 283380 274712
rect 283432 274700 283438 274712
rect 289170 274700 289176 274712
rect 283432 274672 289176 274700
rect 283432 274660 283438 274672
rect 289170 274660 289176 274672
rect 289228 274660 289234 274712
rect 295150 274660 295156 274712
rect 295208 274700 295214 274712
rect 296806 274700 296812 274712
rect 295208 274672 296812 274700
rect 295208 274660 295214 274672
rect 296806 274660 296812 274672
rect 296864 274660 296870 274712
rect 297542 274660 297548 274712
rect 297600 274700 297606 274712
rect 299566 274700 299572 274712
rect 297600 274672 299572 274700
rect 297600 274660 297606 274672
rect 299566 274660 299572 274672
rect 299624 274660 299630 274712
rect 303430 274660 303436 274712
rect 303488 274700 303494 274712
rect 303982 274700 303988 274712
rect 303488 274672 303988 274700
rect 303488 274660 303494 274672
rect 303982 274660 303988 274672
rect 304040 274660 304046 274712
rect 321186 274660 321192 274712
rect 321244 274700 321250 274712
rect 328270 274700 328276 274712
rect 321244 274672 328276 274700
rect 321244 274660 321250 274672
rect 328270 274660 328276 274672
rect 328328 274660 328334 274712
rect 350718 274660 350724 274712
rect 350776 274700 350782 274712
rect 353110 274700 353116 274712
rect 350776 274672 353116 274700
rect 350776 274660 350782 274672
rect 353110 274660 353116 274672
rect 353168 274660 353174 274712
rect 113450 274592 113456 274644
rect 113508 274632 113514 274644
rect 169938 274632 169944 274644
rect 113508 274604 169944 274632
rect 113508 274592 113514 274604
rect 169938 274592 169944 274604
rect 169996 274592 170002 274644
rect 182910 274592 182916 274644
rect 182968 274632 182974 274644
rect 214558 274632 214564 274644
rect 182968 274604 214564 274632
rect 182968 274592 182974 274604
rect 214558 274592 214564 274604
rect 214616 274592 214622 274644
rect 382918 274592 382924 274644
rect 382976 274632 382982 274644
rect 392118 274632 392124 274644
rect 382976 274604 392124 274632
rect 382976 274592 382982 274604
rect 392118 274592 392124 274604
rect 392176 274592 392182 274644
rect 404170 274592 404176 274644
rect 404228 274632 404234 274644
rect 446490 274632 446496 274644
rect 404228 274604 446496 274632
rect 404228 274592 404234 274604
rect 446490 274592 446496 274604
rect 446548 274592 446554 274644
rect 450538 274592 450544 274644
rect 450596 274632 450602 274644
rect 480714 274632 480720 274644
rect 450596 274604 480720 274632
rect 450596 274592 450602 274604
rect 480714 274592 480720 274604
rect 480772 274592 480778 274644
rect 488350 274592 488356 274644
rect 488408 274632 488414 274644
rect 567010 274632 567016 274644
rect 488408 274604 567016 274632
rect 488408 274592 488414 274604
rect 567010 274592 567016 274604
rect 567068 274592 567074 274644
rect 95878 274496 95884 274508
rect 84166 274468 95884 274496
rect 67082 274320 67088 274372
rect 67140 274360 67146 274372
rect 84166 274360 84194 274468
rect 95878 274456 95884 274468
rect 95936 274456 95942 274508
rect 105170 274456 105176 274508
rect 105228 274496 105234 274508
rect 163314 274496 163320 274508
rect 105228 274468 163320 274496
rect 105228 274456 105234 274468
rect 163314 274456 163320 274468
rect 163372 274456 163378 274508
rect 168742 274456 168748 274508
rect 168800 274496 168806 274508
rect 208486 274496 208492 274508
rect 168800 274468 208492 274496
rect 168800 274456 168806 274468
rect 208486 274456 208492 274468
rect 208544 274456 208550 274508
rect 227806 274456 227812 274508
rect 227864 274496 227870 274508
rect 248874 274496 248880 274508
rect 227864 274468 248880 274496
rect 227864 274456 227870 274468
rect 248874 274456 248880 274468
rect 248932 274456 248938 274508
rect 358078 274456 358084 274508
rect 358136 274496 358142 274508
rect 369578 274496 369584 274508
rect 358136 274468 369584 274496
rect 358136 274456 358142 274468
rect 369578 274456 369584 274468
rect 369636 274456 369642 274508
rect 395614 274496 395620 274508
rect 371620 274468 395620 274496
rect 67140 274332 84194 274360
rect 67140 274320 67146 274332
rect 95418 274320 95424 274372
rect 95476 274360 95482 274372
rect 157610 274360 157616 274372
rect 95476 274332 157616 274360
rect 95476 274320 95482 274332
rect 157610 274320 157616 274332
rect 157668 274320 157674 274372
rect 166350 274320 166356 274372
rect 166408 274360 166414 274372
rect 207290 274360 207296 274372
rect 166408 274332 207296 274360
rect 166408 274320 166414 274332
rect 207290 274320 207296 274332
rect 207348 274320 207354 274372
rect 207750 274320 207756 274372
rect 207808 274360 207814 274372
rect 233878 274360 233884 274372
rect 207808 274332 233884 274360
rect 207808 274320 207814 274332
rect 233878 274320 233884 274332
rect 233936 274320 233942 274372
rect 249058 274320 249064 274372
rect 249116 274360 249122 274372
rect 265250 274360 265256 274372
rect 249116 274332 265256 274360
rect 249116 274320 249122 274332
rect 265250 274320 265256 274332
rect 265308 274320 265314 274372
rect 333790 274320 333796 274372
rect 333848 274360 333854 274372
rect 345934 274360 345940 274372
rect 333848 274332 345940 274360
rect 333848 274320 333854 274332
rect 345934 274320 345940 274332
rect 345992 274320 345998 274372
rect 347038 274320 347044 274372
rect 347096 274360 347102 274372
rect 358998 274360 359004 274372
rect 347096 274332 359004 274360
rect 347096 274320 347102 274332
rect 358998 274320 359004 274332
rect 359056 274320 359062 274372
rect 369118 274320 369124 274372
rect 369176 274360 369182 274372
rect 371620 274360 371648 274468
rect 395614 274456 395620 274468
rect 395672 274456 395678 274508
rect 409230 274456 409236 274508
rect 409288 274496 409294 274508
rect 453574 274496 453580 274508
rect 409288 274468 453580 274496
rect 409288 274456 409294 274468
rect 453574 274456 453580 274468
rect 453632 274456 453638 274508
rect 453758 274456 453764 274508
rect 453816 274496 453822 274508
rect 486602 274496 486608 274508
rect 453816 274468 486608 274496
rect 453816 274456 453822 274468
rect 486602 274456 486608 274468
rect 486660 274456 486666 274508
rect 536742 274456 536748 274508
rect 536800 274496 536806 274508
rect 543688 274496 543694 274508
rect 536800 274468 543694 274496
rect 536800 274456 536806 274468
rect 543688 274456 543694 274468
rect 543746 274456 543752 274508
rect 543826 274456 543832 274508
rect 543884 274496 543890 274508
rect 639138 274496 639144 274508
rect 543884 274468 639144 274496
rect 543884 274456 543890 274468
rect 639138 274456 639144 274468
rect 639196 274456 639202 274508
rect 369176 274332 371648 274360
rect 369176 274320 369182 274332
rect 373258 274320 373264 274372
rect 373316 274360 373322 274372
rect 400306 274360 400312 274372
rect 373316 274332 400312 274360
rect 373316 274320 373322 274332
rect 400306 274320 400312 274332
rect 400364 274320 400370 274372
rect 413830 274320 413836 274372
rect 413888 274360 413894 274372
rect 460658 274360 460664 274372
rect 413888 274332 460664 274360
rect 413888 274320 413894 274332
rect 460658 274320 460664 274332
rect 460716 274320 460722 274372
rect 465718 274320 465724 274372
rect 465776 274360 465782 274372
rect 487798 274360 487804 274372
rect 465776 274332 487804 274360
rect 465776 274320 465782 274332
rect 487798 274320 487804 274332
rect 487856 274320 487862 274372
rect 508590 274320 508596 274372
rect 508648 274360 508654 274372
rect 595070 274360 595076 274372
rect 508648 274332 595076 274360
rect 508648 274320 508654 274332
rect 595070 274320 595076 274332
rect 595128 274320 595134 274372
rect 595438 274320 595444 274372
rect 595496 274360 595502 274372
rect 640334 274360 640340 274372
rect 595496 274332 640340 274360
rect 595496 274320 595502 274332
rect 640334 274320 640340 274332
rect 640392 274320 640398 274372
rect 282178 274252 282184 274304
rect 282236 274292 282242 274304
rect 287698 274292 287704 274304
rect 282236 274264 287704 274292
rect 282236 274252 282242 274264
rect 287698 274252 287704 274264
rect 287756 274252 287762 274304
rect 89438 274184 89444 274236
rect 89496 274224 89502 274236
rect 151998 274224 152004 274236
rect 89496 274196 152004 274224
rect 89496 274184 89502 274196
rect 151998 274184 152004 274196
rect 152056 274184 152062 274236
rect 155678 274184 155684 274236
rect 155736 274224 155742 274236
rect 200114 274224 200120 274236
rect 155736 274196 200120 274224
rect 155736 274184 155742 274196
rect 200114 274184 200120 274196
rect 200172 274184 200178 274236
rect 205358 274184 205364 274236
rect 205416 274224 205422 274236
rect 234706 274224 234712 274236
rect 205416 274196 234712 274224
rect 205416 274184 205422 274196
rect 234706 274184 234712 274196
rect 234764 274184 234770 274236
rect 234890 274184 234896 274236
rect 234948 274224 234954 274236
rect 234948 274196 251956 274224
rect 234948 274184 234954 274196
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 144914 274088 144920 274100
rect 77720 274060 144920 274088
rect 77720 274048 77726 274060
rect 144914 274048 144920 274060
rect 144972 274048 144978 274100
rect 147398 274048 147404 274100
rect 147456 274088 147462 274100
rect 193398 274088 193404 274100
rect 147456 274060 193404 274088
rect 147456 274048 147462 274060
rect 193398 274048 193404 274060
rect 193456 274048 193462 274100
rect 198274 274048 198280 274100
rect 198332 274088 198338 274100
rect 229186 274088 229192 274100
rect 198332 274060 229192 274088
rect 198332 274048 198338 274060
rect 229186 274048 229192 274060
rect 229244 274048 229250 274100
rect 237282 274048 237288 274100
rect 237340 274088 237346 274100
rect 251928 274088 251956 274196
rect 255314 274184 255320 274236
rect 255372 274224 255378 274236
rect 261018 274224 261024 274236
rect 255372 274196 261024 274224
rect 255372 274184 255378 274196
rect 261018 274184 261024 274196
rect 261076 274184 261082 274236
rect 325326 274184 325332 274236
rect 325384 274224 325390 274236
rect 332962 274224 332968 274236
rect 325384 274196 332968 274224
rect 325384 274184 325390 274196
rect 332962 274184 332968 274196
rect 333020 274184 333026 274236
rect 343450 274184 343456 274236
rect 343508 274224 343514 274236
rect 360194 274224 360200 274236
rect 343508 274196 360200 274224
rect 343508 274184 343514 274196
rect 360194 274184 360200 274196
rect 360252 274184 360258 274236
rect 364978 274184 364984 274236
rect 365036 274224 365042 274236
rect 374362 274224 374368 274236
rect 365036 274196 374368 274224
rect 365036 274184 365042 274196
rect 374362 274184 374368 274196
rect 374420 274184 374426 274236
rect 379330 274184 379336 274236
rect 379388 274224 379394 274236
rect 410978 274224 410984 274236
rect 379388 274196 410984 274224
rect 379388 274184 379394 274196
rect 410978 274184 410984 274196
rect 411036 274184 411042 274236
rect 416590 274184 416596 274236
rect 416648 274224 416654 274236
rect 464154 274224 464160 274236
rect 416648 274196 464160 274224
rect 416648 274184 416654 274196
rect 464154 274184 464160 274196
rect 464212 274184 464218 274236
rect 474642 274184 474648 274236
rect 474700 274224 474706 274236
rect 507854 274224 507860 274236
rect 474700 274196 507860 274224
rect 474700 274184 474706 274196
rect 507854 274184 507860 274196
rect 507912 274184 507918 274236
rect 511810 274184 511816 274236
rect 511868 274224 511874 274236
rect 598934 274224 598940 274236
rect 511868 274196 598940 274224
rect 511868 274184 511874 274196
rect 598934 274184 598940 274196
rect 598992 274184 598998 274236
rect 255406 274088 255412 274100
rect 237340 274060 251864 274088
rect 251928 274060 255412 274088
rect 237340 274048 237346 274060
rect 65886 273912 65892 273964
rect 65944 273952 65950 273964
rect 136818 273952 136824 273964
rect 65944 273924 136824 273952
rect 65944 273912 65950 273924
rect 136818 273912 136824 273924
rect 136876 273912 136882 273964
rect 145098 273912 145104 273964
rect 145156 273952 145162 273964
rect 192386 273952 192392 273964
rect 145156 273924 192392 273952
rect 145156 273912 145162 273924
rect 192386 273912 192392 273924
rect 192444 273912 192450 273964
rect 195882 273912 195888 273964
rect 195940 273952 195946 273964
rect 227898 273952 227904 273964
rect 195940 273924 227904 273952
rect 195940 273912 195946 273924
rect 227898 273912 227904 273924
rect 227956 273912 227962 273964
rect 229002 273912 229008 273964
rect 229060 273952 229066 273964
rect 250438 273952 250444 273964
rect 229060 273924 250444 273952
rect 229060 273912 229066 273924
rect 250438 273912 250444 273924
rect 250496 273912 250502 273964
rect 251836 273952 251864 274060
rect 255406 274048 255412 274060
rect 255464 274048 255470 274100
rect 261202 274048 261208 274100
rect 261260 274088 261266 274100
rect 273530 274088 273536 274100
rect 261260 274060 273536 274088
rect 261260 274048 261266 274060
rect 273530 274048 273536 274060
rect 273588 274048 273594 274100
rect 275094 274048 275100 274100
rect 275152 274088 275158 274100
rect 283466 274088 283472 274100
rect 275152 274060 283472 274088
rect 275152 274048 275158 274060
rect 283466 274048 283472 274060
rect 283524 274048 283530 274100
rect 332318 274048 332324 274100
rect 332376 274088 332382 274100
rect 343634 274088 343640 274100
rect 332376 274060 343640 274088
rect 332376 274048 332382 274060
rect 343634 274048 343640 274060
rect 343692 274048 343698 274100
rect 350350 274048 350356 274100
rect 350408 274088 350414 274100
rect 368474 274088 368480 274100
rect 350408 274060 368480 274088
rect 350408 274048 350414 274060
rect 368474 274048 368480 274060
rect 368532 274048 368538 274100
rect 369302 274048 369308 274100
rect 369360 274088 369366 274100
rect 387334 274088 387340 274100
rect 369360 274060 387340 274088
rect 369360 274048 369366 274060
rect 387334 274048 387340 274060
rect 387392 274048 387398 274100
rect 394326 274048 394332 274100
rect 394384 274088 394390 274100
rect 432230 274088 432236 274100
rect 394384 274060 432236 274088
rect 394384 274048 394390 274060
rect 432230 274048 432236 274060
rect 432288 274048 432294 274100
rect 432598 274048 432604 274100
rect 432656 274088 432662 274100
rect 485498 274088 485504 274100
rect 432656 274060 485504 274088
rect 432656 274048 432662 274060
rect 485498 274048 485504 274060
rect 485556 274048 485562 274100
rect 491202 274048 491208 274100
rect 491260 274088 491266 274100
rect 569954 274088 569960 274100
rect 491260 274060 569960 274088
rect 491260 274048 491266 274060
rect 569954 274048 569960 274060
rect 570012 274048 570018 274100
rect 571794 274048 571800 274100
rect 571852 274088 571858 274100
rect 583570 274088 583576 274100
rect 571852 274060 583576 274088
rect 571852 274048 571858 274060
rect 583570 274048 583576 274060
rect 583628 274048 583634 274100
rect 256970 273952 256976 273964
rect 251836 273924 256976 273952
rect 256970 273912 256976 273924
rect 257028 273912 257034 273964
rect 258534 273912 258540 273964
rect 258592 273952 258598 273964
rect 272058 273952 272064 273964
rect 258592 273924 272064 273952
rect 258592 273912 258598 273924
rect 272058 273912 272064 273924
rect 272116 273912 272122 273964
rect 272702 273912 272708 273964
rect 272760 273952 272766 273964
rect 281810 273952 281816 273964
rect 272760 273924 281816 273952
rect 272760 273912 272766 273924
rect 281810 273912 281816 273924
rect 281868 273912 281874 273964
rect 324038 273912 324044 273964
rect 324096 273952 324102 273964
rect 331766 273952 331772 273964
rect 324096 273924 331772 273952
rect 324096 273912 324102 273924
rect 331766 273912 331772 273924
rect 331824 273912 331830 273964
rect 331950 273912 331956 273964
rect 332008 273952 332014 273964
rect 341242 273952 341248 273964
rect 332008 273924 341248 273952
rect 332008 273912 332014 273924
rect 341242 273912 341248 273924
rect 341300 273912 341306 273964
rect 342070 273912 342076 273964
rect 342128 273952 342134 273964
rect 357802 273952 357808 273964
rect 342128 273924 357808 273952
rect 342128 273912 342134 273924
rect 357802 273912 357808 273924
rect 357860 273912 357866 273964
rect 360102 273912 360108 273964
rect 360160 273952 360166 273964
rect 382642 273952 382648 273964
rect 360160 273924 382648 273952
rect 360160 273912 360166 273924
rect 382642 273912 382648 273924
rect 382700 273912 382706 273964
rect 387426 273912 387432 273964
rect 387484 273952 387490 273964
rect 421650 273952 421656 273964
rect 387484 273924 421656 273952
rect 387484 273912 387490 273924
rect 421650 273912 421656 273924
rect 421708 273912 421714 273964
rect 421834 273912 421840 273964
rect 421892 273952 421898 273964
rect 471238 273952 471244 273964
rect 421892 273924 471244 273952
rect 421892 273912 421898 273924
rect 471238 273912 471244 273924
rect 471296 273912 471302 273964
rect 475746 273912 475752 273964
rect 475804 273952 475810 273964
rect 543366 273952 543372 273964
rect 475804 273924 543372 273952
rect 475804 273912 475810 273924
rect 543366 273912 543372 273924
rect 543424 273912 543430 273964
rect 543826 273912 543832 273964
rect 543884 273952 543890 273964
rect 634354 273952 634360 273964
rect 543884 273924 634360 273952
rect 543884 273912 543890 273924
rect 634354 273912 634360 273924
rect 634412 273912 634418 273964
rect 96614 273776 96620 273828
rect 96672 273816 96678 273828
rect 117958 273816 117964 273828
rect 96672 273788 117964 273816
rect 96672 273776 96678 273788
rect 117958 273776 117964 273788
rect 118016 273776 118022 273828
rect 118234 273776 118240 273828
rect 118292 273816 118298 273828
rect 174170 273816 174176 273828
rect 118292 273788 174176 273816
rect 118292 273776 118298 273788
rect 174170 273776 174176 273788
rect 174228 273776 174234 273828
rect 175918 273776 175924 273828
rect 175976 273816 175982 273828
rect 204254 273816 204260 273828
rect 175976 273788 204260 273816
rect 175976 273776 175982 273788
rect 204254 273776 204260 273788
rect 204312 273776 204318 273828
rect 206554 273776 206560 273828
rect 206612 273816 206618 273828
rect 235442 273816 235448 273828
rect 206612 273788 235448 273816
rect 206612 273776 206618 273788
rect 235442 273776 235448 273788
rect 235500 273776 235506 273828
rect 400030 273776 400036 273828
rect 400088 273816 400094 273828
rect 439314 273816 439320 273828
rect 400088 273788 439320 273816
rect 400088 273776 400094 273788
rect 439314 273776 439320 273788
rect 439372 273776 439378 273828
rect 442258 273776 442264 273828
rect 442316 273816 442322 273828
rect 481910 273816 481916 273828
rect 442316 273788 481916 273816
rect 442316 273776 442322 273788
rect 481910 273776 481916 273788
rect 481968 273776 481974 273828
rect 487062 273776 487068 273828
rect 487120 273816 487126 273828
rect 560294 273816 560300 273828
rect 487120 273788 560300 273816
rect 487120 273776 487126 273788
rect 560294 273776 560300 273788
rect 560352 273776 560358 273828
rect 571794 273816 571800 273828
rect 562336 273788 571800 273816
rect 123754 273640 123760 273692
rect 123812 273680 123818 273692
rect 177482 273680 177488 273692
rect 123812 273652 177488 273680
rect 123812 273640 123818 273652
rect 177482 273640 177488 273652
rect 177540 273640 177546 273692
rect 392578 273640 392584 273692
rect 392636 273680 392642 273692
rect 409782 273680 409788 273692
rect 392636 273652 409788 273680
rect 392636 273640 392642 273652
rect 409782 273640 409788 273652
rect 409840 273640 409846 273692
rect 440878 273640 440884 273692
rect 440936 273680 440942 273692
rect 474826 273680 474832 273692
rect 440936 273652 474832 273680
rect 440936 273640 440942 273652
rect 474826 273640 474832 273652
rect 474884 273640 474890 273692
rect 481358 273640 481364 273692
rect 481416 273680 481422 273692
rect 556338 273680 556344 273692
rect 481416 273652 556344 273680
rect 481416 273640 481422 273652
rect 556338 273640 556344 273652
rect 556396 273640 556402 273692
rect 562336 273680 562364 273788
rect 571794 273776 571800 273788
rect 571852 273776 571858 273828
rect 571978 273776 571984 273828
rect 572036 273816 572042 273828
rect 597738 273816 597744 273828
rect 572036 273788 597744 273816
rect 572036 273776 572042 273788
rect 597738 273776 597744 273788
rect 597796 273776 597802 273828
rect 590654 273680 590660 273692
rect 556540 273652 562364 273680
rect 562428 273652 590660 273680
rect 134426 273504 134432 273556
rect 134484 273544 134490 273556
rect 185118 273544 185124 273556
rect 134484 273516 185124 273544
rect 134484 273504 134490 273516
rect 185118 273504 185124 273516
rect 185176 273504 185182 273556
rect 446398 273504 446404 273556
rect 446456 273544 446462 273556
rect 475930 273544 475936 273556
rect 446456 273516 475936 273544
rect 446456 273504 446462 273516
rect 475930 273504 475936 273516
rect 475988 273504 475994 273556
rect 484302 273504 484308 273556
rect 484360 273544 484366 273556
rect 484360 273516 545804 273544
rect 484360 273504 484366 273516
rect 545776 273476 545804 273516
rect 549898 273504 549904 273556
rect 549956 273544 549962 273556
rect 556540 273544 556568 273652
rect 549956 273516 556568 273544
rect 549956 273504 549962 273516
rect 556798 273504 556804 273556
rect 556856 273544 556862 273556
rect 562428 273544 562456 273652
rect 590654 273640 590660 273652
rect 590712 273640 590718 273692
rect 556856 273516 562456 273544
rect 556856 273504 556862 273516
rect 563698 273504 563704 273556
rect 563756 273544 563762 273556
rect 571978 273544 571984 273556
rect 563756 273516 571984 273544
rect 563756 273504 563762 273516
rect 571978 273504 571984 273516
rect 572036 273504 572042 273556
rect 545776 273448 546816 273476
rect 135622 273368 135628 273420
rect 135680 273408 135686 273420
rect 146938 273408 146944 273420
rect 135680 273380 146944 273408
rect 135680 273368 135686 273380
rect 146938 273368 146944 273380
rect 146996 273368 147002 273420
rect 460014 273368 460020 273420
rect 460072 273408 460078 273420
rect 465718 273408 465724 273420
rect 460072 273380 465724 273408
rect 460072 273368 460078 273380
rect 465718 273368 465724 273380
rect 465776 273368 465782 273420
rect 467558 273368 467564 273420
rect 467616 273408 467622 273420
rect 476114 273408 476120 273420
rect 467616 273380 476120 273408
rect 467616 273368 467622 273380
rect 476114 273368 476120 273380
rect 476172 273368 476178 273420
rect 478690 273368 478696 273420
rect 478748 273408 478754 273420
rect 543688 273408 543694 273420
rect 478748 273380 543694 273408
rect 478748 273368 478754 273380
rect 543688 273368 543694 273380
rect 543746 273368 543752 273420
rect 546788 273408 546816 273448
rect 559926 273408 559932 273420
rect 546788 273380 559932 273408
rect 559926 273368 559932 273380
rect 559984 273368 559990 273420
rect 560294 273368 560300 273420
rect 560352 273408 560358 273420
rect 563422 273408 563428 273420
rect 560352 273380 563428 273408
rect 560352 273368 560358 273380
rect 563422 273368 563428 273380
rect 563480 273368 563486 273420
rect 374638 273300 374644 273352
rect 374696 273340 374702 273352
rect 377858 273340 377864 273352
rect 374696 273312 377864 273340
rect 374696 273300 374702 273312
rect 377858 273300 377864 273312
rect 377916 273300 377922 273352
rect 453298 273300 453304 273352
rect 453356 273340 453362 273352
rect 453758 273340 453764 273352
rect 453356 273312 453764 273340
rect 453356 273300 453362 273312
rect 453758 273300 453764 273312
rect 453816 273300 453822 273352
rect 318610 273232 318616 273284
rect 318668 273272 318674 273284
rect 324682 273272 324688 273284
rect 318668 273244 324688 273272
rect 318668 273232 318674 273244
rect 324682 273232 324688 273244
rect 324740 273232 324746 273284
rect 327534 273232 327540 273284
rect 327592 273272 327598 273284
rect 329466 273272 329472 273284
rect 327592 273244 329472 273272
rect 327592 273232 327598 273244
rect 329466 273232 329472 273244
rect 329524 273232 329530 273284
rect 114370 273164 114376 273216
rect 114428 273204 114434 273216
rect 171594 273204 171600 273216
rect 114428 273176 171600 273204
rect 114428 273164 114434 273176
rect 171594 273164 171600 273176
rect 171652 273164 171658 273216
rect 184106 273164 184112 273216
rect 184164 273204 184170 273216
rect 218882 273204 218888 273216
rect 184164 273176 218888 273204
rect 184164 273164 184170 273176
rect 218882 273164 218888 273176
rect 218940 273164 218946 273216
rect 366358 273164 366364 273216
rect 366416 273204 366422 273216
rect 383838 273204 383844 273216
rect 366416 273176 383844 273204
rect 366416 273164 366422 273176
rect 383838 273164 383844 273176
rect 383896 273164 383902 273216
rect 401502 273164 401508 273216
rect 401560 273204 401566 273216
rect 442902 273204 442908 273216
rect 401560 273176 442908 273204
rect 401560 273164 401566 273176
rect 442902 273164 442908 273176
rect 442960 273164 442966 273216
rect 451182 273164 451188 273216
rect 451240 273204 451246 273216
rect 513834 273204 513840 273216
rect 451240 273176 513840 273204
rect 451240 273164 451246 273176
rect 513834 273164 513840 273176
rect 513892 273164 513898 273216
rect 514018 273164 514024 273216
rect 514076 273204 514082 273216
rect 519722 273204 519728 273216
rect 514076 273176 519728 273204
rect 514076 273164 514082 273176
rect 519722 273164 519728 273176
rect 519780 273164 519786 273216
rect 521470 273164 521476 273216
rect 521528 273204 521534 273216
rect 614298 273204 614304 273216
rect 521528 273176 614304 273204
rect 521528 273164 521534 273176
rect 614298 273164 614304 273176
rect 614356 273164 614362 273216
rect 278590 273096 278596 273148
rect 278648 273136 278654 273148
rect 285858 273136 285864 273148
rect 278648 273108 285864 273136
rect 278648 273096 278654 273108
rect 285858 273096 285864 273108
rect 285916 273096 285922 273148
rect 101306 273028 101312 273080
rect 101364 273068 101370 273080
rect 160922 273068 160928 273080
rect 101364 273040 160928 273068
rect 101364 273028 101370 273040
rect 160922 273028 160928 273040
rect 160980 273028 160986 273080
rect 172238 273028 172244 273080
rect 172296 273068 172302 273080
rect 210602 273068 210608 273080
rect 172296 273040 210608 273068
rect 172296 273028 172302 273040
rect 210602 273028 210608 273040
rect 210660 273028 210666 273080
rect 224034 273028 224040 273080
rect 224092 273068 224098 273080
rect 243262 273068 243268 273080
rect 224092 273040 243268 273068
rect 224092 273028 224098 273040
rect 243262 273028 243268 273040
rect 243320 273028 243326 273080
rect 329466 273028 329472 273080
rect 329524 273068 329530 273080
rect 338850 273068 338856 273080
rect 329524 273040 338856 273068
rect 329524 273028 329530 273040
rect 338850 273028 338856 273040
rect 338908 273028 338914 273080
rect 349798 273028 349804 273080
rect 349856 273068 349862 273080
rect 366082 273068 366088 273080
rect 349856 273040 366088 273068
rect 349856 273028 349862 273040
rect 366082 273028 366088 273040
rect 366140 273028 366146 273080
rect 377398 273028 377404 273080
rect 377456 273068 377462 273080
rect 399202 273068 399208 273080
rect 377456 273040 399208 273068
rect 377456 273028 377462 273040
rect 399202 273028 399208 273040
rect 399260 273028 399266 273080
rect 408218 273028 408224 273080
rect 408276 273068 408282 273080
rect 450814 273068 450820 273080
rect 408276 273040 450820 273068
rect 408276 273028 408282 273040
rect 450814 273028 450820 273040
rect 450872 273028 450878 273080
rect 452286 273028 452292 273080
rect 452344 273068 452350 273080
rect 452344 273040 457392 273068
rect 452344 273028 452350 273040
rect 99006 272892 99012 272944
rect 99064 272932 99070 272944
rect 160094 272932 160100 272944
rect 99064 272904 160100 272932
rect 99064 272892 99070 272904
rect 160094 272892 160100 272904
rect 160152 272892 160158 272944
rect 162762 272892 162768 272944
rect 162820 272932 162826 272944
rect 204714 272932 204720 272944
rect 162820 272904 204720 272932
rect 162820 272892 162826 272904
rect 204714 272892 204720 272904
rect 204772 272892 204778 272944
rect 219526 272892 219532 272944
rect 219584 272932 219590 272944
rect 244458 272932 244464 272944
rect 219584 272904 244464 272932
rect 219584 272892 219590 272904
rect 244458 272892 244464 272904
rect 244516 272892 244522 272944
rect 252646 272892 252652 272944
rect 252704 272932 252710 272944
rect 267918 272932 267924 272944
rect 252704 272904 267924 272932
rect 252704 272892 252710 272904
rect 267918 272892 267924 272904
rect 267976 272892 267982 272944
rect 335262 272892 335268 272944
rect 335320 272932 335326 272944
rect 346854 272932 346860 272944
rect 335320 272904 346860 272932
rect 335320 272892 335326 272904
rect 346854 272892 346860 272904
rect 346912 272892 346918 272944
rect 362770 272892 362776 272944
rect 362828 272932 362834 272944
rect 385862 272932 385868 272944
rect 362828 272904 385868 272932
rect 362828 272892 362834 272904
rect 385862 272892 385868 272904
rect 385920 272892 385926 272944
rect 406838 272892 406844 272944
rect 406896 272932 406902 272944
rect 449986 272932 449992 272944
rect 406896 272904 449992 272932
rect 406896 272892 406902 272904
rect 449986 272892 449992 272904
rect 450044 272892 450050 272944
rect 455230 272892 455236 272944
rect 455288 272932 455294 272944
rect 457364 272932 457392 273040
rect 458082 273028 458088 273080
rect 458140 273068 458146 273080
rect 465534 273068 465540 273080
rect 458140 273040 465540 273068
rect 458140 273028 458146 273040
rect 465534 273028 465540 273040
rect 465592 273028 465598 273080
rect 465718 273028 465724 273080
rect 465776 273068 465782 273080
rect 518526 273068 518532 273080
rect 465776 273040 518532 273068
rect 465776 273028 465782 273040
rect 518526 273028 518532 273040
rect 518584 273028 518590 273080
rect 526806 273028 526812 273080
rect 526864 273068 526870 273080
rect 621382 273068 621388 273080
rect 526864 273040 621388 273068
rect 526864 273028 526870 273040
rect 621382 273028 621388 273040
rect 621440 273028 621446 273080
rect 515030 272932 515036 272944
rect 455288 272904 457300 272932
rect 457364 272904 515036 272932
rect 455288 272892 455294 272904
rect 82446 272756 82452 272808
rect 82504 272796 82510 272808
rect 148410 272796 148416 272808
rect 82504 272768 148416 272796
rect 82504 272756 82510 272768
rect 148410 272756 148416 272768
rect 148468 272756 148474 272808
rect 158070 272756 158076 272808
rect 158128 272796 158134 272808
rect 200666 272796 200672 272808
rect 158128 272768 200672 272796
rect 158128 272756 158134 272768
rect 200666 272756 200672 272768
rect 200724 272756 200730 272808
rect 208854 272756 208860 272808
rect 208912 272796 208918 272808
rect 237374 272796 237380 272808
rect 208912 272768 237380 272796
rect 208912 272756 208918 272768
rect 237374 272756 237380 272768
rect 237432 272756 237438 272808
rect 251450 272756 251456 272808
rect 251508 272796 251514 272808
rect 266998 272796 267004 272808
rect 251508 272768 267004 272796
rect 251508 272756 251514 272768
rect 266998 272756 267004 272768
rect 267056 272756 267062 272808
rect 271506 272756 271512 272808
rect 271564 272796 271570 272808
rect 280338 272796 280344 272808
rect 271564 272768 280344 272796
rect 271564 272756 271570 272768
rect 280338 272756 280344 272768
rect 280396 272756 280402 272808
rect 336366 272756 336372 272808
rect 336424 272796 336430 272808
rect 349522 272796 349528 272808
rect 336424 272768 349528 272796
rect 336424 272756 336430 272768
rect 349522 272756 349528 272768
rect 349580 272756 349586 272808
rect 352558 272756 352564 272808
rect 352616 272796 352622 272808
rect 370774 272796 370780 272808
rect 352616 272768 370780 272796
rect 352616 272756 352622 272768
rect 370774 272756 370780 272768
rect 370832 272756 370838 272808
rect 375190 272756 375196 272808
rect 375248 272796 375254 272808
rect 403894 272796 403900 272808
rect 375248 272768 403900 272796
rect 375248 272756 375254 272768
rect 403894 272756 403900 272768
rect 403952 272756 403958 272808
rect 412266 272756 412272 272808
rect 412324 272796 412330 272808
rect 457070 272796 457076 272808
rect 412324 272768 457076 272796
rect 412324 272756 412330 272768
rect 457070 272756 457076 272768
rect 457128 272756 457134 272808
rect 457272 272796 457300 272904
rect 515030 272892 515036 272904
rect 515088 272892 515094 272944
rect 529842 272892 529848 272944
rect 529900 272932 529906 272944
rect 624970 272932 624976 272944
rect 529900 272904 624976 272932
rect 529900 272892 529906 272904
rect 624970 272892 624976 272904
rect 625028 272892 625034 272944
rect 465718 272796 465724 272808
rect 457272 272768 465724 272796
rect 465718 272756 465724 272768
rect 465776 272756 465782 272808
rect 522114 272796 522120 272808
rect 465920 272768 522120 272796
rect 69382 272620 69388 272672
rect 69440 272660 69446 272672
rect 139394 272660 139400 272672
rect 69440 272632 139400 272660
rect 69440 272620 69446 272632
rect 139394 272620 139400 272632
rect 139452 272620 139458 272672
rect 141510 272620 141516 272672
rect 141568 272660 141574 272672
rect 184934 272660 184940 272672
rect 141568 272632 184940 272660
rect 141568 272620 141574 272632
rect 184934 272620 184940 272632
rect 184992 272620 184998 272672
rect 189074 272620 189080 272672
rect 189132 272660 189138 272672
rect 194042 272660 194048 272672
rect 189132 272632 194048 272660
rect 189132 272620 189138 272632
rect 194042 272620 194048 272632
rect 194100 272620 194106 272672
rect 194686 272620 194692 272672
rect 194744 272660 194750 272672
rect 227162 272660 227168 272672
rect 194744 272632 227168 272660
rect 194744 272620 194750 272632
rect 227162 272620 227168 272632
rect 227220 272620 227226 272672
rect 238478 272620 238484 272672
rect 238536 272660 238542 272672
rect 258074 272660 258080 272672
rect 238536 272632 258080 272660
rect 238536 272620 238542 272632
rect 258074 272620 258080 272632
rect 258132 272620 258138 272672
rect 266814 272620 266820 272672
rect 266872 272660 266878 272672
rect 277578 272660 277584 272672
rect 266872 272632 277584 272660
rect 266872 272620 266878 272632
rect 277578 272620 277584 272632
rect 277636 272620 277642 272672
rect 280982 272620 280988 272672
rect 281040 272660 281046 272672
rect 286318 272660 286324 272672
rect 281040 272632 286324 272660
rect 281040 272620 281046 272632
rect 286318 272620 286324 272632
rect 286376 272620 286382 272672
rect 322750 272620 322756 272672
rect 322808 272660 322814 272672
rect 330570 272660 330576 272672
rect 322808 272632 330576 272660
rect 322808 272620 322814 272632
rect 330570 272620 330576 272632
rect 330628 272620 330634 272672
rect 338022 272620 338028 272672
rect 338080 272660 338086 272672
rect 351914 272660 351920 272672
rect 338080 272632 351920 272660
rect 338080 272620 338086 272632
rect 351914 272620 351920 272632
rect 351972 272620 351978 272672
rect 354490 272620 354496 272672
rect 354548 272660 354554 272672
rect 375558 272660 375564 272672
rect 354548 272632 375564 272660
rect 354548 272620 354554 272632
rect 375558 272620 375564 272632
rect 375616 272620 375622 272672
rect 381998 272620 382004 272672
rect 382056 272660 382062 272672
rect 414566 272660 414572 272672
rect 382056 272632 414572 272660
rect 382056 272620 382062 272632
rect 414566 272620 414572 272632
rect 414624 272620 414630 272672
rect 419166 272620 419172 272672
rect 419224 272660 419230 272672
rect 465350 272660 465356 272672
rect 419224 272632 465356 272660
rect 419224 272620 419230 272632
rect 465350 272620 465356 272632
rect 465408 272620 465414 272672
rect 465534 272620 465540 272672
rect 465592 272660 465598 272672
rect 465920 272660 465948 272768
rect 522114 272756 522120 272768
rect 522172 272756 522178 272808
rect 522758 272756 522764 272808
rect 522816 272796 522822 272808
rect 524138 272796 524144 272808
rect 522816 272768 524144 272796
rect 522816 272756 522822 272768
rect 524138 272756 524144 272768
rect 524196 272756 524202 272808
rect 532510 272756 532516 272808
rect 532568 272796 532574 272808
rect 628466 272796 628472 272808
rect 532568 272768 628472 272796
rect 532568 272756 532574 272768
rect 628466 272756 628472 272768
rect 628524 272756 628530 272808
rect 465592 272632 465948 272660
rect 465592 272620 465598 272632
rect 466086 272620 466092 272672
rect 466144 272660 466150 272672
rect 467374 272660 467380 272672
rect 466144 272632 467380 272660
rect 466144 272620 466150 272632
rect 467374 272620 467380 272632
rect 467432 272620 467438 272672
rect 467742 272620 467748 272672
rect 467800 272660 467806 272672
rect 470410 272660 470416 272672
rect 467800 272632 470416 272660
rect 467800 272620 467806 272632
rect 470410 272620 470416 272632
rect 470468 272620 470474 272672
rect 470594 272620 470600 272672
rect 470652 272660 470658 272672
rect 536282 272660 536288 272672
rect 470652 272632 536288 272660
rect 470652 272620 470658 272632
rect 536282 272620 536288 272632
rect 536340 272620 536346 272672
rect 536558 272620 536564 272672
rect 536616 272660 536622 272672
rect 635550 272660 635556 272672
rect 536616 272632 635556 272660
rect 536616 272620 536622 272632
rect 635550 272620 635556 272632
rect 635608 272620 635614 272672
rect 72970 272484 72976 272536
rect 73028 272524 73034 272536
rect 142154 272524 142160 272536
rect 73028 272496 142160 272524
rect 73028 272484 73034 272496
rect 142154 272484 142160 272496
rect 142212 272484 142218 272536
rect 152182 272484 152188 272536
rect 152240 272524 152246 272536
rect 197538 272524 197544 272536
rect 152240 272496 197544 272524
rect 152240 272484 152246 272496
rect 197538 272484 197544 272496
rect 197596 272484 197602 272536
rect 199470 272484 199476 272536
rect 199528 272524 199534 272536
rect 230566 272524 230572 272536
rect 199528 272496 230572 272524
rect 199528 272484 199534 272496
rect 230566 272484 230572 272496
rect 230624 272484 230630 272536
rect 233694 272484 233700 272536
rect 233752 272524 233758 272536
rect 253934 272524 253940 272536
rect 233752 272496 253940 272524
rect 233752 272484 233758 272496
rect 253934 272484 253940 272496
rect 253992 272484 253998 272536
rect 264422 272484 264428 272536
rect 264480 272524 264486 272536
rect 276014 272524 276020 272536
rect 264480 272496 276020 272524
rect 264480 272484 264486 272496
rect 276014 272484 276020 272496
rect 276072 272484 276078 272536
rect 325510 272484 325516 272536
rect 325568 272524 325574 272536
rect 334158 272524 334164 272536
rect 325568 272496 334164 272524
rect 325568 272484 325574 272496
rect 334158 272484 334164 272496
rect 334216 272484 334222 272536
rect 344646 272484 344652 272536
rect 344704 272524 344710 272536
rect 361390 272524 361396 272536
rect 344704 272496 361396 272524
rect 344704 272484 344710 272496
rect 361390 272484 361396 272496
rect 361448 272484 361454 272536
rect 363782 272484 363788 272536
rect 363840 272524 363846 272536
rect 388530 272524 388536 272536
rect 363840 272496 388536 272524
rect 363840 272484 363846 272496
rect 388530 272484 388536 272496
rect 388588 272484 388594 272536
rect 397270 272484 397276 272536
rect 397328 272524 397334 272536
rect 435818 272524 435824 272536
rect 397328 272496 435824 272524
rect 397328 272484 397334 272496
rect 435818 272484 435824 272496
rect 435876 272484 435882 272536
rect 438762 272484 438768 272536
rect 438820 272524 438826 272536
rect 489868 272524 489874 272536
rect 438820 272496 489874 272524
rect 438820 272484 438826 272496
rect 489868 272484 489874 272496
rect 489926 272484 489932 272536
rect 490006 272484 490012 272536
rect 490064 272524 490070 272536
rect 529198 272524 529204 272536
rect 490064 272496 529204 272524
rect 490064 272484 490070 272496
rect 529198 272484 529204 272496
rect 529256 272484 529262 272536
rect 533706 272484 533712 272536
rect 533764 272524 533770 272536
rect 632054 272524 632060 272536
rect 533764 272496 632060 272524
rect 533764 272484 533770 272496
rect 632054 272484 632060 272496
rect 632112 272484 632118 272536
rect 120258 272348 120264 272400
rect 120316 272388 120322 272400
rect 175274 272388 175280 272400
rect 120316 272360 175280 272388
rect 120316 272348 120322 272360
rect 175274 272348 175280 272360
rect 175332 272348 175338 272400
rect 184934 272348 184940 272400
rect 184992 272388 184998 272400
rect 189166 272388 189172 272400
rect 184992 272360 189172 272388
rect 184992 272348 184998 272360
rect 189166 272348 189172 272360
rect 189224 272348 189230 272400
rect 193582 272348 193588 272400
rect 193640 272388 193646 272400
rect 224218 272388 224224 272400
rect 193640 272360 224224 272388
rect 193640 272348 193646 272360
rect 224218 272348 224224 272360
rect 224276 272348 224282 272400
rect 388990 272348 388996 272400
rect 389048 272388 389054 272400
rect 425146 272388 425152 272400
rect 389048 272360 425152 272388
rect 389048 272348 389054 272360
rect 425146 272348 425152 272360
rect 425204 272348 425210 272400
rect 449802 272348 449808 272400
rect 449860 272388 449866 272400
rect 511442 272388 511448 272400
rect 449860 272360 511448 272388
rect 449860 272348 449866 272360
rect 511442 272348 511448 272360
rect 511500 272348 511506 272400
rect 512638 272348 512644 272400
rect 512696 272388 512702 272400
rect 514018 272388 514024 272400
rect 512696 272360 514024 272388
rect 512696 272348 512702 272360
rect 514018 272348 514024 272360
rect 514076 272348 514082 272400
rect 517330 272348 517336 272400
rect 517388 272388 517394 272400
rect 607214 272388 607220 272400
rect 517388 272360 607220 272388
rect 517388 272348 517394 272360
rect 607214 272348 607220 272360
rect 607272 272348 607278 272400
rect 119062 272212 119068 272264
rect 119120 272252 119126 272264
rect 172514 272252 172520 272264
rect 119120 272224 172520 272252
rect 119120 272212 119126 272224
rect 172514 272212 172520 272224
rect 172572 272212 172578 272264
rect 174446 272212 174452 272264
rect 174504 272252 174510 272264
rect 189350 272252 189356 272264
rect 174504 272224 189356 272252
rect 174504 272212 174510 272224
rect 189350 272212 189356 272224
rect 189408 272212 189414 272264
rect 446950 272212 446956 272264
rect 447008 272252 447014 272264
rect 508038 272252 508044 272264
rect 447008 272224 508044 272252
rect 447008 272212 447014 272224
rect 508038 272212 508044 272224
rect 508096 272212 508102 272264
rect 520090 272212 520096 272264
rect 520148 272252 520154 272264
rect 610710 272252 610716 272264
rect 520148 272224 610716 272252
rect 520148 272212 520154 272224
rect 610710 272212 610716 272224
rect 610768 272212 610774 272264
rect 130838 272076 130844 272128
rect 130896 272116 130902 272128
rect 182450 272116 182456 272128
rect 130896 272088 182456 272116
rect 130896 272076 130902 272088
rect 182450 272076 182456 272088
rect 182508 272076 182514 272128
rect 426342 272076 426348 272128
rect 426400 272116 426406 272128
rect 470548 272116 470554 272128
rect 426400 272088 470554 272116
rect 426400 272076 426406 272088
rect 470548 272076 470554 272088
rect 470606 272076 470612 272128
rect 470778 272076 470784 272128
rect 470836 272116 470842 272128
rect 489868 272116 489874 272128
rect 470836 272088 489874 272116
rect 470836 272076 470842 272088
rect 489868 272076 489874 272088
rect 489926 272076 489932 272128
rect 490006 272076 490012 272128
rect 490064 272116 490070 272128
rect 558730 272116 558736 272128
rect 490064 272088 558736 272116
rect 490064 272076 490070 272088
rect 558730 272076 558736 272088
rect 558788 272076 558794 272128
rect 191466 271940 191472 271992
rect 191524 271980 191530 271992
rect 191524 271952 192800 271980
rect 191524 271940 191530 271952
rect 108390 271804 108396 271856
rect 108448 271844 108454 271856
rect 165890 271844 165896 271856
rect 108448 271816 165896 271844
rect 108448 271804 108454 271816
rect 165890 271804 165896 271816
rect 165948 271804 165954 271856
rect 188798 271804 188804 271856
rect 188856 271844 188862 271856
rect 192570 271844 192576 271856
rect 188856 271816 192576 271844
rect 188856 271804 188862 271816
rect 192570 271804 192576 271816
rect 192628 271804 192634 271856
rect 192772 271844 192800 271952
rect 447778 271940 447784 271992
rect 447836 271980 447842 271992
rect 506750 271980 506756 271992
rect 447836 271952 506756 271980
rect 447836 271940 447842 271952
rect 506750 271940 506756 271952
rect 506808 271940 506814 271992
rect 507118 271940 507124 271992
rect 507176 271980 507182 271992
rect 569402 271980 569408 271992
rect 507176 271952 569408 271980
rect 507176 271940 507182 271952
rect 569402 271940 569408 271952
rect 569460 271940 569466 271992
rect 268838 271872 268844 271924
rect 268896 271912 268902 271924
rect 270494 271912 270500 271924
rect 268896 271884 270500 271912
rect 268896 271872 268902 271884
rect 270494 271872 270500 271884
rect 270552 271872 270558 271924
rect 225046 271844 225052 271856
rect 192772 271816 225052 271844
rect 225046 271804 225052 271816
rect 225104 271804 225110 271856
rect 225414 271804 225420 271856
rect 225472 271844 225478 271856
rect 228358 271844 228364 271856
rect 225472 271816 228364 271844
rect 225472 271804 225478 271816
rect 228358 271804 228364 271816
rect 228416 271804 228422 271856
rect 355318 271804 355324 271856
rect 355376 271844 355382 271856
rect 356606 271844 356612 271856
rect 355376 271816 356612 271844
rect 355376 271804 355382 271816
rect 356606 271804 356612 271816
rect 356664 271804 356670 271856
rect 376570 271804 376576 271856
rect 376628 271844 376634 271856
rect 407482 271844 407488 271856
rect 376628 271816 407488 271844
rect 376628 271804 376634 271816
rect 407482 271804 407488 271816
rect 407540 271804 407546 271856
rect 407758 271804 407764 271856
rect 407816 271844 407822 271856
rect 437014 271844 437020 271856
rect 407816 271816 437020 271844
rect 407816 271804 407822 271816
rect 437014 271804 437020 271816
rect 437072 271804 437078 271856
rect 437198 271804 437204 271856
rect 437256 271844 437262 271856
rect 493686 271844 493692 271856
rect 437256 271816 493692 271844
rect 437256 271804 437262 271816
rect 493686 271804 493692 271816
rect 493744 271804 493750 271856
rect 496538 271804 496544 271856
rect 496596 271844 496602 271856
rect 578510 271844 578516 271856
rect 496596 271816 578516 271844
rect 496596 271804 496602 271816
rect 578510 271804 578516 271816
rect 578568 271804 578574 271856
rect 578878 271804 578884 271856
rect 578936 271844 578942 271856
rect 611906 271844 611912 271856
rect 578936 271816 611912 271844
rect 578936 271804 578942 271816
rect 611906 271804 611912 271816
rect 611964 271804 611970 271856
rect 106090 271668 106096 271720
rect 106148 271708 106154 271720
rect 164970 271708 164976 271720
rect 106148 271680 164976 271708
rect 106148 271668 106154 271680
rect 164970 271668 164976 271680
rect 165028 271668 165034 271720
rect 175734 271668 175740 271720
rect 175792 271708 175798 271720
rect 212994 271708 213000 271720
rect 175792 271680 213000 271708
rect 175792 271668 175798 271680
rect 212994 271668 213000 271680
rect 213052 271668 213058 271720
rect 239858 271668 239864 271720
rect 239916 271708 239922 271720
rect 254118 271708 254124 271720
rect 239916 271680 254124 271708
rect 239916 271668 239922 271680
rect 254118 271668 254124 271680
rect 254176 271668 254182 271720
rect 353938 271668 353944 271720
rect 353996 271708 354002 271720
rect 372798 271708 372804 271720
rect 353996 271680 372804 271708
rect 353996 271668 354002 271680
rect 372798 271668 372804 271680
rect 372856 271668 372862 271720
rect 384942 271668 384948 271720
rect 385000 271708 385006 271720
rect 418062 271708 418068 271720
rect 385000 271680 418068 271708
rect 385000 271668 385006 271680
rect 418062 271668 418068 271680
rect 418120 271668 418126 271720
rect 420178 271668 420184 271720
rect 420236 271708 420242 271720
rect 431126 271708 431132 271720
rect 420236 271680 431132 271708
rect 420236 271668 420242 271680
rect 431126 271668 431132 271680
rect 431184 271668 431190 271720
rect 434622 271668 434628 271720
rect 434680 271708 434686 271720
rect 485222 271708 485228 271720
rect 434680 271680 485228 271708
rect 434680 271668 434686 271680
rect 485222 271668 485228 271680
rect 485280 271668 485286 271720
rect 485406 271668 485412 271720
rect 485464 271708 485470 271720
rect 490006 271708 490012 271720
rect 485464 271680 490012 271708
rect 485464 271668 485470 271680
rect 490006 271668 490012 271680
rect 490064 271668 490070 271720
rect 501966 271668 501972 271720
rect 502024 271708 502030 271720
rect 585962 271708 585968 271720
rect 502024 271680 585968 271708
rect 502024 271668 502030 271680
rect 585962 271668 585968 271680
rect 586020 271668 586026 271720
rect 94222 271532 94228 271584
rect 94280 271572 94286 271584
rect 156138 271572 156144 271584
rect 94280 271544 156144 271572
rect 94280 271532 94286 271544
rect 156138 271532 156144 271544
rect 156196 271532 156202 271584
rect 170122 271532 170128 271584
rect 170180 271572 170186 271584
rect 209774 271572 209780 271584
rect 170180 271544 209780 271572
rect 170180 271532 170186 271544
rect 209774 271532 209780 271544
rect 209832 271532 209838 271584
rect 223114 271532 223120 271584
rect 223172 271572 223178 271584
rect 247218 271572 247224 271584
rect 223172 271544 247224 271572
rect 223172 271532 223178 271544
rect 247218 271532 247224 271544
rect 247276 271532 247282 271584
rect 357158 271532 357164 271584
rect 357216 271572 357222 271584
rect 379054 271572 379060 271584
rect 357216 271544 379060 271572
rect 357216 271532 357222 271544
rect 379054 271532 379060 271544
rect 379112 271532 379118 271584
rect 387610 271532 387616 271584
rect 387668 271572 387674 271584
rect 422846 271572 422852 271584
rect 387668 271544 422852 271572
rect 387668 271532 387674 271544
rect 422846 271532 422852 271544
rect 422904 271532 422910 271584
rect 439958 271532 439964 271584
rect 440016 271572 440022 271584
rect 497274 271572 497280 271584
rect 440016 271544 497280 271572
rect 440016 271532 440022 271544
rect 497274 271532 497280 271544
rect 497332 271532 497338 271584
rect 499298 271532 499304 271584
rect 499356 271572 499362 271584
rect 582374 271572 582380 271584
rect 499356 271544 582380 271572
rect 499356 271532 499362 271544
rect 582374 271532 582380 271544
rect 582432 271532 582438 271584
rect 585778 271532 585784 271584
rect 585836 271572 585842 271584
rect 626074 271572 626080 271584
rect 585836 271544 626080 271572
rect 585836 271532 585842 271544
rect 626074 271532 626080 271544
rect 626132 271532 626138 271584
rect 87138 271396 87144 271448
rect 87196 271436 87202 271448
rect 152182 271436 152188 271448
rect 87196 271408 152188 271436
rect 87196 271396 87202 271408
rect 152182 271396 152188 271408
rect 152240 271396 152246 271448
rect 159266 271396 159272 271448
rect 159324 271436 159330 271448
rect 202322 271436 202328 271448
rect 159324 271408 202328 271436
rect 159324 271396 159330 271408
rect 202322 271396 202328 271408
rect 202380 271396 202386 271448
rect 213638 271396 213644 271448
rect 213696 271436 213702 271448
rect 240410 271436 240416 271448
rect 213696 271408 240416 271436
rect 213696 271396 213702 271408
rect 240410 271396 240416 271408
rect 240468 271396 240474 271448
rect 250254 271396 250260 271448
rect 250312 271436 250318 271448
rect 250312 271408 262444 271436
rect 250312 271396 250318 271408
rect 75362 271260 75368 271312
rect 75420 271300 75426 271312
rect 75420 271272 142154 271300
rect 75420 271260 75426 271272
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 142126 271164 142154 271272
rect 142706 271260 142712 271312
rect 142764 271300 142770 271312
rect 144178 271300 144184 271312
rect 142764 271272 144184 271300
rect 142764 271260 142770 271272
rect 144178 271260 144184 271272
rect 144236 271260 144242 271312
rect 154298 271260 154304 271312
rect 154356 271300 154362 271312
rect 198090 271300 198096 271312
rect 154356 271272 198096 271300
rect 154356 271260 154362 271272
rect 198090 271260 198096 271272
rect 198148 271260 198154 271312
rect 212258 271260 212264 271312
rect 212316 271300 212322 271312
rect 239306 271300 239312 271312
rect 212316 271272 239312 271300
rect 212316 271260 212322 271272
rect 239306 271260 239312 271272
rect 239364 271260 239370 271312
rect 244642 271260 244648 271312
rect 244700 271300 244706 271312
rect 262214 271300 262220 271312
rect 244700 271272 262220 271300
rect 244700 271260 244706 271272
rect 262214 271260 262220 271272
rect 262272 271260 262278 271312
rect 262416 271300 262444 271408
rect 265618 271396 265624 271448
rect 265676 271436 265682 271448
rect 276842 271436 276848 271448
rect 265676 271408 276848 271436
rect 265676 271396 265682 271408
rect 276842 271396 276848 271408
rect 276900 271396 276906 271448
rect 339218 271396 339224 271448
rect 339276 271436 339282 271448
rect 354214 271436 354220 271448
rect 339276 271408 354220 271436
rect 339276 271396 339282 271408
rect 354214 271396 354220 271408
rect 354272 271396 354278 271448
rect 358722 271396 358728 271448
rect 358780 271436 358786 271448
rect 381446 271436 381452 271448
rect 358780 271408 381452 271436
rect 358780 271396 358786 271408
rect 381446 271396 381452 271408
rect 381504 271396 381510 271448
rect 393958 271396 393964 271448
rect 394016 271436 394022 271448
rect 429930 271436 429936 271448
rect 394016 271408 429936 271436
rect 394016 271396 394022 271408
rect 429930 271396 429936 271408
rect 429988 271396 429994 271448
rect 442902 271396 442908 271448
rect 442960 271436 442966 271448
rect 500862 271436 500868 271448
rect 442960 271408 500868 271436
rect 442960 271396 442966 271408
rect 500862 271396 500868 271408
rect 500920 271396 500926 271448
rect 505002 271396 505008 271448
rect 505060 271436 505066 271448
rect 589458 271436 589464 271448
rect 505060 271408 589464 271436
rect 505060 271396 505066 271408
rect 589458 271396 589464 271408
rect 589516 271396 589522 271448
rect 266446 271300 266452 271312
rect 262416 271272 266452 271300
rect 266446 271260 266452 271272
rect 266504 271260 266510 271312
rect 276658 271260 276664 271312
rect 276716 271300 276722 271312
rect 284478 271300 284484 271312
rect 276716 271272 284484 271300
rect 276716 271260 276722 271272
rect 284478 271260 284484 271272
rect 284536 271260 284542 271312
rect 329650 271260 329656 271312
rect 329708 271300 329714 271312
rect 340046 271300 340052 271312
rect 329708 271272 340052 271300
rect 329708 271260 329714 271272
rect 340046 271260 340052 271272
rect 340104 271260 340110 271312
rect 340598 271260 340604 271312
rect 340656 271300 340662 271312
rect 355134 271300 355140 271312
rect 340656 271272 355140 271300
rect 340656 271260 340662 271272
rect 355134 271260 355140 271272
rect 355192 271260 355198 271312
rect 365438 271260 365444 271312
rect 365496 271300 365502 271312
rect 390922 271300 390928 271312
rect 365496 271272 390928 271300
rect 365496 271260 365502 271272
rect 390922 271260 390928 271272
rect 390980 271260 390986 271312
rect 391842 271260 391848 271312
rect 391900 271300 391906 271312
rect 428734 271300 428740 271312
rect 391900 271272 428740 271300
rect 391900 271260 391906 271272
rect 428734 271260 428740 271272
rect 428792 271260 428798 271312
rect 445662 271260 445668 271312
rect 445720 271300 445726 271312
rect 504358 271300 504364 271312
rect 445720 271272 504364 271300
rect 445720 271260 445726 271272
rect 504358 271260 504364 271272
rect 504416 271260 504422 271312
rect 507670 271260 507676 271312
rect 507728 271300 507734 271312
rect 593046 271300 593052 271312
rect 507728 271272 593052 271300
rect 507728 271260 507734 271272
rect 593046 271260 593052 271272
rect 593104 271260 593110 271312
rect 611998 271260 612004 271312
rect 612056 271300 612062 271312
rect 618622 271300 618628 271312
rect 612056 271272 618628 271300
rect 612056 271260 612062 271272
rect 618622 271260 618628 271272
rect 618680 271260 618686 271312
rect 618898 271260 618904 271312
rect 618956 271300 618962 271312
rect 633250 271300 633256 271312
rect 618956 271272 633256 271300
rect 618956 271260 618962 271272
rect 633250 271260 633256 271272
rect 633308 271260 633314 271312
rect 142706 271164 142712 271176
rect 142126 271136 142712 271164
rect 142706 271124 142712 271136
rect 142764 271124 142770 271176
rect 148594 271124 148600 271176
rect 148652 271164 148658 271176
rect 194778 271164 194784 271176
rect 148652 271136 194784 271164
rect 148652 271124 148658 271136
rect 194778 271124 194784 271136
rect 194836 271124 194842 271176
rect 197078 271124 197084 271176
rect 197136 271164 197142 271176
rect 229278 271164 229284 271176
rect 197136 271136 229284 271164
rect 197136 271124 197142 271136
rect 229278 271124 229284 271136
rect 229336 271124 229342 271176
rect 230198 271124 230204 271176
rect 230256 271164 230262 271176
rect 251726 271164 251732 271176
rect 230256 271136 251732 271164
rect 230256 271124 230262 271136
rect 251726 271124 251732 271136
rect 251784 271124 251790 271176
rect 254946 271124 254952 271176
rect 255004 271164 255010 271176
rect 269298 271164 269304 271176
rect 255004 271136 269304 271164
rect 255004 271124 255010 271136
rect 269298 271124 269304 271136
rect 269356 271124 269362 271176
rect 270310 271124 270316 271176
rect 270368 271164 270374 271176
rect 280522 271164 280528 271176
rect 270368 271136 280528 271164
rect 270368 271124 270374 271136
rect 280522 271124 280528 271136
rect 280580 271124 280586 271176
rect 331122 271124 331128 271176
rect 331180 271164 331186 271176
rect 342438 271164 342444 271176
rect 331180 271136 342444 271164
rect 331180 271124 331186 271136
rect 342438 271124 342444 271136
rect 342496 271124 342502 271176
rect 347590 271124 347596 271176
rect 347648 271164 347654 271176
rect 364518 271164 364524 271176
rect 347648 271136 364524 271164
rect 347648 271124 347654 271136
rect 364518 271124 364524 271136
rect 364576 271124 364582 271176
rect 366910 271124 366916 271176
rect 366968 271164 366974 271176
rect 393314 271164 393320 271176
rect 366968 271136 393320 271164
rect 366968 271124 366974 271136
rect 393314 271124 393320 271136
rect 393372 271124 393378 271176
rect 402606 271124 402612 271176
rect 402664 271164 402670 271176
rect 444098 271164 444104 271176
rect 402664 271136 444104 271164
rect 402664 271124 402670 271136
rect 444098 271124 444104 271136
rect 444156 271124 444162 271176
rect 459462 271124 459468 271176
rect 459520 271164 459526 271176
rect 523862 271164 523868 271176
rect 459520 271136 523868 271164
rect 459520 271124 459526 271136
rect 523862 271124 523868 271136
rect 523920 271124 523926 271176
rect 524046 271124 524052 271176
rect 524104 271164 524110 271176
rect 617794 271164 617800 271176
rect 524104 271136 617800 271164
rect 524104 271124 524110 271136
rect 617794 271124 617800 271136
rect 617852 271124 617858 271176
rect 625798 271124 625804 271176
rect 625856 271164 625862 271176
rect 645026 271164 645032 271176
rect 625856 271136 645032 271164
rect 625856 271124 625862 271136
rect 645026 271124 645032 271136
rect 645084 271124 645090 271176
rect 116670 270988 116676 271040
rect 116728 271028 116734 271040
rect 172698 271028 172704 271040
rect 116728 271000 172704 271028
rect 116728 270988 116734 271000
rect 172698 270988 172704 271000
rect 172756 270988 172762 271040
rect 192754 270988 192760 271040
rect 192812 271028 192818 271040
rect 225506 271028 225512 271040
rect 192812 271000 225512 271028
rect 192812 270988 192818 271000
rect 225506 270988 225512 271000
rect 225564 270988 225570 271040
rect 326430 270988 326436 271040
rect 326488 271028 326494 271040
rect 335078 271028 335084 271040
rect 326488 271000 335084 271028
rect 326488 270988 326494 271000
rect 335078 270988 335084 271000
rect 335136 270988 335142 271040
rect 381538 270988 381544 271040
rect 381596 271028 381602 271040
rect 411806 271028 411812 271040
rect 381596 271000 411812 271028
rect 381596 270988 381602 271000
rect 411806 270988 411812 271000
rect 411864 270988 411870 271040
rect 414474 270988 414480 271040
rect 414532 271028 414538 271040
rect 438118 271028 438124 271040
rect 414532 271000 438124 271028
rect 414532 270988 414538 271000
rect 438118 270988 438124 271000
rect 438176 270988 438182 271040
rect 438302 270988 438308 271040
rect 438360 271028 438366 271040
rect 438360 271000 485084 271028
rect 438360 270988 438366 271000
rect 124950 270852 124956 270904
rect 125008 270892 125014 270904
rect 178678 270892 178684 270904
rect 125008 270864 178684 270892
rect 125008 270852 125014 270864
rect 178678 270852 178684 270864
rect 178736 270852 178742 270904
rect 417418 270852 417424 270904
rect 417476 270892 417482 270904
rect 427538 270892 427544 270904
rect 417476 270864 427544 270892
rect 417476 270852 417482 270864
rect 427538 270852 427544 270864
rect 427596 270852 427602 270904
rect 430390 270852 430396 270904
rect 430448 270892 430454 270904
rect 483106 270892 483112 270904
rect 430448 270864 483112 270892
rect 430448 270852 430454 270864
rect 483106 270852 483112 270864
rect 483164 270852 483170 270904
rect 485056 270892 485084 271000
rect 485222 270988 485228 271040
rect 485280 271028 485286 271040
rect 490190 271028 490196 271040
rect 485280 271000 490196 271028
rect 485280 270988 485286 271000
rect 490190 270988 490196 271000
rect 490248 270988 490254 271040
rect 495250 270988 495256 271040
rect 495308 271028 495314 271040
rect 575290 271028 575296 271040
rect 495308 271000 575296 271028
rect 495308 270988 495314 271000
rect 575290 270988 575296 271000
rect 575348 270988 575354 271040
rect 492398 270892 492404 270904
rect 485056 270864 492404 270892
rect 492398 270852 492404 270864
rect 492456 270852 492462 270904
rect 492582 270852 492588 270904
rect 492640 270892 492646 270904
rect 571610 270892 571616 270904
rect 492640 270864 571616 270892
rect 492640 270852 492646 270864
rect 571610 270852 571616 270864
rect 571668 270852 571674 270904
rect 571978 270852 571984 270904
rect 572036 270892 572042 270904
rect 604822 270892 604828 270904
rect 572036 270864 604828 270892
rect 572036 270852 572042 270864
rect 604822 270852 604828 270864
rect 604880 270852 604886 270904
rect 127342 270716 127348 270768
rect 127400 270756 127406 270768
rect 179874 270756 179880 270768
rect 127400 270728 179880 270756
rect 127400 270716 127406 270728
rect 179874 270716 179880 270728
rect 179932 270716 179938 270768
rect 321370 270716 321376 270768
rect 321428 270756 321434 270768
rect 327074 270756 327080 270768
rect 321428 270728 327080 270756
rect 321428 270716 321434 270728
rect 327074 270716 327080 270728
rect 327132 270716 327138 270768
rect 427446 270716 427452 270768
rect 427504 270756 427510 270768
rect 479150 270756 479156 270768
rect 427504 270728 479156 270756
rect 427504 270716 427510 270728
rect 479150 270716 479156 270728
rect 479208 270716 479214 270768
rect 486878 270716 486884 270768
rect 486936 270756 486942 270768
rect 564618 270756 564624 270768
rect 486936 270728 564624 270756
rect 486936 270716 486942 270728
rect 564618 270716 564624 270728
rect 564676 270716 564682 270768
rect 137922 270580 137928 270632
rect 137980 270620 137986 270632
rect 187694 270620 187700 270632
rect 137980 270592 187700 270620
rect 137980 270580 137986 270592
rect 187694 270580 187700 270592
rect 187752 270580 187758 270632
rect 422938 270580 422944 270632
rect 422996 270620 423002 270632
rect 445294 270620 445300 270632
rect 422996 270592 445300 270620
rect 422996 270580 423002 270592
rect 445294 270580 445300 270592
rect 445352 270580 445358 270632
rect 489638 270580 489644 270632
rect 489696 270620 489702 270632
rect 568206 270620 568212 270632
rect 489696 270592 568212 270620
rect 489696 270580 489702 270592
rect 568206 270580 568212 270592
rect 568264 270580 568270 270632
rect 129458 270444 129464 270496
rect 129516 270484 129522 270496
rect 181162 270484 181168 270496
rect 129516 270456 181168 270484
rect 129516 270444 129522 270456
rect 181162 270444 181168 270456
rect 181220 270444 181226 270496
rect 191742 270444 191748 270496
rect 191800 270484 191806 270496
rect 196894 270484 196900 270496
rect 191800 270456 196900 270484
rect 191800 270444 191806 270456
rect 196894 270444 196900 270456
rect 196952 270444 196958 270496
rect 201770 270444 201776 270496
rect 201828 270484 201834 270496
rect 232222 270484 232228 270496
rect 201828 270456 232228 270484
rect 201828 270444 201834 270456
rect 232222 270444 232228 270456
rect 232280 270444 232286 270496
rect 395614 270444 395620 270496
rect 395672 270484 395678 270496
rect 433610 270484 433616 270496
rect 395672 270456 433616 270484
rect 395672 270444 395678 270456
rect 433610 270444 433616 270456
rect 433668 270444 433674 270496
rect 453574 270444 453580 270496
rect 453632 270484 453638 270496
rect 516778 270484 516784 270496
rect 453632 270456 516784 270484
rect 453632 270444 453638 270456
rect 516778 270444 516784 270456
rect 516836 270444 516842 270496
rect 517514 270444 517520 270496
rect 517572 270484 517578 270496
rect 579614 270484 579620 270496
rect 517572 270456 579620 270484
rect 517572 270444 517578 270456
rect 579614 270444 579620 270456
rect 579672 270444 579678 270496
rect 581638 270444 581644 270496
rect 581696 270484 581702 270496
rect 620278 270484 620284 270496
rect 581696 270456 620284 270484
rect 581696 270444 581702 270456
rect 620278 270444 620284 270456
rect 620336 270444 620342 270496
rect 88334 270308 88340 270360
rect 88392 270348 88398 270360
rect 121454 270348 121460 270360
rect 88392 270320 121460 270348
rect 88392 270308 88398 270320
rect 121454 270308 121460 270320
rect 121512 270308 121518 270360
rect 122558 270308 122564 270360
rect 122616 270348 122622 270360
rect 176194 270348 176200 270360
rect 122616 270320 176200 270348
rect 122616 270308 122622 270320
rect 176194 270308 176200 270320
rect 176252 270308 176258 270360
rect 180702 270308 180708 270360
rect 180760 270348 180766 270360
rect 215294 270348 215300 270360
rect 180760 270320 215300 270348
rect 180760 270308 180766 270320
rect 215294 270308 215300 270320
rect 215352 270308 215358 270360
rect 232774 270308 232780 270360
rect 232832 270348 232838 270360
rect 247862 270348 247868 270360
rect 232832 270320 247868 270348
rect 232832 270308 232838 270320
rect 247862 270308 247868 270320
rect 247920 270308 247926 270360
rect 262858 270308 262864 270360
rect 262916 270348 262922 270360
rect 262916 270320 267734 270348
rect 262916 270308 262922 270320
rect 97902 270172 97908 270224
rect 97960 270212 97966 270224
rect 158806 270212 158812 270224
rect 97960 270184 158812 270212
rect 97960 270172 97966 270184
rect 158806 270172 158812 270184
rect 158864 270172 158870 270224
rect 179322 270172 179328 270224
rect 179380 270212 179386 270224
rect 214098 270212 214104 270224
rect 179380 270184 214104 270212
rect 179380 270172 179386 270184
rect 214098 270172 214104 270184
rect 214156 270172 214162 270224
rect 226610 270172 226616 270224
rect 226668 270212 226674 270224
rect 249886 270212 249892 270224
rect 226668 270184 249892 270212
rect 226668 270172 226674 270184
rect 249886 270172 249892 270184
rect 249944 270172 249950 270224
rect 259730 270172 259736 270224
rect 259788 270212 259794 270224
rect 267706 270212 267734 270320
rect 367462 270308 367468 270360
rect 367520 270348 367526 270360
rect 393498 270348 393504 270360
rect 367520 270320 393504 270348
rect 367520 270308 367526 270320
rect 393498 270308 393504 270320
rect 393556 270308 393562 270360
rect 400858 270308 400864 270360
rect 400916 270348 400922 270360
rect 441614 270348 441620 270360
rect 400916 270320 441620 270348
rect 400916 270308 400922 270320
rect 441614 270308 441620 270320
rect 441672 270308 441678 270360
rect 456058 270308 456064 270360
rect 456116 270348 456122 270360
rect 520274 270348 520280 270360
rect 456116 270320 520280 270348
rect 456116 270308 456122 270320
rect 520274 270308 520280 270320
rect 520332 270308 520338 270360
rect 524414 270348 524420 270360
rect 521672 270320 524420 270348
rect 271414 270212 271420 270224
rect 259788 270184 265020 270212
rect 267706 270184 271420 270212
rect 259788 270172 259794 270184
rect 85482 270036 85488 270088
rect 85540 270076 85546 270088
rect 149422 270076 149428 270088
rect 85540 270048 149428 270076
rect 85540 270036 85546 270048
rect 149422 270036 149428 270048
rect 149480 270036 149486 270088
rect 173710 270036 173716 270088
rect 173768 270076 173774 270088
rect 212626 270076 212632 270088
rect 173768 270048 212632 270076
rect 173768 270036 173774 270048
rect 212626 270036 212632 270048
rect 212684 270036 212690 270088
rect 216490 270036 216496 270088
rect 216548 270076 216554 270088
rect 242434 270076 242440 270088
rect 216548 270048 242440 270076
rect 216548 270036 216554 270048
rect 242434 270036 242440 270048
rect 242492 270036 242498 270088
rect 248322 270036 248328 270088
rect 248380 270076 248386 270088
rect 264790 270076 264796 270088
rect 248380 270048 264796 270076
rect 248380 270036 248386 270048
rect 264790 270036 264796 270048
rect 264848 270036 264854 270088
rect 70578 269900 70584 269952
rect 70636 269940 70642 269952
rect 79962 269940 79968 269952
rect 70636 269912 79968 269940
rect 70636 269900 70642 269912
rect 79962 269900 79968 269912
rect 80020 269900 80026 269952
rect 80146 269900 80152 269952
rect 80204 269940 80210 269952
rect 146386 269940 146392 269952
rect 80204 269912 146392 269940
rect 80204 269900 80210 269912
rect 146386 269900 146392 269912
rect 146444 269900 146450 269952
rect 165430 269900 165436 269952
rect 165488 269940 165494 269952
rect 206002 269940 206008 269952
rect 165488 269912 206008 269940
rect 165488 269900 165494 269912
rect 206002 269900 206008 269912
rect 206060 269900 206066 269952
rect 210050 269900 210056 269952
rect 210108 269940 210114 269952
rect 238294 269940 238300 269952
rect 210108 269912 238300 269940
rect 210108 269900 210114 269912
rect 238294 269900 238300 269912
rect 238352 269900 238358 269952
rect 241974 269900 241980 269952
rect 242032 269940 242038 269952
rect 260374 269940 260380 269952
rect 242032 269912 260380 269940
rect 242032 269900 242038 269912
rect 260374 269900 260380 269912
rect 260432 269900 260438 269952
rect 264992 269940 265020 270184
rect 271414 270172 271420 270184
rect 271472 270172 271478 270224
rect 345106 270172 345112 270224
rect 345164 270212 345170 270224
rect 361574 270212 361580 270224
rect 345164 270184 361580 270212
rect 345164 270172 345170 270184
rect 361574 270172 361580 270184
rect 361632 270172 361638 270224
rect 364150 270172 364156 270224
rect 364208 270212 364214 270224
rect 389174 270212 389180 270224
rect 364208 270184 389180 270212
rect 364208 270172 364214 270184
rect 389174 270172 389180 270184
rect 389232 270172 389238 270224
rect 390094 270172 390100 270224
rect 390152 270212 390158 270224
rect 405734 270212 405740 270224
rect 390152 270184 405740 270212
rect 390152 270172 390158 270184
rect 405734 270172 405740 270184
rect 405792 270172 405798 270224
rect 409690 270172 409696 270224
rect 409748 270212 409754 270224
rect 454034 270212 454040 270224
rect 409748 270184 454040 270212
rect 409748 270172 409754 270184
rect 454034 270172 454040 270184
rect 454092 270172 454098 270224
rect 458542 270172 458548 270224
rect 458600 270212 458606 270224
rect 521672 270212 521700 270320
rect 524414 270308 524420 270320
rect 524472 270308 524478 270360
rect 525610 270308 525616 270360
rect 525668 270348 525674 270360
rect 525668 270320 533384 270348
rect 525668 270308 525674 270320
rect 458600 270184 521700 270212
rect 458600 270172 458606 270184
rect 523126 270172 523132 270224
rect 523184 270212 523190 270224
rect 533154 270212 533160 270224
rect 523184 270184 533160 270212
rect 523184 270172 523190 270184
rect 533154 270172 533160 270184
rect 533212 270172 533218 270224
rect 533356 270212 533384 270320
rect 533522 270308 533528 270360
rect 533580 270348 533586 270360
rect 626534 270348 626540 270360
rect 533580 270320 626540 270348
rect 533580 270308 533586 270320
rect 626534 270308 626540 270320
rect 626592 270308 626598 270360
rect 619634 270212 619640 270224
rect 533356 270184 619640 270212
rect 619634 270172 619640 270184
rect 619692 270172 619698 270224
rect 623958 270212 623964 270224
rect 619836 270184 623964 270212
rect 327718 270036 327724 270088
rect 327776 270076 327782 270088
rect 336734 270076 336740 270088
rect 327776 270048 336740 270076
rect 327776 270036 327782 270048
rect 336734 270036 336740 270048
rect 336792 270036 336798 270088
rect 345934 270036 345940 270088
rect 345992 270076 345998 270088
rect 362954 270076 362960 270088
rect 345992 270048 362960 270076
rect 345992 270036 345998 270048
rect 362954 270036 362960 270048
rect 363012 270036 363018 270088
rect 369854 270036 369860 270088
rect 369912 270076 369918 270088
rect 396074 270076 396080 270088
rect 369912 270048 396080 270076
rect 369912 270036 369918 270048
rect 396074 270036 396080 270048
rect 396132 270036 396138 270088
rect 399846 270036 399852 270088
rect 399904 270076 399910 270088
rect 412634 270076 412640 270088
rect 399904 270048 412640 270076
rect 399904 270036 399910 270048
rect 412634 270036 412640 270048
rect 412692 270036 412698 270088
rect 414658 270036 414664 270088
rect 414716 270076 414722 270088
rect 460934 270076 460940 270088
rect 414716 270048 460940 270076
rect 414716 270036 414722 270048
rect 460934 270036 460940 270048
rect 460992 270036 460998 270088
rect 461394 270036 461400 270088
rect 461452 270076 461458 270088
rect 527174 270076 527180 270088
rect 461452 270048 527180 270076
rect 461452 270036 461458 270048
rect 527174 270036 527180 270048
rect 527232 270036 527238 270088
rect 528370 270036 528376 270088
rect 528428 270076 528434 270088
rect 619836 270076 619864 270184
rect 623958 270172 623964 270184
rect 624016 270172 624022 270224
rect 528428 270048 619864 270076
rect 528428 270036 528434 270048
rect 620278 270036 620284 270088
rect 620336 270076 620342 270088
rect 630674 270076 630680 270088
rect 620336 270048 630680 270076
rect 620336 270036 620342 270048
rect 630674 270036 630680 270048
rect 630732 270036 630738 270088
rect 273070 269940 273076 269952
rect 264992 269912 273076 269940
rect 273070 269900 273076 269912
rect 273128 269900 273134 269952
rect 326890 269900 326896 269952
rect 326948 269940 326954 269952
rect 335538 269940 335544 269952
rect 326948 269912 335544 269940
rect 326948 269900 326954 269912
rect 335538 269900 335544 269912
rect 335596 269900 335602 269952
rect 336826 269900 336832 269952
rect 336884 269940 336890 269952
rect 350534 269940 350540 269952
rect 336884 269912 350540 269940
rect 336884 269900 336890 269912
rect 350534 269900 350540 269912
rect 350592 269900 350598 269952
rect 351730 269900 351736 269952
rect 351788 269940 351794 269952
rect 371234 269940 371240 269952
rect 351788 269912 371240 269940
rect 351788 269900 351794 269912
rect 371234 269900 371240 269912
rect 371292 269900 371298 269952
rect 372430 269900 372436 269952
rect 372488 269940 372494 269952
rect 400490 269940 400496 269952
rect 372488 269912 400496 269940
rect 372488 269900 372494 269912
rect 400490 269900 400496 269912
rect 400548 269900 400554 269952
rect 401870 269900 401876 269952
rect 401928 269940 401934 269952
rect 416774 269940 416780 269952
rect 401928 269912 416780 269940
rect 401928 269900 401934 269912
rect 416774 269900 416780 269912
rect 416832 269900 416838 269952
rect 417142 269900 417148 269952
rect 417200 269940 417206 269952
rect 465074 269940 465080 269952
rect 417200 269912 465080 269940
rect 417200 269900 417206 269912
rect 465074 269900 465080 269912
rect 465132 269900 465138 269952
rect 468478 269900 468484 269952
rect 468536 269940 468542 269952
rect 468536 269912 531820 269940
rect 468536 269900 468542 269912
rect 76742 269764 76748 269816
rect 76800 269804 76806 269816
rect 143902 269804 143908 269816
rect 76800 269776 143908 269804
rect 76800 269764 76806 269776
rect 143902 269764 143908 269776
rect 143960 269764 143966 269816
rect 144362 269764 144368 269816
rect 144420 269804 144426 269816
rect 190822 269804 190828 269816
rect 144420 269776 190828 269804
rect 144420 269764 144426 269776
rect 190822 269764 190828 269776
rect 190880 269764 190886 269816
rect 202966 269764 202972 269816
rect 203024 269804 203030 269816
rect 233326 269804 233332 269816
rect 203024 269776 233332 269804
rect 203024 269764 203030 269776
rect 233326 269764 233332 269776
rect 233384 269764 233390 269816
rect 241422 269764 241428 269816
rect 241480 269804 241486 269816
rect 259822 269804 259828 269816
rect 241480 269776 259828 269804
rect 241480 269764 241486 269776
rect 259822 269764 259828 269776
rect 259880 269764 259886 269816
rect 261938 269764 261944 269816
rect 261996 269804 262002 269816
rect 274726 269804 274732 269816
rect 261996 269776 274732 269804
rect 261996 269764 262002 269776
rect 274726 269764 274732 269776
rect 274784 269764 274790 269816
rect 280062 269764 280068 269816
rect 280120 269804 280126 269816
rect 287146 269804 287152 269816
rect 280120 269776 287152 269804
rect 280120 269764 280126 269776
rect 287146 269764 287152 269776
rect 287204 269764 287210 269816
rect 335078 269764 335084 269816
rect 335136 269804 335142 269816
rect 347774 269804 347780 269816
rect 335136 269776 347780 269804
rect 335136 269764 335142 269776
rect 347774 269764 347780 269776
rect 347832 269764 347838 269816
rect 355042 269764 355048 269816
rect 355100 269804 355106 269816
rect 376938 269804 376944 269816
rect 355100 269776 376944 269804
rect 355100 269764 355106 269776
rect 376938 269764 376944 269776
rect 376996 269764 377002 269816
rect 377674 269764 377680 269816
rect 377732 269804 377738 269816
rect 408494 269804 408500 269816
rect 377732 269776 408500 269804
rect 377732 269764 377738 269776
rect 408494 269764 408500 269776
rect 408552 269764 408558 269816
rect 412450 269764 412456 269816
rect 412508 269804 412514 269816
rect 458266 269804 458272 269816
rect 412508 269776 458272 269804
rect 412508 269764 412514 269776
rect 458266 269764 458272 269776
rect 458324 269764 458330 269816
rect 463510 269764 463516 269816
rect 463568 269804 463574 269816
rect 531314 269804 531320 269816
rect 463568 269776 531320 269804
rect 463568 269764 463574 269776
rect 531314 269764 531320 269776
rect 531372 269764 531378 269816
rect 531792 269804 531820 269912
rect 531958 269900 531964 269952
rect 532016 269940 532022 269952
rect 533522 269940 533528 269952
rect 532016 269912 533528 269940
rect 532016 269900 532022 269912
rect 533522 269900 533528 269912
rect 533580 269900 533586 269952
rect 533982 269900 533988 269952
rect 534040 269940 534046 269952
rect 537754 269940 537760 269952
rect 534040 269912 537760 269940
rect 534040 269900 534046 269912
rect 537754 269900 537760 269912
rect 537812 269900 537818 269952
rect 537938 269900 537944 269952
rect 537996 269940 538002 269952
rect 537996 269912 543044 269940
rect 537996 269900 538002 269912
rect 538490 269804 538496 269816
rect 531792 269776 538496 269804
rect 538490 269764 538496 269776
rect 538548 269764 538554 269816
rect 538674 269764 538680 269816
rect 538732 269804 538738 269816
rect 542814 269804 542820 269816
rect 538732 269776 542820 269804
rect 538732 269764 538738 269776
rect 542814 269764 542820 269776
rect 542872 269764 542878 269816
rect 543016 269804 543044 269912
rect 543182 269900 543188 269952
rect 543240 269940 543246 269952
rect 640518 269940 640524 269952
rect 543240 269912 640524 269940
rect 543240 269900 543246 269912
rect 640518 269900 640524 269912
rect 640576 269900 640582 269952
rect 637574 269804 637580 269816
rect 543016 269776 637580 269804
rect 637574 269764 637580 269776
rect 637632 269764 637638 269816
rect 126882 269628 126888 269680
rect 126940 269668 126946 269680
rect 178310 269668 178316 269680
rect 126940 269640 178316 269668
rect 126940 269628 126946 269640
rect 178310 269628 178316 269640
rect 178368 269628 178374 269680
rect 200482 269628 200488 269680
rect 200540 269668 200546 269680
rect 226886 269668 226892 269680
rect 200540 269640 226892 269668
rect 200540 269628 200546 269640
rect 226886 269628 226892 269640
rect 226944 269628 226950 269680
rect 384758 269628 384764 269680
rect 384816 269668 384822 269680
rect 418246 269668 418252 269680
rect 384816 269640 418252 269668
rect 384816 269628 384822 269640
rect 418246 269628 418252 269640
rect 418304 269628 418310 269680
rect 422110 269628 422116 269680
rect 422168 269668 422174 269680
rect 471974 269668 471980 269680
rect 422168 269640 471980 269668
rect 422168 269628 422174 269640
rect 471974 269628 471980 269640
rect 472032 269628 472038 269680
rect 472618 269628 472624 269680
rect 472676 269668 472682 269680
rect 473354 269668 473360 269680
rect 472676 269640 473360 269668
rect 472676 269628 472682 269640
rect 473354 269628 473360 269640
rect 473412 269628 473418 269680
rect 530394 269668 530400 269680
rect 480226 269640 530400 269668
rect 78858 269492 78864 269544
rect 78916 269532 78922 269544
rect 130378 269532 130384 269544
rect 78916 269504 130384 269532
rect 78916 269492 78922 269504
rect 130378 269492 130384 269504
rect 130436 269492 130442 269544
rect 133782 269492 133788 269544
rect 133840 269532 133846 269544
rect 183646 269532 183652 269544
rect 133840 269504 183652 269532
rect 133840 269492 133846 269504
rect 183646 269492 183652 269504
rect 183704 269492 183710 269544
rect 186406 269492 186412 269544
rect 186464 269532 186470 269544
rect 204070 269532 204076 269544
rect 186464 269504 204076 269532
rect 186464 269492 186470 269504
rect 204070 269492 204076 269504
rect 204128 269492 204134 269544
rect 392026 269492 392032 269544
rect 392084 269532 392090 269544
rect 401686 269532 401692 269544
rect 392084 269504 401692 269532
rect 392084 269492 392090 269504
rect 401686 269492 401692 269504
rect 401744 269492 401750 269544
rect 404538 269492 404544 269544
rect 404596 269532 404602 269544
rect 423674 269532 423680 269544
rect 404596 269504 423680 269532
rect 404596 269492 404602 269504
rect 423674 269492 423680 269504
rect 423732 269492 423738 269544
rect 432230 269492 432236 269544
rect 432288 269532 432294 269544
rect 466454 269532 466460 269544
rect 432288 269504 466460 269532
rect 432288 269492 432294 269504
rect 466454 269492 466460 269504
rect 466512 269492 466518 269544
rect 480226 269532 480254 269640
rect 530394 269628 530400 269640
rect 530452 269628 530458 269680
rect 530578 269628 530584 269680
rect 530636 269668 530642 269680
rect 531958 269668 531964 269680
rect 530636 269640 531964 269668
rect 530636 269628 530642 269640
rect 531958 269628 531964 269640
rect 532016 269628 532022 269680
rect 533154 269628 533160 269680
rect 533212 269668 533218 269680
rect 616138 269668 616144 269680
rect 533212 269640 616144 269668
rect 533212 269628 533218 269640
rect 616138 269628 616144 269640
rect 616196 269628 616202 269680
rect 470566 269504 480254 269532
rect 140682 269356 140688 269408
rect 140740 269396 140746 269408
rect 188614 269396 188620 269408
rect 140740 269368 188620 269396
rect 140740 269356 140746 269368
rect 188614 269356 188620 269368
rect 188672 269356 188678 269408
rect 429102 269356 429108 269408
rect 429160 269396 429166 269408
rect 455414 269396 455420 269408
rect 429160 269368 455420 269396
rect 429160 269356 429166 269368
rect 455414 269356 455420 269368
rect 455472 269356 455478 269408
rect 465994 269356 466000 269408
rect 466052 269396 466058 269408
rect 470566 269396 470594 269504
rect 509050 269492 509056 269544
rect 509108 269532 509114 269544
rect 596174 269532 596180 269544
rect 509108 269504 596180 269532
rect 509108 269492 509114 269504
rect 596174 269492 596180 269504
rect 596232 269492 596238 269544
rect 466052 269368 470594 269396
rect 466052 269356 466058 269368
rect 474274 269356 474280 269408
rect 474332 269396 474338 269408
rect 538122 269396 538128 269408
rect 474332 269368 538128 269396
rect 474332 269356 474338 269368
rect 538122 269356 538128 269368
rect 538180 269356 538186 269408
rect 538306 269356 538312 269408
rect 538364 269396 538370 269408
rect 581638 269396 581644 269408
rect 538364 269368 581644 269396
rect 538364 269356 538370 269368
rect 581638 269356 581644 269368
rect 581696 269356 581702 269408
rect 121638 269220 121644 269272
rect 121696 269260 121702 269272
rect 167822 269260 167828 269272
rect 121696 269232 167828 269260
rect 121696 269220 121702 269232
rect 167822 269220 167828 269232
rect 167880 269220 167886 269272
rect 272426 269220 272432 269272
rect 272484 269260 272490 269272
rect 278866 269260 278872 269272
rect 272484 269232 278872 269260
rect 272484 269220 272490 269232
rect 278866 269220 278872 269232
rect 278924 269220 278930 269272
rect 423950 269220 423956 269272
rect 424008 269260 424014 269272
rect 448514 269260 448520 269272
rect 424008 269232 448520 269260
rect 424008 269220 424014 269232
rect 448514 269220 448520 269232
rect 448572 269220 448578 269272
rect 470962 269220 470968 269272
rect 471020 269260 471026 269272
rect 540606 269260 540612 269272
rect 471020 269232 540612 269260
rect 471020 269220 471026 269232
rect 540606 269220 540612 269232
rect 540664 269220 540670 269272
rect 540790 269220 540796 269272
rect 540848 269260 540854 269272
rect 543182 269260 543188 269272
rect 540848 269232 543188 269260
rect 540848 269220 540854 269232
rect 543182 269220 543188 269232
rect 543240 269220 543246 269272
rect 543366 269152 543372 269204
rect 543424 269192 543430 269204
rect 546494 269192 546500 269204
rect 543424 269164 546500 269192
rect 543424 269152 543430 269164
rect 546494 269152 546500 269164
rect 546552 269152 546558 269204
rect 274910 269084 274916 269136
rect 274968 269124 274974 269136
rect 279694 269124 279700 269136
rect 274968 269096 279700 269124
rect 274968 269084 274974 269096
rect 279694 269084 279700 269096
rect 279752 269084 279758 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 42150 269016 42156 269068
rect 42208 269056 42214 269068
rect 43162 269056 43168 269068
rect 42208 269028 43168 269056
rect 42208 269016 42214 269028
rect 43162 269016 43168 269028
rect 43220 269016 43226 269068
rect 84102 269016 84108 269068
rect 84160 269056 84166 269068
rect 137462 269056 137468 269068
rect 84160 269028 137468 269056
rect 84160 269016 84166 269028
rect 137462 269016 137468 269028
rect 137520 269016 137526 269068
rect 137646 269016 137652 269068
rect 137704 269056 137710 269068
rect 186130 269056 186136 269068
rect 137704 269028 186136 269056
rect 137704 269016 137710 269028
rect 186130 269016 186136 269028
rect 186188 269016 186194 269068
rect 379698 269016 379704 269068
rect 379756 269056 379762 269068
rect 404354 269056 404360 269068
rect 379756 269028 404360 269056
rect 379756 269016 379762 269028
rect 404354 269016 404360 269028
rect 404412 269016 404418 269068
rect 436186 269016 436192 269068
rect 436244 269056 436250 269068
rect 491754 269056 491760 269068
rect 436244 269028 491760 269056
rect 436244 269016 436250 269028
rect 491754 269016 491760 269028
rect 491812 269016 491818 269068
rect 498286 269016 498292 269068
rect 498344 269056 498350 269068
rect 580994 269056 581000 269068
rect 498344 269028 581000 269056
rect 498344 269016 498350 269028
rect 580994 269016 581000 269028
rect 581052 269016 581058 269068
rect 273254 268948 273260 269000
rect 273312 268988 273318 269000
rect 275554 268988 275560 269000
rect 273312 268960 275560 268988
rect 273312 268948 273318 268960
rect 275554 268948 275560 268960
rect 275612 268948 275618 269000
rect 111978 268880 111984 268932
rect 112036 268920 112042 268932
rect 168742 268920 168748 268932
rect 112036 268892 168748 268920
rect 112036 268880 112042 268892
rect 168742 268880 168748 268892
rect 168800 268880 168806 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 415394 268920 415400 268932
rect 382424 268892 415400 268920
rect 382424 268880 382430 268892
rect 415394 268880 415400 268892
rect 415452 268880 415458 268932
rect 433702 268880 433708 268932
rect 433760 268920 433766 268932
rect 488534 268920 488540 268932
rect 433760 268892 488540 268920
rect 433760 268880 433766 268892
rect 488534 268880 488540 268892
rect 488592 268880 488598 268932
rect 500770 268880 500776 268932
rect 500828 268920 500834 268932
rect 583754 268920 583760 268932
rect 500828 268892 583760 268920
rect 500828 268880 500834 268892
rect 583754 268880 583760 268892
rect 583812 268880 583818 268932
rect 115842 268744 115848 268796
rect 115900 268784 115906 268796
rect 115900 268756 166304 268784
rect 115900 268744 115906 268756
rect 110230 268608 110236 268660
rect 110288 268648 110294 268660
rect 110288 268620 164648 268648
rect 110288 268608 110294 268620
rect 102502 268472 102508 268524
rect 102560 268512 102566 268524
rect 162946 268512 162952 268524
rect 102560 268484 162952 268512
rect 102560 268472 102566 268484
rect 162946 268472 162952 268484
rect 163004 268472 163010 268524
rect 92382 268336 92388 268388
rect 92440 268376 92446 268388
rect 155494 268376 155500 268388
rect 92440 268348 155500 268376
rect 92440 268336 92446 268348
rect 155494 268336 155500 268348
rect 155552 268336 155558 268388
rect 164620 268376 164648 268620
rect 166276 268512 166304 268756
rect 211338 268744 211344 268796
rect 211396 268784 211402 268796
rect 223482 268784 223488 268796
rect 211396 268756 223488 268784
rect 211396 268744 211402 268756
rect 223482 268744 223488 268756
rect 223540 268744 223546 268796
rect 389818 268744 389824 268796
rect 389876 268784 389882 268796
rect 425330 268784 425336 268796
rect 389876 268756 425336 268784
rect 389876 268744 389882 268756
rect 425330 268744 425336 268756
rect 425388 268744 425394 268796
rect 441154 268744 441160 268796
rect 441212 268784 441218 268796
rect 499574 268784 499580 268796
rect 441212 268756 499580 268784
rect 441212 268744 441218 268756
rect 499574 268744 499580 268756
rect 499632 268744 499638 268796
rect 503254 268744 503260 268796
rect 503312 268784 503318 268796
rect 587894 268784 587900 268796
rect 503312 268756 587900 268784
rect 503312 268744 503318 268756
rect 587894 268744 587900 268756
rect 587952 268744 587958 268796
rect 166994 268608 167000 268660
rect 167052 268648 167058 268660
rect 184474 268648 184480 268660
rect 167052 268620 184480 268648
rect 167052 268608 167058 268620
rect 184474 268608 184480 268620
rect 184532 268608 184538 268660
rect 187326 268608 187332 268660
rect 187384 268648 187390 268660
rect 219434 268648 219440 268660
rect 187384 268620 219440 268648
rect 187384 268608 187390 268620
rect 219434 268608 219440 268620
rect 219492 268608 219498 268660
rect 245562 268608 245568 268660
rect 245620 268648 245626 268660
rect 263134 268648 263140 268660
rect 245620 268620 263140 268648
rect 245620 268608 245626 268620
rect 263134 268608 263140 268620
rect 263192 268608 263198 268660
rect 403250 268608 403256 268660
rect 403308 268648 403314 268660
rect 440234 268648 440240 268660
rect 403308 268620 440240 268648
rect 403308 268608 403314 268620
rect 440234 268608 440240 268620
rect 440292 268608 440298 268660
rect 443638 268608 443644 268660
rect 443696 268648 443702 268660
rect 502334 268648 502340 268660
rect 443696 268620 502340 268648
rect 443696 268608 443702 268620
rect 502334 268608 502340 268620
rect 502392 268608 502398 268660
rect 505738 268608 505744 268660
rect 505796 268648 505802 268660
rect 590838 268648 590844 268660
rect 505796 268620 590844 268648
rect 505796 268608 505802 268620
rect 590838 268608 590844 268620
rect 590896 268608 590902 268660
rect 171226 268512 171232 268524
rect 166276 268484 171232 268512
rect 171226 268472 171232 268484
rect 171284 268472 171290 268524
rect 176930 268472 176936 268524
rect 176988 268512 176994 268524
rect 215110 268512 215116 268524
rect 176988 268484 215116 268512
rect 176988 268472 176994 268484
rect 215110 268472 215116 268484
rect 215168 268472 215174 268524
rect 220446 268472 220452 268524
rect 220504 268512 220510 268524
rect 245746 268512 245752 268524
rect 220504 268484 245752 268512
rect 220504 268472 220510 268484
rect 245746 268472 245752 268484
rect 245804 268472 245810 268524
rect 338482 268472 338488 268524
rect 338540 268512 338546 268524
rect 350718 268512 350724 268524
rect 338540 268484 350724 268512
rect 338540 268472 338546 268484
rect 350718 268472 350724 268484
rect 350776 268472 350782 268524
rect 359826 268472 359832 268524
rect 359884 268512 359890 268524
rect 379514 268512 379520 268524
rect 359884 268484 379520 268512
rect 359884 268472 359890 268484
rect 379514 268472 379520 268484
rect 379572 268472 379578 268524
rect 397086 268472 397092 268524
rect 397144 268512 397150 268524
rect 433334 268512 433340 268524
rect 397144 268484 433340 268512
rect 397144 268472 397150 268484
rect 433334 268472 433340 268484
rect 433392 268472 433398 268524
rect 448606 268472 448612 268524
rect 448664 268512 448670 268524
rect 509234 268512 509240 268524
rect 448664 268484 509240 268512
rect 448664 268472 448670 268484
rect 509234 268472 509240 268484
rect 509292 268472 509298 268524
rect 513190 268472 513196 268524
rect 513248 268512 513254 268524
rect 601694 268512 601700 268524
rect 513248 268484 601700 268512
rect 513248 268472 513254 268484
rect 601694 268472 601700 268484
rect 601752 268472 601758 268524
rect 167638 268376 167644 268388
rect 164620 268348 167644 268376
rect 167638 268336 167644 268348
rect 167696 268336 167702 268388
rect 168006 268336 168012 268388
rect 168064 268376 168070 268388
rect 203518 268376 203524 268388
rect 168064 268348 203524 268376
rect 168064 268336 168070 268348
rect 203518 268336 203524 268348
rect 203576 268336 203582 268388
rect 203886 268336 203892 268388
rect 203944 268376 203950 268388
rect 230750 268376 230756 268388
rect 203944 268348 230756 268376
rect 203944 268336 203950 268348
rect 230750 268336 230756 268348
rect 230808 268336 230814 268388
rect 231670 268336 231676 268388
rect 231728 268376 231734 268388
rect 253198 268376 253204 268388
rect 231728 268348 253204 268376
rect 231728 268336 231734 268348
rect 253198 268336 253204 268348
rect 253256 268336 253262 268388
rect 258350 268336 258356 268388
rect 258408 268376 258414 268388
rect 268930 268376 268936 268388
rect 258408 268348 268936 268376
rect 258408 268336 258414 268348
rect 268930 268336 268936 268348
rect 268988 268336 268994 268388
rect 348418 268336 348424 268388
rect 348476 268376 348482 268388
rect 367094 268376 367100 268388
rect 348476 268348 367100 268376
rect 348476 268336 348482 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 372154 268336 372160 268388
rect 372212 268376 372218 268388
rect 397454 268376 397460 268388
rect 372212 268348 397460 268376
rect 372212 268336 372218 268348
rect 397454 268336 397460 268348
rect 397512 268336 397518 268388
rect 408034 268336 408040 268388
rect 408092 268376 408098 268388
rect 451366 268376 451372 268388
rect 408092 268348 451372 268376
rect 408092 268336 408098 268348
rect 451366 268336 451372 268348
rect 451424 268336 451430 268388
rect 464338 268336 464344 268388
rect 464396 268376 464402 268388
rect 532694 268376 532700 268388
rect 464396 268348 532700 268376
rect 464396 268336 464402 268348
rect 532694 268336 532700 268348
rect 532752 268336 532758 268388
rect 541342 268336 541348 268388
rect 541400 268376 541406 268388
rect 641714 268376 641720 268388
rect 541400 268348 641720 268376
rect 541400 268336 541406 268348
rect 641714 268336 641720 268348
rect 641772 268336 641778 268388
rect 128538 268200 128544 268252
rect 128596 268240 128602 268252
rect 150434 268240 150440 268252
rect 128596 268212 150440 268240
rect 128596 268200 128602 268212
rect 150434 268200 150440 268212
rect 150492 268200 150498 268252
rect 151722 268200 151728 268252
rect 151780 268240 151786 268252
rect 196066 268240 196072 268252
rect 151780 268212 196072 268240
rect 151780 268200 151786 268212
rect 196066 268200 196072 268212
rect 196124 268200 196130 268252
rect 419626 268200 419632 268252
rect 419684 268240 419690 268252
rect 467926 268240 467932 268252
rect 419684 268212 467932 268240
rect 419684 268200 419690 268212
rect 467926 268200 467932 268212
rect 467984 268200 467990 268252
rect 493594 268200 493600 268252
rect 493652 268240 493658 268252
rect 574094 268240 574100 268252
rect 493652 268212 574100 268240
rect 493652 268200 493658 268212
rect 574094 268200 574100 268212
rect 574152 268200 574158 268252
rect 163130 268064 163136 268116
rect 163188 268104 163194 268116
rect 168006 268104 168012 268116
rect 163188 268076 168012 268104
rect 163188 268064 163194 268076
rect 168006 268064 168012 268076
rect 168064 268064 168070 268116
rect 412634 268064 412640 268116
rect 412692 268104 412698 268116
rect 447134 268104 447140 268116
rect 412692 268076 447140 268104
rect 412692 268064 412698 268076
rect 447134 268064 447140 268076
rect 447192 268064 447198 268116
rect 495802 268064 495808 268116
rect 495860 268104 495866 268116
rect 576854 268104 576860 268116
rect 495860 268076 576860 268104
rect 495860 268064 495866 268076
rect 576854 268064 576860 268076
rect 576912 268064 576918 268116
rect 198734 267792 198740 267844
rect 198792 267832 198798 267844
rect 201862 267832 201868 267844
rect 198792 267804 201868 267832
rect 198792 267792 198798 267804
rect 201862 267792 201868 267804
rect 201920 267792 201926 267844
rect 117958 267656 117964 267708
rect 118016 267696 118022 267708
rect 159634 267696 159640 267708
rect 118016 267668 159640 267696
rect 118016 267656 118022 267668
rect 159634 267656 159640 267668
rect 159692 267656 159698 267708
rect 167822 267656 167828 267708
rect 167880 267696 167886 267708
rect 177022 267696 177028 267708
rect 167880 267668 177028 267696
rect 167880 267656 167886 267668
rect 177022 267656 177028 267668
rect 177080 267656 177086 267708
rect 181990 267656 181996 267708
rect 182048 267696 182054 267708
rect 182048 267668 182312 267696
rect 182048 267656 182054 267668
rect 95878 267520 95884 267572
rect 95936 267560 95942 267572
rect 138106 267560 138112 267572
rect 95936 267532 138112 267560
rect 95936 267520 95942 267532
rect 138106 267520 138112 267532
rect 138164 267520 138170 267572
rect 150434 267520 150440 267572
rect 150492 267560 150498 267572
rect 181990 267560 181996 267572
rect 150492 267532 181996 267560
rect 150492 267520 150498 267532
rect 181990 267520 181996 267532
rect 182048 267520 182054 267572
rect 182284 267560 182312 267668
rect 182726 267656 182732 267708
rect 182784 267696 182790 267708
rect 214282 267696 214288 267708
rect 182784 267668 214288 267696
rect 182784 267656 182790 267668
rect 214282 267656 214288 267668
rect 214340 267656 214346 267708
rect 378226 267656 378232 267708
rect 378284 267696 378290 267708
rect 392578 267696 392584 267708
rect 378284 267668 392584 267696
rect 378284 267656 378290 267668
rect 392578 267656 392584 267668
rect 392636 267656 392642 267708
rect 398098 267656 398104 267708
rect 398156 267696 398162 267708
rect 414474 267696 414480 267708
rect 398156 267668 414480 267696
rect 398156 267656 398162 267668
rect 414474 267656 414480 267668
rect 414532 267656 414538 267708
rect 423766 267656 423772 267708
rect 423824 267696 423830 267708
rect 440878 267696 440884 267708
rect 423824 267668 440884 267696
rect 423824 267656 423830 267668
rect 440878 267656 440884 267668
rect 440936 267656 440942 267708
rect 442718 267656 442724 267708
rect 442776 267696 442782 267708
rect 493318 267696 493324 267708
rect 442776 267668 493324 267696
rect 442776 267656 442782 267668
rect 493318 267656 493324 267668
rect 493376 267656 493382 267708
rect 497826 267656 497832 267708
rect 497884 267696 497890 267708
rect 517514 267696 517520 267708
rect 497884 267668 517520 267696
rect 497884 267656 497890 267668
rect 517514 267656 517520 267668
rect 517572 267656 517578 267708
rect 529658 267656 529664 267708
rect 529716 267696 529722 267708
rect 585778 267696 585784 267708
rect 529716 267668 585784 267696
rect 529716 267656 529722 267668
rect 585778 267656 585784 267668
rect 585836 267656 585842 267708
rect 219250 267560 219256 267572
rect 182284 267532 219256 267560
rect 219250 267520 219256 267532
rect 219308 267520 219314 267572
rect 340966 267520 340972 267572
rect 341024 267560 341030 267572
rect 355318 267560 355324 267572
rect 341024 267532 355324 267560
rect 341024 267520 341030 267532
rect 355318 267520 355324 267532
rect 355376 267520 355382 267572
rect 370774 267520 370780 267572
rect 370832 267560 370838 267572
rect 377398 267560 377404 267572
rect 370832 267532 377404 267560
rect 370832 267520 370838 267532
rect 377398 267520 377404 267532
rect 377456 267520 377462 267572
rect 380710 267520 380716 267572
rect 380768 267560 380774 267572
rect 399846 267560 399852 267572
rect 380768 267532 399852 267560
rect 380768 267520 380774 267532
rect 399846 267520 399852 267532
rect 399904 267520 399910 267572
rect 410518 267520 410524 267572
rect 410576 267560 410582 267572
rect 429102 267560 429108 267572
rect 410576 267532 429108 267560
rect 410576 267520 410582 267532
rect 429102 267520 429108 267532
rect 429160 267520 429166 267572
rect 445294 267520 445300 267572
rect 445352 267560 445358 267572
rect 497458 267560 497464 267572
rect 445352 267532 497464 267560
rect 445352 267520 445358 267532
rect 497458 267520 497464 267532
rect 497516 267520 497522 267572
rect 514846 267520 514852 267572
rect 514904 267560 514910 267572
rect 571978 267560 571984 267572
rect 514904 267532 571984 267560
rect 514904 267520 514910 267532
rect 571978 267520 571984 267532
rect 572036 267520 572042 267572
rect 86218 267384 86224 267436
rect 86276 267424 86282 267436
rect 144730 267424 144736 267436
rect 86276 267396 144736 267424
rect 86276 267384 86282 267396
rect 144730 267384 144736 267396
rect 144788 267384 144794 267436
rect 146938 267384 146944 267436
rect 146996 267424 147002 267436
rect 186958 267424 186964 267436
rect 146996 267396 186964 267424
rect 146996 267384 147002 267396
rect 186958 267384 186964 267396
rect 187016 267384 187022 267436
rect 236638 267384 236644 267436
rect 236696 267424 236702 267436
rect 241606 267424 241612 267436
rect 236696 267396 241612 267424
rect 236696 267384 236702 267396
rect 241606 267384 241612 267396
rect 241664 267384 241670 267436
rect 315298 267384 315304 267436
rect 315356 267424 315362 267436
rect 318978 267424 318984 267436
rect 315356 267396 318984 267424
rect 315356 267384 315362 267396
rect 318978 267384 318984 267396
rect 319036 267384 319042 267436
rect 350074 267384 350080 267436
rect 350132 267424 350138 267436
rect 358078 267424 358084 267436
rect 350132 267396 358084 267424
rect 350132 267384 350138 267396
rect 358078 267384 358084 267396
rect 358136 267384 358142 267436
rect 362494 267384 362500 267436
rect 362552 267424 362558 267436
rect 369302 267424 369308 267436
rect 362552 267396 369308 267424
rect 362552 267384 362558 267396
rect 369302 267384 369308 267396
rect 369360 267384 369366 267436
rect 371602 267384 371608 267436
rect 371660 267424 371666 267436
rect 373258 267424 373264 267436
rect 371660 267396 373264 267424
rect 371660 267384 371666 267396
rect 373258 267384 373264 267396
rect 373316 267384 373322 267436
rect 383194 267384 383200 267436
rect 383252 267424 383258 267436
rect 401870 267424 401876 267436
rect 383252 267396 401876 267424
rect 383252 267384 383258 267396
rect 401870 267384 401876 267396
rect 401928 267384 401934 267436
rect 405550 267384 405556 267436
rect 405608 267424 405614 267436
rect 423950 267424 423956 267436
rect 405608 267396 423956 267424
rect 405608 267384 405614 267396
rect 423950 267384 423956 267396
rect 424008 267384 424014 267436
rect 432046 267384 432052 267436
rect 432104 267424 432110 267436
rect 453298 267424 453304 267436
rect 432104 267396 453304 267424
rect 432104 267384 432110 267396
rect 453298 267384 453304 267396
rect 453356 267384 453362 267436
rect 460198 267384 460204 267436
rect 460256 267424 460262 267436
rect 515398 267424 515404 267436
rect 460256 267396 515404 267424
rect 460256 267384 460262 267396
rect 515398 267384 515404 267396
rect 515456 267384 515462 267436
rect 519814 267384 519820 267436
rect 519872 267424 519878 267436
rect 578878 267424 578884 267436
rect 519872 267396 578884 267424
rect 519872 267384 519878 267396
rect 578878 267384 578884 267396
rect 578936 267384 578942 267436
rect 104802 267248 104808 267300
rect 104860 267288 104866 267300
rect 164602 267288 164608 267300
rect 104860 267260 164608 267288
rect 104860 267248 104866 267260
rect 164602 267248 164608 267260
rect 164660 267248 164666 267300
rect 169018 267248 169024 267300
rect 169076 267288 169082 267300
rect 209314 267288 209320 267300
rect 169076 267260 209320 267288
rect 169076 267248 169082 267260
rect 209314 267248 209320 267260
rect 209372 267248 209378 267300
rect 218698 267248 218704 267300
rect 218756 267288 218762 267300
rect 223022 267288 223028 267300
rect 218756 267260 223028 267288
rect 218756 267248 218762 267260
rect 223022 267248 223028 267260
rect 223080 267248 223086 267300
rect 223482 267248 223488 267300
rect 223540 267288 223546 267300
rect 239122 267288 239128 267300
rect 223540 267260 239128 267288
rect 223540 267248 223546 267260
rect 239122 267248 239128 267260
rect 239180 267248 239186 267300
rect 314470 267248 314476 267300
rect 314528 267288 314534 267300
rect 318794 267288 318800 267300
rect 314528 267260 318800 267288
rect 314528 267248 314534 267260
rect 318794 267248 318800 267260
rect 318852 267248 318858 267300
rect 353386 267248 353392 267300
rect 353444 267288 353450 267300
rect 364978 267288 364984 267300
rect 353444 267260 364984 267288
rect 353444 267248 353450 267260
rect 364978 267248 364984 267260
rect 365036 267248 365042 267300
rect 373258 267248 373264 267300
rect 373316 267288 373322 267300
rect 392026 267288 392032 267300
rect 373316 267260 392032 267288
rect 373316 267248 373322 267260
rect 392026 267248 392032 267260
rect 392084 267248 392090 267300
rect 403066 267248 403072 267300
rect 403124 267288 403130 267300
rect 422938 267288 422944 267300
rect 403124 267260 422944 267288
rect 403124 267248 403130 267260
rect 422938 267248 422944 267260
rect 422996 267248 423002 267300
rect 424594 267248 424600 267300
rect 424652 267288 424658 267300
rect 446398 267288 446404 267300
rect 424652 267260 446404 267288
rect 424652 267248 424658 267260
rect 446398 267248 446404 267260
rect 446456 267248 446462 267300
rect 448146 267248 448152 267300
rect 448204 267288 448210 267300
rect 457438 267288 457444 267300
rect 448204 267260 457444 267288
rect 448204 267248 448210 267260
rect 457438 267248 457444 267260
rect 457496 267248 457502 267300
rect 470134 267248 470140 267300
rect 470192 267288 470198 267300
rect 534718 267288 534724 267300
rect 470192 267260 534724 267288
rect 470192 267248 470198 267260
rect 534718 267248 534724 267260
rect 534776 267248 534782 267300
rect 542998 267248 543004 267300
rect 543056 267288 543062 267300
rect 625798 267288 625804 267300
rect 543056 267260 625804 267288
rect 543056 267248 543062 267260
rect 625798 267248 625804 267260
rect 625856 267248 625862 267300
rect 79962 267112 79968 267164
rect 80020 267152 80026 267164
rect 140590 267152 140596 267164
rect 80020 267124 140596 267152
rect 80020 267112 80026 267124
rect 140590 267112 140596 267124
rect 140648 267112 140654 267164
rect 144178 267112 144184 267164
rect 144236 267152 144242 267164
rect 191926 267152 191932 267164
rect 144236 267124 191932 267152
rect 144236 267112 144242 267124
rect 191926 267112 191932 267124
rect 191984 267112 191990 267164
rect 192570 267112 192576 267164
rect 192628 267152 192634 267164
rect 223942 267152 223948 267164
rect 192628 267124 223948 267152
rect 192628 267112 192634 267124
rect 223942 267112 223948 267124
rect 224000 267112 224006 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 312814 267112 312820 267164
rect 312872 267152 312878 267164
rect 316034 267152 316040 267164
rect 312872 267124 316040 267152
rect 312872 267112 312878 267124
rect 316034 267112 316040 267124
rect 316092 267112 316098 267164
rect 365806 267112 365812 267164
rect 365864 267152 365870 267164
rect 382918 267152 382924 267164
rect 365864 267124 382924 267152
rect 365864 267112 365870 267124
rect 382918 267112 382924 267124
rect 382976 267112 382982 267164
rect 390646 267112 390652 267164
rect 390704 267152 390710 267164
rect 417418 267152 417424 267164
rect 390704 267124 417424 267152
rect 390704 267112 390710 267124
rect 417418 267112 417424 267124
rect 417476 267112 417482 267164
rect 417970 267112 417976 267164
rect 418028 267152 418034 267164
rect 432230 267152 432236 267164
rect 418028 267124 432236 267152
rect 418028 267112 418034 267124
rect 432230 267112 432236 267124
rect 432288 267112 432294 267164
rect 432874 267112 432880 267164
rect 432932 267152 432938 267164
rect 460014 267152 460020 267164
rect 432932 267124 460020 267152
rect 432932 267112 432938 267124
rect 460014 267112 460020 267124
rect 460072 267112 460078 267164
rect 465166 267112 465172 267164
rect 465224 267152 465230 267164
rect 526438 267152 526444 267164
rect 465224 267124 526444 267152
rect 465224 267112 465230 267124
rect 526438 267112 526444 267124
rect 526496 267112 526502 267164
rect 534718 267112 534724 267164
rect 534776 267152 534782 267164
rect 618898 267152 618904 267164
rect 534776 267124 618904 267152
rect 534776 267112 534782 267124
rect 618898 267112 618904 267124
rect 618956 267112 618962 267164
rect 90358 266976 90364 267028
rect 90416 267016 90422 267028
rect 151354 267016 151360 267028
rect 90416 266988 151360 267016
rect 90416 266976 90422 266988
rect 151354 266976 151360 266988
rect 151412 266976 151418 267028
rect 154482 266976 154488 267028
rect 154540 267016 154546 267028
rect 199378 267016 199384 267028
rect 154540 266988 199384 267016
rect 154540 266976 154546 266988
rect 199378 266976 199384 266988
rect 199436 266976 199442 267028
rect 218882 266976 218888 267028
rect 218940 267016 218946 267028
rect 220078 267016 220084 267028
rect 218940 266988 220084 267016
rect 218940 266976 218946 266988
rect 220078 266976 220084 266988
rect 220136 266976 220142 267028
rect 228358 266976 228364 267028
rect 228416 267016 228422 267028
rect 228416 266988 238754 267016
rect 228416 266976 228422 266988
rect 121454 266840 121460 266892
rect 121512 266880 121518 266892
rect 144914 266880 144920 266892
rect 121512 266852 144920 266880
rect 121512 266840 121518 266852
rect 144914 266840 144920 266852
rect 144972 266840 144978 266892
rect 145374 266840 145380 266892
rect 145432 266880 145438 266892
rect 150526 266880 150532 266892
rect 145432 266852 150532 266880
rect 145432 266840 145438 266852
rect 150526 266840 150532 266852
rect 150584 266840 150590 266892
rect 204070 266840 204076 266892
rect 204128 266880 204134 266892
rect 220906 266880 220912 266892
rect 204128 266852 220912 266880
rect 204128 266840 204134 266852
rect 220906 266840 220912 266852
rect 220964 266840 220970 266892
rect 238726 266880 238754 266988
rect 316954 266976 316960 267028
rect 317012 267016 317018 267028
rect 321922 267016 321928 267028
rect 317012 266988 321928 267016
rect 317012 266976 317018 266988
rect 321922 266976 321928 266988
rect 321980 266976 321986 267028
rect 375742 266976 375748 267028
rect 375800 267016 375806 267028
rect 390094 267016 390100 267028
rect 375800 266988 390100 267016
rect 375800 266976 375806 266988
rect 390094 266976 390100 266988
rect 390152 266976 390158 267028
rect 393130 266976 393136 267028
rect 393188 267016 393194 267028
rect 420178 267016 420184 267028
rect 393188 266988 420184 267016
rect 393188 266976 393194 266988
rect 420178 266976 420184 266988
rect 420236 266976 420242 267028
rect 431218 266976 431224 267028
rect 431276 267016 431282 267028
rect 432598 267016 432604 267028
rect 431276 266988 432604 267016
rect 431276 266976 431282 266988
rect 432598 266976 432604 266988
rect 432656 266976 432662 267028
rect 450538 267016 450544 267028
rect 441586 266988 450544 267016
rect 249058 266880 249064 266892
rect 238726 266852 249064 266880
rect 249058 266840 249064 266852
rect 249116 266840 249122 266892
rect 286318 266840 286324 266892
rect 286376 266880 286382 266892
rect 287974 266880 287980 266892
rect 286376 266852 287980 266880
rect 286376 266840 286382 266852
rect 287974 266840 287980 266852
rect 288032 266840 288038 266892
rect 321922 266840 321928 266892
rect 321980 266880 321986 266892
rect 327534 266880 327540 266892
rect 321980 266852 327540 266880
rect 321980 266840 321986 266852
rect 327534 266840 327540 266852
rect 327592 266840 327598 266892
rect 332686 266840 332692 266892
rect 332744 266880 332750 266892
rect 343818 266880 343824 266892
rect 332744 266852 343824 266880
rect 332744 266840 332750 266852
rect 343818 266840 343824 266852
rect 343876 266840 343882 266892
rect 392302 266840 392308 266892
rect 392360 266880 392366 266892
rect 393958 266880 393964 266892
rect 392360 266852 393964 266880
rect 392360 266840 392366 266852
rect 393958 266840 393964 266852
rect 394016 266840 394022 266892
rect 427906 266840 427912 266892
rect 427964 266880 427970 266892
rect 441586 266880 441614 266988
rect 450538 266976 450544 266988
rect 450596 266976 450602 267028
rect 455046 266976 455052 267028
rect 455104 267016 455110 267028
rect 512638 267016 512644 267028
rect 455104 266988 512644 267016
rect 455104 266976 455110 266988
rect 512638 266976 512644 266988
rect 512696 266976 512702 267028
rect 524782 266976 524788 267028
rect 524840 267016 524846 267028
rect 611998 267016 612004 267028
rect 524840 266988 612004 267016
rect 524840 266976 524846 266988
rect 611998 266976 612004 266988
rect 612056 266976 612062 267028
rect 427964 266852 441614 266880
rect 427964 266840 427970 266852
rect 450262 266840 450268 266892
rect 450320 266880 450326 266892
rect 450320 266852 489914 266880
rect 450320 266840 450326 266852
rect 355870 266772 355876 266824
rect 355928 266812 355934 266824
rect 374638 266812 374644 266824
rect 355928 266784 374644 266812
rect 355928 266772 355934 266784
rect 374638 266772 374644 266784
rect 374696 266772 374702 266824
rect 130378 266704 130384 266756
rect 130436 266744 130442 266756
rect 147214 266744 147220 266756
rect 130436 266716 147220 266744
rect 130436 266704 130442 266716
rect 147214 266704 147220 266716
rect 147272 266704 147278 266756
rect 149698 266704 149704 266756
rect 149756 266744 149762 266756
rect 169570 266744 169576 266756
rect 149756 266716 169576 266744
rect 149756 266704 149762 266716
rect 169570 266704 169576 266716
rect 169628 266704 169634 266756
rect 230750 266704 230756 266756
rect 230808 266744 230814 266756
rect 234154 266744 234160 266756
rect 230808 266716 234160 266744
rect 230808 266704 230814 266716
rect 234154 266704 234160 266716
rect 234212 266704 234218 266756
rect 252002 266704 252008 266756
rect 252060 266744 252066 266756
rect 258994 266744 259000 266756
rect 252060 266716 259000 266744
rect 252060 266704 252066 266716
rect 258994 266704 259000 266716
rect 259052 266704 259058 266756
rect 313642 266704 313648 266756
rect 313700 266744 313706 266756
rect 317414 266744 317420 266756
rect 313700 266716 317420 266744
rect 313700 266704 313706 266716
rect 317414 266704 317420 266716
rect 317472 266704 317478 266756
rect 388162 266704 388168 266756
rect 388220 266744 388226 266756
rect 388220 266716 393314 266744
rect 388220 266704 388226 266716
rect 214558 266636 214564 266688
rect 214616 266676 214622 266688
rect 218422 266676 218428 266688
rect 214616 266648 218428 266676
rect 214616 266636 214622 266648
rect 218422 266636 218428 266648
rect 218480 266636 218486 266688
rect 308674 266636 308680 266688
rect 308732 266676 308738 266688
rect 310514 266676 310520 266688
rect 308732 266648 310520 266676
rect 308732 266636 308738 266648
rect 310514 266636 310520 266648
rect 310572 266636 310578 266688
rect 317782 266636 317788 266688
rect 317840 266676 317846 266688
rect 322934 266676 322940 266688
rect 317840 266648 322940 266676
rect 317840 266636 317846 266648
rect 322934 266636 322940 266648
rect 322992 266636 322998 266688
rect 342622 266636 342628 266688
rect 342680 266676 342686 266688
rect 347038 266676 347044 266688
rect 342680 266648 347044 266676
rect 342680 266636 342686 266648
rect 347038 266636 347044 266648
rect 347096 266636 347102 266688
rect 137462 266568 137468 266620
rect 137520 266608 137526 266620
rect 145374 266608 145380 266620
rect 137520 266580 145380 266608
rect 137520 266568 137526 266580
rect 145374 266568 145380 266580
rect 145432 266568 145438 266620
rect 145558 266568 145564 266620
rect 145616 266608 145622 266620
rect 148042 266608 148048 266620
rect 145616 266580 148048 266608
rect 145616 266568 145622 266580
rect 148042 266568 148048 266580
rect 148100 266568 148106 266620
rect 226886 266568 226892 266620
rect 226944 266608 226950 266620
rect 231670 266608 231676 266620
rect 226944 266580 231676 266608
rect 226944 266568 226950 266580
rect 231670 266568 231676 266580
rect 231728 266568 231734 266620
rect 393286 266608 393314 266716
rect 394786 266704 394792 266756
rect 394844 266744 394850 266756
rect 397086 266744 397092 266756
rect 394844 266716 397092 266744
rect 394844 266704 394850 266716
rect 397086 266704 397092 266716
rect 397144 266704 397150 266756
rect 397454 266704 397460 266756
rect 397512 266744 397518 266756
rect 407758 266744 407764 266756
rect 397512 266716 407764 266744
rect 397512 266704 397518 266716
rect 407758 266704 407764 266716
rect 407816 266704 407822 266756
rect 428734 266704 428740 266756
rect 428792 266744 428798 266756
rect 428792 266716 431954 266744
rect 428792 266704 428798 266716
rect 404538 266608 404544 266620
rect 393286 266580 404544 266608
rect 404538 266568 404544 266580
rect 404596 266568 404602 266620
rect 404722 266568 404728 266620
rect 404780 266608 404786 266620
rect 412634 266608 412640 266620
rect 404780 266580 412640 266608
rect 404780 266568 404786 266580
rect 412634 266568 412640 266580
rect 412692 266568 412698 266620
rect 431926 266608 431954 266716
rect 440326 266704 440332 266756
rect 440384 266744 440390 266756
rect 445018 266744 445024 266756
rect 440384 266716 445024 266744
rect 440384 266704 440390 266716
rect 445018 266704 445024 266716
rect 445076 266704 445082 266756
rect 457714 266704 457720 266756
rect 457772 266744 457778 266756
rect 479518 266744 479524 266756
rect 457772 266716 479524 266744
rect 457772 266704 457778 266716
rect 479518 266704 479524 266716
rect 479576 266704 479582 266756
rect 442258 266608 442264 266620
rect 431926 266580 442264 266608
rect 442258 266568 442264 266580
rect 442316 266568 442322 266620
rect 452746 266568 452752 266620
rect 452804 266608 452810 266620
rect 469858 266608 469864 266620
rect 452804 266580 469864 266608
rect 452804 266568 452810 266580
rect 469858 266568 469864 266580
rect 469916 266568 469922 266620
rect 489886 266608 489914 266852
rect 504818 266840 504824 266892
rect 504876 266880 504882 266892
rect 513926 266880 513932 266892
rect 504876 266852 513932 266880
rect 504876 266840 504882 266852
rect 513926 266840 513932 266852
rect 513984 266840 513990 266892
rect 514128 266852 518894 266880
rect 490006 266704 490012 266756
rect 490064 266744 490070 266756
rect 507118 266744 507124 266756
rect 490064 266716 507124 266744
rect 490064 266704 490070 266716
rect 507118 266704 507124 266716
rect 507176 266704 507182 266756
rect 509878 266704 509884 266756
rect 509936 266744 509942 266756
rect 514128 266744 514156 266852
rect 509936 266716 514156 266744
rect 509936 266704 509942 266716
rect 516502 266704 516508 266756
rect 516560 266744 516566 266756
rect 517330 266744 517336 266756
rect 516560 266716 517336 266744
rect 516560 266704 516566 266716
rect 517330 266704 517336 266716
rect 517388 266704 517394 266756
rect 518866 266744 518894 266852
rect 518986 266840 518992 266892
rect 519044 266880 519050 266892
rect 520090 266880 520096 266892
rect 519044 266852 520096 266880
rect 519044 266840 519050 266852
rect 520090 266840 520096 266852
rect 520148 266840 520154 266892
rect 527266 266840 527272 266892
rect 527324 266880 527330 266892
rect 528186 266880 528192 266892
rect 527324 266852 528192 266880
rect 527324 266840 527330 266852
rect 528186 266840 528192 266852
rect 528244 266840 528250 266892
rect 528922 266840 528928 266892
rect 528980 266880 528986 266892
rect 529842 266880 529848 266892
rect 528980 266852 529848 266880
rect 528980 266840 528986 266852
rect 529842 266840 529848 266852
rect 529900 266840 529906 266892
rect 531406 266840 531412 266892
rect 531464 266880 531470 266892
rect 532510 266880 532516 266892
rect 531464 266852 532516 266880
rect 531464 266840 531470 266852
rect 532510 266840 532516 266852
rect 532568 266840 532574 266892
rect 533062 266840 533068 266892
rect 533120 266880 533126 266892
rect 533982 266880 533988 266892
rect 533120 266852 533988 266880
rect 533120 266840 533126 266852
rect 533982 266840 533988 266852
rect 534040 266840 534046 266892
rect 535546 266840 535552 266892
rect 535604 266880 535610 266892
rect 536742 266880 536748 266892
rect 535604 266852 536748 266880
rect 535604 266840 535610 266852
rect 536742 266840 536748 266852
rect 536800 266840 536806 266892
rect 539686 266840 539692 266892
rect 539744 266880 539750 266892
rect 595438 266880 595444 266892
rect 539744 266852 595444 266880
rect 539744 266840 539750 266852
rect 595438 266840 595444 266852
rect 595496 266840 595502 266892
rect 563698 266744 563704 266756
rect 518866 266716 563704 266744
rect 563698 266704 563704 266716
rect 563756 266704 563762 266756
rect 501598 266608 501604 266620
rect 489886 266580 501604 266608
rect 501598 266568 501604 266580
rect 501656 266568 501662 266620
rect 501800 266580 509234 266608
rect 214098 266500 214104 266552
rect 214156 266540 214162 266552
rect 215938 266540 215944 266552
rect 214156 266512 215944 266540
rect 214156 266500 214162 266512
rect 215938 266500 215944 266512
rect 215996 266500 216002 266552
rect 248874 266500 248880 266552
rect 248932 266540 248938 266552
rect 250714 266540 250720 266552
rect 248932 266512 250720 266540
rect 248932 266500 248938 266512
rect 250714 266500 250720 266512
rect 250772 266500 250778 266552
rect 310330 266500 310336 266552
rect 310388 266540 310394 266552
rect 311894 266540 311900 266552
rect 310388 266512 311900 266540
rect 310388 266500 310394 266512
rect 311894 266500 311900 266512
rect 311952 266500 311958 266552
rect 312262 266500 312268 266552
rect 312320 266540 312326 266552
rect 314654 266540 314660 266552
rect 312320 266512 314660 266540
rect 312320 266500 312326 266512
rect 314654 266500 314660 266512
rect 314712 266500 314718 266552
rect 316126 266500 316132 266552
rect 316184 266540 316190 266552
rect 320174 266540 320180 266552
rect 316184 266512 320180 266540
rect 316184 266500 316190 266512
rect 320174 266500 320180 266512
rect 320232 266500 320238 266552
rect 347406 266500 347412 266552
rect 347464 266540 347470 266552
rect 349798 266540 349804 266552
rect 347464 266512 349804 266540
rect 347464 266500 347470 266512
rect 349798 266500 349804 266512
rect 349856 266500 349862 266552
rect 350902 266500 350908 266552
rect 350960 266540 350966 266552
rect 352558 266540 352564 266552
rect 350960 266512 352564 266540
rect 350960 266500 350966 266512
rect 352558 266500 352564 266512
rect 352616 266500 352622 266552
rect 357526 266500 357532 266552
rect 357584 266540 357590 266552
rect 359826 266540 359832 266552
rect 357584 266512 359832 266540
rect 357584 266500 357590 266512
rect 359826 266500 359832 266512
rect 359884 266500 359890 266552
rect 366358 266540 366364 266552
rect 360304 266512 366364 266540
rect 144914 266432 144920 266484
rect 144972 266472 144978 266484
rect 153838 266472 153844 266484
rect 144972 266444 153844 266472
rect 144972 266432 144978 266444
rect 153838 266432 153844 266444
rect 153896 266432 153902 266484
rect 162118 266364 162124 266416
rect 162176 266404 162182 266416
rect 167086 266404 167092 266416
rect 162176 266376 167092 266404
rect 162176 266364 162182 266376
rect 167086 266364 167092 266376
rect 167144 266364 167150 266416
rect 178678 266364 178684 266416
rect 178736 266404 178742 266416
rect 179506 266404 179512 266416
rect 178736 266376 179512 266404
rect 178736 266364 178742 266376
rect 179506 266364 179512 266376
rect 179564 266364 179570 266416
rect 215294 266364 215300 266416
rect 215352 266404 215358 266416
rect 217594 266404 217600 266416
rect 215352 266376 217600 266404
rect 215352 266364 215358 266376
rect 217594 266364 217600 266376
rect 217652 266364 217658 266416
rect 219434 266364 219440 266416
rect 219492 266404 219498 266416
rect 222562 266404 222568 266416
rect 219492 266376 222568 266404
rect 219492 266364 219498 266376
rect 222562 266364 222568 266376
rect 222620 266364 222626 266416
rect 224218 266364 224224 266416
rect 224276 266404 224282 266416
rect 226702 266404 226708 266416
rect 224276 266376 226708 266404
rect 224276 266364 224282 266376
rect 226702 266364 226708 266376
rect 226760 266364 226766 266416
rect 233878 266364 233884 266416
rect 233936 266404 233942 266416
rect 236638 266404 236644 266416
rect 233936 266376 236644 266404
rect 233936 266364 233942 266376
rect 236638 266364 236644 266376
rect 236696 266364 236702 266416
rect 239582 266364 239588 266416
rect 239640 266404 239646 266416
rect 246574 266404 246580 266416
rect 239640 266376 246580 266404
rect 239640 266364 239646 266376
rect 246574 266364 246580 266376
rect 246632 266364 246638 266416
rect 250438 266364 250444 266416
rect 250496 266404 250502 266416
rect 251542 266404 251548 266416
rect 250496 266376 251548 266404
rect 250496 266364 250502 266376
rect 251542 266364 251548 266376
rect 251600 266364 251606 266416
rect 253382 266364 253388 266416
rect 253440 266404 253446 266416
rect 256510 266404 256516 266416
rect 253440 266376 256516 266404
rect 253440 266364 253446 266376
rect 256510 266364 256516 266376
rect 256568 266364 256574 266416
rect 287698 266364 287704 266416
rect 287756 266404 287762 266416
rect 288802 266404 288808 266416
rect 287756 266376 288808 266404
rect 287756 266364 287762 266376
rect 288802 266364 288808 266376
rect 288860 266364 288866 266416
rect 301038 266364 301044 266416
rect 301096 266404 301102 266416
rect 302050 266404 302056 266416
rect 301096 266376 302056 266404
rect 301096 266364 301102 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304534 266404 304540 266416
rect 303764 266376 304540 266404
rect 303764 266364 303770 266376
rect 304534 266364 304540 266376
rect 304592 266364 304598 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309134 266404 309140 266416
rect 307904 266376 309140 266404
rect 307904 266364 307910 266376
rect 309134 266364 309140 266376
rect 309192 266364 309198 266416
rect 309502 266364 309508 266416
rect 309560 266404 309566 266416
rect 310974 266404 310980 266416
rect 309560 266376 310980 266404
rect 309560 266364 309566 266376
rect 310974 266364 310980 266376
rect 311032 266364 311038 266416
rect 311158 266364 311164 266416
rect 311216 266404 311222 266416
rect 313274 266404 313280 266416
rect 311216 266376 313280 266404
rect 311216 266364 311222 266376
rect 313274 266364 313280 266376
rect 313332 266364 313338 266416
rect 320266 266364 320272 266416
rect 320324 266404 320330 266416
rect 321370 266404 321376 266416
rect 320324 266376 321376 266404
rect 320324 266364 320330 266376
rect 321370 266364 321376 266376
rect 321428 266364 321434 266416
rect 324406 266364 324412 266416
rect 324464 266404 324470 266416
rect 325326 266404 325332 266416
rect 324464 266376 325332 266404
rect 324464 266364 324470 266376
rect 325326 266364 325332 266376
rect 325384 266364 325390 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329466 266404 329472 266416
rect 328604 266376 329472 266404
rect 328604 266364 328610 266376
rect 329466 266364 329472 266376
rect 329524 266364 329530 266416
rect 330202 266364 330208 266416
rect 330260 266404 330266 266416
rect 331950 266404 331956 266416
rect 330260 266376 331956 266404
rect 330260 266364 330266 266376
rect 331950 266364 331956 266376
rect 332008 266364 332014 266416
rect 334342 266364 334348 266416
rect 334400 266404 334406 266416
rect 335262 266404 335268 266416
rect 334400 266376 335268 266404
rect 334400 266364 334406 266376
rect 335262 266364 335268 266376
rect 335320 266364 335326 266416
rect 346762 266364 346768 266416
rect 346820 266404 346826 266416
rect 347590 266404 347596 266416
rect 346820 266376 347596 266404
rect 346820 266364 346826 266376
rect 347590 266364 347596 266376
rect 347648 266364 347654 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350350 266404 350356 266416
rect 349304 266376 350356 266404
rect 349304 266364 349310 266376
rect 350350 266364 350356 266376
rect 350408 266364 350414 266416
rect 352558 266364 352564 266416
rect 352616 266404 352622 266416
rect 353938 266404 353944 266416
rect 352616 266376 353944 266404
rect 352616 266364 352622 266376
rect 353938 266364 353944 266376
rect 353996 266364 354002 266416
rect 359182 266364 359188 266416
rect 359240 266404 359246 266416
rect 360102 266404 360108 266416
rect 359240 266376 360108 266404
rect 359240 266364 359246 266376
rect 360102 266364 360108 266376
rect 360160 266364 360166 266416
rect 360010 266228 360016 266280
rect 360068 266268 360074 266280
rect 360304 266268 360332 266512
rect 366358 266500 366364 266512
rect 366416 266500 366422 266552
rect 374914 266500 374920 266552
rect 374972 266540 374978 266552
rect 379698 266540 379704 266552
rect 374972 266512 379704 266540
rect 374972 266500 374978 266512
rect 379698 266500 379704 266512
rect 379756 266500 379762 266552
rect 482554 266500 482560 266552
rect 482612 266540 482618 266552
rect 485038 266540 485044 266552
rect 482612 266512 485044 266540
rect 482612 266500 482618 266512
rect 485038 266500 485044 266512
rect 485096 266500 485102 266552
rect 491662 266432 491668 266484
rect 491720 266472 491726 266484
rect 492582 266472 492588 266484
rect 491720 266444 492588 266472
rect 491720 266432 491726 266444
rect 492582 266432 492588 266444
rect 492640 266432 492646 266484
rect 494146 266432 494152 266484
rect 494204 266472 494210 266484
rect 495250 266472 495256 266484
rect 494204 266444 495256 266472
rect 494204 266432 494210 266444
rect 495250 266432 495256 266444
rect 495308 266432 495314 266484
rect 499942 266432 499948 266484
rect 500000 266472 500006 266484
rect 501800 266472 501828 266580
rect 500000 266444 501828 266472
rect 500000 266432 500006 266444
rect 502426 266432 502432 266484
rect 502484 266472 502490 266484
rect 503438 266472 503444 266484
rect 502484 266444 503444 266472
rect 502484 266432 502490 266444
rect 503438 266432 503444 266444
rect 503496 266432 503502 266484
rect 504082 266432 504088 266484
rect 504140 266472 504146 266484
rect 505002 266472 505008 266484
rect 504140 266444 505008 266472
rect 504140 266432 504146 266444
rect 505002 266432 505008 266444
rect 505060 266432 505066 266484
rect 506566 266432 506572 266484
rect 506624 266472 506630 266484
rect 507670 266472 507676 266484
rect 506624 266444 507676 266472
rect 506624 266432 506630 266444
rect 507670 266432 507676 266444
rect 507728 266432 507734 266484
rect 509206 266472 509234 266580
rect 510706 266568 510712 266620
rect 510764 266608 510770 266620
rect 511810 266608 511816 266620
rect 510764 266580 511816 266608
rect 510764 266568 510770 266580
rect 511810 266568 511816 266580
rect 511868 266568 511874 266620
rect 513926 266568 513932 266620
rect 513984 266608 513990 266620
rect 556798 266608 556804 266620
rect 513984 266580 556804 266608
rect 513984 266568 513990 266580
rect 556798 266568 556804 266580
rect 556856 266568 556862 266620
rect 549898 266472 549904 266484
rect 509206 266444 549904 266472
rect 549898 266432 549904 266444
rect 549956 266432 549962 266484
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362770 266404 362776 266416
rect 361724 266376 362776 266404
rect 361724 266364 361730 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 368290 266364 368296 266416
rect 368348 266404 368354 266416
rect 369118 266404 369124 266416
rect 368348 266376 369124 266404
rect 368348 266364 368354 266376
rect 369118 266364 369124 266376
rect 369176 266364 369182 266416
rect 369394 266364 369400 266416
rect 369452 266404 369458 266416
rect 369854 266404 369860 266416
rect 369452 266376 369860 266404
rect 369452 266364 369458 266376
rect 369854 266364 369860 266376
rect 369912 266364 369918 266416
rect 370314 266364 370320 266416
rect 370372 266404 370378 266416
rect 372154 266404 372160 266416
rect 370372 266376 372160 266404
rect 370372 266364 370378 266376
rect 372154 266364 372160 266376
rect 372212 266364 372218 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375190 266404 375196 266416
rect 374144 266376 375196 266404
rect 374144 266364 374150 266376
rect 375190 266364 375196 266376
rect 375248 266364 375254 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 381538 266404 381544 266416
rect 379940 266376 381544 266404
rect 379940 266364 379946 266376
rect 381538 266364 381544 266376
rect 381596 266364 381602 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387426 266404 387432 266416
rect 386564 266376 387432 266404
rect 386564 266364 386570 266376
rect 387426 266364 387432 266376
rect 387484 266364 387490 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400030 266404 400036 266416
rect 398984 266376 400036 266404
rect 398984 266364 398990 266376
rect 400030 266364 400036 266376
rect 400088 266364 400094 266416
rect 403250 266404 403256 266416
rect 400232 266376 403256 266404
rect 360068 266240 360332 266268
rect 360068 266228 360074 266240
rect 400030 266228 400036 266280
rect 400088 266268 400094 266280
rect 400232 266268 400260 266376
rect 403250 266364 403256 266376
rect 403308 266364 403314 266416
rect 407206 266364 407212 266416
rect 407264 266404 407270 266416
rect 408218 266404 408224 266416
rect 407264 266376 408224 266404
rect 407264 266364 407270 266376
rect 408218 266364 408224 266376
rect 408276 266364 408282 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 427078 266404 427084 266416
rect 425480 266376 427084 266404
rect 425480 266364 425486 266376
rect 427078 266364 427084 266376
rect 427136 266364 427142 266416
rect 429562 266364 429568 266416
rect 429620 266404 429626 266416
rect 430390 266404 430396 266416
rect 429620 266376 430396 266404
rect 429620 266364 429626 266376
rect 430390 266364 430396 266376
rect 430448 266364 430454 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 446122 266364 446128 266416
rect 446180 266404 446186 266416
rect 447778 266404 447784 266416
rect 446180 266376 447784 266404
rect 446180 266364 446186 266376
rect 447778 266364 447784 266376
rect 447836 266364 447842 266416
rect 454402 266364 454408 266416
rect 454460 266404 454466 266416
rect 455230 266404 455236 266416
rect 454460 266376 455236 266404
rect 454460 266364 454466 266376
rect 455230 266364 455236 266376
rect 455288 266364 455294 266416
rect 456886 266364 456892 266416
rect 456944 266404 456950 266416
rect 458082 266404 458088 266416
rect 456944 266376 458088 266404
rect 456944 266364 456950 266376
rect 458082 266364 458088 266376
rect 458140 266364 458146 266416
rect 466822 266364 466828 266416
rect 466880 266404 466886 266416
rect 467742 266404 467748 266416
rect 466880 266376 467748 266404
rect 466880 266364 466886 266376
rect 467742 266364 467748 266376
rect 467800 266364 467806 266416
rect 473446 266364 473452 266416
rect 473504 266404 473510 266416
rect 474642 266404 474648 266416
rect 473504 266376 474648 266404
rect 473504 266364 473510 266376
rect 474642 266364 474648 266376
rect 474700 266364 474706 266416
rect 477586 266364 477592 266416
rect 477644 266404 477650 266416
rect 478506 266404 478512 266416
rect 477644 266376 478512 266404
rect 477644 266364 477650 266376
rect 478506 266364 478512 266376
rect 478564 266364 478570 266416
rect 481726 266364 481732 266416
rect 481784 266404 481790 266416
rect 482830 266404 482836 266416
rect 481784 266376 482836 266404
rect 481784 266364 481790 266376
rect 482830 266364 482836 266376
rect 482888 266364 482894 266416
rect 483382 266364 483388 266416
rect 483440 266404 483446 266416
rect 484302 266404 484308 266416
rect 483440 266376 484308 266404
rect 483440 266364 483446 266376
rect 484302 266364 484308 266376
rect 484360 266364 484366 266416
rect 485866 266364 485872 266416
rect 485924 266404 485930 266416
rect 487062 266404 487068 266416
rect 485924 266376 487068 266404
rect 485924 266364 485930 266376
rect 487062 266364 487068 266376
rect 487120 266364 487126 266416
rect 560478 266336 560484 266348
rect 487264 266308 560484 266336
rect 400088 266240 400260 266268
rect 400088 266228 400094 266240
rect 484210 266228 484216 266280
rect 484268 266268 484274 266280
rect 487264 266268 487292 266308
rect 560478 266296 560484 266308
rect 560536 266296 560542 266348
rect 484268 266240 487292 266268
rect 484268 266228 484274 266240
rect 487522 266160 487528 266212
rect 487580 266200 487586 266212
rect 565814 266200 565820 266212
rect 487580 266172 565820 266200
rect 487580 266160 487586 266172
rect 565814 266160 565820 266172
rect 565872 266160 565878 266212
rect 492490 266024 492496 266076
rect 492548 266064 492554 266076
rect 572714 266064 572720 266076
rect 492548 266036 572720 266064
rect 492548 266024 492554 266036
rect 572714 266024 572720 266036
rect 572772 266024 572778 266076
rect 512362 265888 512368 265940
rect 512420 265928 512426 265940
rect 600314 265928 600320 265940
rect 512420 265900 600320 265928
rect 512420 265888 512426 265900
rect 600314 265888 600320 265900
rect 600372 265888 600378 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 151998 265616 152004 265668
rect 152056 265656 152062 265668
rect 152734 265656 152740 265668
rect 152056 265628 152740 265656
rect 152056 265616 152062 265628
rect 152734 265616 152740 265628
rect 152792 265616 152798 265668
rect 155954 265616 155960 265668
rect 156012 265656 156018 265668
rect 156782 265656 156788 265668
rect 156012 265628 156788 265656
rect 156012 265616 156018 265628
rect 156782 265616 156788 265628
rect 156840 265616 156846 265668
rect 172514 265616 172520 265668
rect 172572 265656 172578 265668
rect 173342 265656 173348 265668
rect 172572 265628 173348 265656
rect 172572 265616 172578 265628
rect 173342 265616 173348 265628
rect 173400 265616 173406 265668
rect 189166 265616 189172 265668
rect 189224 265656 189230 265668
rect 189902 265656 189908 265668
rect 189224 265628 189908 265656
rect 189224 265616 189230 265628
rect 189902 265616 189908 265628
rect 189960 265616 189966 265668
rect 229094 265616 229100 265668
rect 229152 265656 229158 265668
rect 229646 265656 229652 265668
rect 229152 265628 229652 265656
rect 229152 265616 229158 265628
rect 229646 265616 229652 265628
rect 229704 265616 229710 265668
rect 243078 265616 243084 265668
rect 243136 265656 243142 265668
rect 243814 265656 243820 265668
rect 243136 265628 243820 265656
rect 243136 265616 243142 265628
rect 243814 265616 243820 265628
rect 243872 265616 243878 265668
rect 253934 265616 253940 265668
rect 253992 265656 253998 265668
rect 254486 265656 254492 265668
rect 253992 265628 254492 265656
rect 253992 265616 253998 265628
rect 254486 265616 254492 265628
rect 254544 265616 254550 265668
rect 280338 265616 280344 265668
rect 280396 265656 280402 265668
rect 280982 265656 280988 265668
rect 280396 265628 280988 265656
rect 280396 265616 280402 265628
rect 280982 265616 280988 265628
rect 281040 265616 281046 265668
rect 284294 265616 284300 265668
rect 284352 265656 284358 265668
rect 285214 265656 285220 265668
rect 284352 265628 285220 265656
rect 284352 265616 284358 265628
rect 285214 265616 285220 265628
rect 285272 265616 285278 265668
rect 296806 265616 296812 265668
rect 296864 265656 296870 265668
rect 297542 265656 297548 265668
rect 296864 265628 297548 265656
rect 296864 265616 296870 265628
rect 297542 265616 297548 265628
rect 297600 265616 297606 265668
rect 520642 265616 520648 265668
rect 520700 265656 520706 265668
rect 612734 265656 612740 265668
rect 520700 265628 612740 265656
rect 520700 265616 520706 265628
rect 612734 265616 612740 265628
rect 612792 265616 612798 265668
rect 480070 265480 480076 265532
rect 480128 265520 480134 265532
rect 554774 265520 554780 265532
rect 480128 265492 554780 265520
rect 480128 265480 480134 265492
rect 554774 265480 554780 265492
rect 554832 265480 554838 265532
rect 479242 265344 479248 265396
rect 479300 265384 479306 265396
rect 553394 265384 553400 265396
rect 479300 265356 553400 265384
rect 479300 265344 479306 265356
rect 553394 265344 553400 265356
rect 553452 265344 553458 265396
rect 475102 265208 475108 265260
rect 475160 265248 475166 265260
rect 547966 265248 547972 265260
rect 475160 265220 547972 265248
rect 475160 265208 475166 265220
rect 547966 265208 547972 265220
rect 548024 265208 548030 265260
rect 469306 265072 469312 265124
rect 469364 265112 469370 265124
rect 539962 265112 539968 265124
rect 469364 265084 539968 265112
rect 469364 265072 469370 265084
rect 539962 265072 539968 265084
rect 540020 265072 540026 265124
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 676030 259564 676036 259616
rect 676088 259604 676094 259616
rect 676214 259604 676220 259616
rect 676088 259576 676220 259604
rect 676088 259564 676094 259576
rect 676214 259564 676220 259576
rect 676272 259564 676278 259616
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 560938 259468 560944 259480
rect 554372 259440 560944 259468
rect 554372 259428 554378 259440
rect 560938 259428 560944 259440
rect 560996 259428 561002 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 563698 256748 563704 256760
rect 554004 256720 563704 256748
rect 554004 256708 554010 256720
rect 563698 256708 563704 256720
rect 563756 256708 563762 256760
rect 553486 255552 553492 255604
rect 553544 255592 553550 255604
rect 555418 255592 555424 255604
rect 553544 255564 555424 255592
rect 553544 255552 553550 255564
rect 555418 255552 555424 255564
rect 555476 255552 555482 255604
rect 35802 255416 35808 255468
rect 35860 255456 35866 255468
rect 39758 255456 39764 255468
rect 35860 255428 39764 255456
rect 35860 255416 35866 255428
rect 39758 255416 39764 255428
rect 39816 255416 39822 255468
rect 675846 254600 675852 254652
rect 675904 254640 675910 254652
rect 683022 254640 683028 254652
rect 675904 254612 683028 254640
rect 675904 254600 675910 254612
rect 683022 254600 683028 254612
rect 683080 254600 683086 254652
rect 675018 254260 675024 254312
rect 675076 254300 675082 254312
rect 675478 254300 675484 254312
rect 675076 254272 675484 254300
rect 675076 254260 675082 254272
rect 675478 254260 675484 254272
rect 675536 254260 675542 254312
rect 35802 254056 35808 254108
rect 35860 254096 35866 254108
rect 39574 254096 39580 254108
rect 35860 254068 39580 254096
rect 35860 254056 35866 254068
rect 39574 254056 39580 254068
rect 39632 254056 39638 254108
rect 35802 252696 35808 252748
rect 35860 252736 35866 252748
rect 41690 252736 41696 252748
rect 35860 252708 41696 252736
rect 35860 252696 35866 252708
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 35618 252560 35624 252612
rect 35676 252600 35682 252612
rect 40954 252600 40960 252612
rect 35676 252572 40960 252600
rect 35676 252560 35682 252572
rect 40954 252560 40960 252572
rect 41012 252560 41018 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 35802 251336 35808 251388
rect 35860 251376 35866 251388
rect 40494 251376 40500 251388
rect 35860 251348 40500 251376
rect 35860 251336 35866 251348
rect 40494 251336 40500 251348
rect 40552 251336 40558 251388
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 35802 249908 35808 249960
rect 35860 249948 35866 249960
rect 39390 249948 39396 249960
rect 35860 249920 39396 249948
rect 35860 249908 35866 249920
rect 39390 249908 39396 249920
rect 39448 249908 39454 249960
rect 35802 248480 35808 248532
rect 35860 248520 35866 248532
rect 39206 248520 39212 248532
rect 35860 248492 39212 248520
rect 35860 248480 35866 248492
rect 39206 248480 39212 248492
rect 39264 248480 39270 248532
rect 35802 247188 35808 247240
rect 35860 247228 35866 247240
rect 41690 247228 41696 247240
rect 35860 247200 41696 247228
rect 35860 247188 35866 247200
rect 41690 247188 41696 247200
rect 41748 247188 41754 247240
rect 35618 247052 35624 247104
rect 35676 247092 35682 247104
rect 41506 247092 41512 247104
rect 35676 247064 41512 247092
rect 35676 247052 35682 247064
rect 41506 247052 41512 247064
rect 41564 247052 41570 247104
rect 558178 246304 558184 246356
rect 558236 246344 558242 246356
rect 647234 246344 647240 246356
rect 558236 246316 647240 246344
rect 558236 246304 558242 246316
rect 647234 246304 647240 246316
rect 647292 246304 647298 246356
rect 553854 245624 553860 245676
rect 553912 245664 553918 245676
rect 596818 245664 596824 245676
rect 553912 245636 596824 245664
rect 553912 245624 553918 245636
rect 596818 245624 596824 245636
rect 596876 245624 596882 245676
rect 554498 244264 554504 244316
rect 554556 244304 554562 244316
rect 573358 244304 573364 244316
rect 554556 244276 573364 244304
rect 554556 244264 554562 244276
rect 573358 244264 573364 244276
rect 573416 244264 573422 244316
rect 674742 242700 674748 242752
rect 674800 242740 674806 242752
rect 675294 242740 675300 242752
rect 674800 242712 675300 242740
rect 674800 242700 674806 242712
rect 675294 242700 675300 242712
rect 675352 242700 675358 242752
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553670 241476 553676 241528
rect 553728 241516 553734 241528
rect 629938 241516 629944 241528
rect 553728 241488 629944 241516
rect 553728 241476 553734 241488
rect 629938 241476 629944 241488
rect 629996 241476 630002 241528
rect 554498 240116 554504 240168
rect 554556 240156 554562 240168
rect 577498 240156 577504 240168
rect 554556 240128 577504 240156
rect 554556 240116 554562 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 668762 236988 668768 237040
rect 668820 237028 668826 237040
rect 671522 237028 671528 237040
rect 668820 237000 671528 237028
rect 668820 236988 668826 237000
rect 671522 236988 671528 237000
rect 671580 236988 671586 237040
rect 672756 236892 672784 237082
rect 672736 236864 672784 236892
rect 672074 236784 672080 236836
rect 672132 236824 672138 236836
rect 672736 236824 672764 236864
rect 672132 236796 672764 236824
rect 672132 236784 672138 236796
rect 672874 236756 672902 236878
rect 672828 236728 672902 236756
rect 671522 236580 671528 236632
rect 671580 236620 671586 236632
rect 672828 236620 672856 236728
rect 672954 236700 673006 236706
rect 672954 236642 673006 236648
rect 671580 236592 672856 236620
rect 671580 236580 671586 236592
rect 671706 236444 671712 236496
rect 671764 236484 671770 236496
rect 671764 236456 673118 236484
rect 671764 236444 671770 236456
rect 673184 236292 673236 236298
rect 673184 236234 673236 236240
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 672184 236048 673330 236076
rect 670970 235900 670976 235952
rect 671028 235940 671034 235952
rect 672184 235940 672212 236048
rect 671028 235912 672212 235940
rect 671028 235900 671034 235912
rect 673270 235900 673276 235952
rect 673328 235940 673334 235952
rect 673328 235912 673440 235940
rect 673328 235900 673334 235912
rect 670142 235764 670148 235816
rect 670200 235804 670206 235816
rect 672074 235804 672080 235816
rect 670200 235776 672080 235804
rect 670200 235764 670206 235776
rect 672074 235764 672080 235776
rect 672132 235764 672138 235816
rect 672626 235696 672632 235748
rect 672684 235736 672690 235748
rect 672684 235708 673554 235736
rect 672684 235696 672690 235708
rect 673086 235492 673092 235544
rect 673144 235532 673150 235544
rect 673144 235504 673670 235532
rect 673144 235492 673150 235504
rect 669590 235288 669596 235340
rect 669648 235328 669654 235340
rect 669648 235300 673778 235328
rect 669648 235288 669654 235300
rect 668210 235084 668216 235136
rect 668268 235124 668274 235136
rect 668268 235096 673900 235124
rect 668268 235084 668274 235096
rect 668394 234812 668400 234864
rect 668452 234852 668458 234864
rect 673978 234852 674006 234906
rect 668452 234824 674006 234852
rect 668452 234812 668458 234824
rect 674088 234728 674140 234734
rect 674088 234670 674140 234676
rect 661678 234608 661684 234660
rect 661736 234648 661742 234660
rect 670418 234648 670424 234660
rect 661736 234620 670424 234648
rect 661736 234608 661742 234620
rect 670418 234608 670424 234620
rect 670476 234608 670482 234660
rect 42426 234540 42432 234592
rect 42484 234580 42490 234592
rect 42978 234580 42984 234592
rect 42484 234552 42984 234580
rect 42484 234540 42490 234552
rect 42978 234540 42984 234552
rect 43036 234540 43042 234592
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 669406 234472 669412 234524
rect 669464 234512 669470 234524
rect 669464 234484 674222 234512
rect 669464 234472 669470 234484
rect 675110 234472 675116 234524
rect 675168 234472 675174 234524
rect 671890 234336 671896 234388
rect 671948 234376 671954 234388
rect 675128 234376 675156 234472
rect 671948 234348 675156 234376
rect 671948 234336 671954 234348
rect 671154 234200 671160 234252
rect 671212 234240 671218 234252
rect 674098 234240 674104 234252
rect 671212 234212 674104 234240
rect 671212 234200 671218 234212
rect 674098 234200 674104 234212
rect 674156 234200 674162 234252
rect 675846 233928 675852 233980
rect 675904 233968 675910 233980
rect 683390 233968 683396 233980
rect 675904 233940 683396 233968
rect 675904 233928 675910 233940
rect 683390 233928 683396 233940
rect 683448 233928 683454 233980
rect 652386 233860 652392 233912
rect 652444 233900 652450 233912
rect 652444 233872 663794 233900
rect 652444 233860 652450 233872
rect 663766 233764 663794 233872
rect 674098 233832 674104 233844
rect 666526 233804 674104 233832
rect 666526 233764 666554 233804
rect 674098 233792 674104 233804
rect 674156 233792 674162 233844
rect 676030 233792 676036 233844
rect 676088 233832 676094 233844
rect 678238 233832 678244 233844
rect 676088 233804 678244 233832
rect 676088 233792 676094 233804
rect 678238 233792 678244 233804
rect 678296 233792 678302 233844
rect 663766 233736 666554 233764
rect 670326 233180 670332 233232
rect 670384 233220 670390 233232
rect 672626 233220 672632 233232
rect 670384 233192 672632 233220
rect 670384 233180 670390 233192
rect 672626 233180 672632 233192
rect 672684 233180 672690 233232
rect 639598 232500 639604 232552
rect 639656 232540 639662 232552
rect 654778 232540 654784 232552
rect 639656 232512 654784 232540
rect 639656 232500 639662 232512
rect 654778 232500 654784 232512
rect 654836 232500 654842 232552
rect 660298 232500 660304 232552
rect 660356 232540 660362 232552
rect 660356 232512 663794 232540
rect 660356 232500 660362 232512
rect 663766 232472 663794 232512
rect 675846 232500 675852 232552
rect 675904 232540 675910 232552
rect 683206 232540 683212 232552
rect 675904 232512 683212 232540
rect 675904 232500 675910 232512
rect 683206 232500 683212 232512
rect 683264 232500 683270 232552
rect 671890 232472 671896 232484
rect 663766 232444 671896 232472
rect 671890 232432 671896 232444
rect 671948 232432 671954 232484
rect 665450 231616 665456 231668
rect 665508 231656 665514 231668
rect 674926 231656 674932 231668
rect 665508 231628 674932 231656
rect 665508 231616 665514 231628
rect 674926 231616 674932 231628
rect 674984 231616 674990 231668
rect 146202 231548 146208 231600
rect 146260 231588 146266 231600
rect 150526 231588 150532 231600
rect 146260 231560 150532 231588
rect 146260 231548 146266 231560
rect 150526 231548 150532 231560
rect 150584 231548 150590 231600
rect 663058 231480 663064 231532
rect 663116 231520 663122 231532
rect 671890 231520 671896 231532
rect 663116 231492 671896 231520
rect 663116 231480 663122 231492
rect 671890 231480 671896 231492
rect 671948 231480 671954 231532
rect 675846 231480 675852 231532
rect 675904 231520 675910 231532
rect 683574 231520 683580 231532
rect 675904 231492 683580 231520
rect 675904 231480 675910 231492
rect 683574 231480 683580 231492
rect 683632 231480 683638 231532
rect 146754 231412 146760 231464
rect 146812 231452 146818 231464
rect 147214 231452 147220 231464
rect 146812 231424 147220 231452
rect 146812 231412 146818 231424
rect 147214 231412 147220 231424
rect 147272 231412 147278 231464
rect 662322 231344 662328 231396
rect 662380 231384 662386 231396
rect 675110 231384 675116 231396
rect 662380 231356 675116 231384
rect 662380 231344 662386 231356
rect 675110 231344 675116 231356
rect 675168 231344 675174 231396
rect 137922 231276 137928 231328
rect 137980 231316 137986 231328
rect 152458 231316 152464 231328
rect 137980 231288 152464 231316
rect 137980 231276 137986 231288
rect 152458 231276 152464 231288
rect 152516 231276 152522 231328
rect 156506 231276 156512 231328
rect 156564 231316 156570 231328
rect 163682 231316 163688 231328
rect 156564 231288 163688 231316
rect 156564 231276 156570 231288
rect 163682 231276 163688 231288
rect 163740 231276 163746 231328
rect 91738 231140 91744 231192
rect 91796 231180 91802 231192
rect 168834 231180 168840 231192
rect 91796 231152 168840 231180
rect 91796 231140 91802 231152
rect 168834 231140 168840 231152
rect 168892 231140 168898 231192
rect 664990 231140 664996 231192
rect 665048 231180 665054 231192
rect 665048 231152 675326 231180
rect 665048 231140 665054 231152
rect 596818 231072 596824 231124
rect 596876 231112 596882 231124
rect 633618 231112 633624 231124
rect 596876 231084 633624 231112
rect 596876 231072 596882 231084
rect 633618 231072 633624 231084
rect 633676 231072 633682 231124
rect 636838 231072 636844 231124
rect 636896 231112 636902 231124
rect 650638 231112 650644 231124
rect 636896 231084 650644 231112
rect 636896 231072 636902 231084
rect 650638 231072 650644 231084
rect 650696 231072 650702 231124
rect 675116 231056 675168 231062
rect 128262 231004 128268 231056
rect 128320 231044 128326 231056
rect 195882 231044 195888 231056
rect 128320 231016 195888 231044
rect 128320 231004 128326 231016
rect 195882 231004 195888 231016
rect 195940 231004 195946 231056
rect 675116 230998 675168 231004
rect 118602 230868 118608 230920
rect 118660 230908 118666 230920
rect 188154 230908 188160 230920
rect 118660 230880 188160 230908
rect 118660 230868 118666 230880
rect 188154 230868 188160 230880
rect 188212 230868 188218 230920
rect 674956 230852 675008 230858
rect 674956 230794 675008 230800
rect 110322 230732 110328 230784
rect 110380 230772 110386 230784
rect 184290 230772 184296 230784
rect 110380 230744 184296 230772
rect 110380 230732 110386 230744
rect 184290 230732 184296 230744
rect 184348 230732 184354 230784
rect 97902 230596 97908 230648
rect 97960 230636 97966 230648
rect 173986 230636 173992 230648
rect 97960 230608 173992 230636
rect 97960 230596 97966 230608
rect 173986 230596 173992 230608
rect 174044 230596 174050 230648
rect 195054 230596 195060 230648
rect 195112 230636 195118 230648
rect 196894 230636 196900 230648
rect 195112 230608 196900 230636
rect 195112 230596 195118 230608
rect 196894 230596 196900 230608
rect 196952 230596 196958 230648
rect 672074 230596 672080 230648
rect 672132 230636 672138 230648
rect 672132 230608 674820 230636
rect 672132 230596 672138 230608
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 152458 230460 152464 230512
rect 152516 230500 152522 230512
rect 203610 230500 203616 230512
rect 152516 230472 203616 230500
rect 152516 230460 152522 230472
rect 203610 230460 203616 230472
rect 203668 230460 203674 230512
rect 42426 230392 42432 230444
rect 42484 230432 42490 230444
rect 43070 230432 43076 230444
rect 42484 230404 43076 230432
rect 42484 230392 42490 230404
rect 43070 230392 43076 230404
rect 43128 230392 43134 230444
rect 130378 230392 130384 230444
rect 130436 230432 130442 230444
rect 142430 230432 142436 230444
rect 130436 230404 142436 230432
rect 130436 230392 130442 230404
rect 142430 230392 142436 230404
rect 142488 230392 142494 230444
rect 142614 230392 142620 230444
rect 142672 230432 142678 230444
rect 146202 230432 146208 230444
rect 142672 230404 146208 230432
rect 142672 230392 142678 230404
rect 146202 230392 146208 230404
rect 146260 230392 146266 230444
rect 147628 230392 147634 230444
rect 147686 230432 147692 230444
rect 149514 230432 149520 230444
rect 147686 230404 149520 230432
rect 147686 230392 147692 230404
rect 149514 230392 149520 230404
rect 149572 230392 149578 230444
rect 206278 230392 206284 230444
rect 206336 230432 206342 230444
rect 256418 230432 256424 230444
rect 206336 230404 256424 230432
rect 206336 230392 206342 230404
rect 256418 230392 256424 230404
rect 256476 230392 256482 230444
rect 276290 230392 276296 230444
rect 276348 230432 276354 230444
rect 292482 230432 292488 230444
rect 276348 230404 292488 230432
rect 276348 230392 276354 230404
rect 292482 230392 292488 230404
rect 292540 230392 292546 230444
rect 308398 230392 308404 230444
rect 308456 230432 308462 230444
rect 334986 230432 334992 230444
rect 308456 230404 334992 230432
rect 308456 230392 308462 230404
rect 334986 230392 334992 230404
rect 335044 230392 335050 230444
rect 439516 230432 439544 230540
rect 674676 230444 674728 230450
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 526898 230392 526904 230444
rect 526956 230432 526962 230444
rect 536098 230432 536104 230444
rect 526956 230404 536104 230432
rect 526956 230392 526962 230404
rect 536098 230392 536104 230404
rect 536156 230392 536162 230444
rect 674676 230386 674728 230392
rect 387426 230324 387432 230376
rect 387484 230364 387490 230376
rect 388438 230364 388444 230376
rect 387484 230336 388444 230364
rect 387484 230324 387490 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 398098 230324 398104 230376
rect 398156 230364 398162 230376
rect 399386 230364 399392 230376
rect 398156 230336 399392 230364
rect 398156 230324 398162 230336
rect 399386 230324 399392 230336
rect 399444 230324 399450 230376
rect 436094 230324 436100 230376
rect 436152 230364 436158 230376
rect 436738 230364 436744 230376
rect 436152 230336 436744 230364
rect 436152 230324 436158 230336
rect 436738 230324 436744 230336
rect 436796 230324 436802 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 443822 230324 443828 230376
rect 443880 230364 443886 230376
rect 444834 230364 444840 230376
rect 443880 230336 444840 230364
rect 443880 230324 443886 230336
rect 444834 230324 444840 230336
rect 444892 230324 444898 230376
rect 446398 230324 446404 230376
rect 446456 230364 446462 230376
rect 448698 230364 448704 230376
rect 446456 230336 448704 230364
rect 446456 230324 446462 230336
rect 448698 230324 448704 230336
rect 448756 230324 448762 230376
rect 449618 230324 449624 230376
rect 449676 230364 449682 230376
rect 450538 230364 450544 230376
rect 449676 230336 450544 230364
rect 449676 230324 449682 230336
rect 450538 230324 450544 230336
rect 450596 230324 450602 230376
rect 452838 230324 452844 230376
rect 452896 230364 452902 230376
rect 454310 230364 454316 230376
rect 452896 230336 454316 230364
rect 452896 230324 452902 230336
rect 454310 230324 454316 230336
rect 454368 230324 454374 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 470870 230324 470876 230376
rect 470928 230364 470934 230376
rect 471882 230364 471888 230376
rect 470928 230336 471888 230364
rect 470928 230324 470934 230336
rect 471882 230324 471888 230336
rect 471940 230324 471946 230376
rect 472158 230324 472164 230376
rect 472216 230364 472222 230376
rect 473170 230364 473176 230376
rect 472216 230336 473176 230364
rect 472216 230324 472222 230336
rect 473170 230324 473176 230336
rect 473228 230324 473234 230376
rect 487614 230324 487620 230376
rect 487672 230364 487678 230376
rect 488442 230364 488448 230376
rect 487672 230336 488448 230364
rect 487672 230324 487678 230336
rect 488442 230324 488448 230336
rect 488500 230324 488506 230376
rect 493410 230324 493416 230376
rect 493468 230364 493474 230376
rect 496354 230364 496360 230376
rect 493468 230336 496360 230364
rect 493468 230324 493474 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 497274 230324 497280 230376
rect 497332 230364 497338 230376
rect 498102 230364 498108 230376
rect 497332 230336 498108 230364
rect 497332 230324 497338 230336
rect 498102 230324 498108 230336
rect 498160 230324 498166 230376
rect 511442 230324 511448 230376
rect 511500 230364 511506 230376
rect 517514 230364 517520 230376
rect 511500 230336 517520 230364
rect 511500 230324 511506 230336
rect 517514 230324 517520 230336
rect 517572 230324 517578 230376
rect 133782 230256 133788 230308
rect 133840 230296 133846 230308
rect 202322 230296 202328 230308
rect 133840 230268 202328 230296
rect 133840 230256 133846 230268
rect 202322 230256 202328 230268
rect 202380 230256 202386 230308
rect 210418 230256 210424 230308
rect 210476 230296 210482 230308
rect 261570 230296 261576 230308
rect 210476 230268 261576 230296
rect 210476 230256 210482 230268
rect 261570 230256 261576 230268
rect 261628 230256 261634 230308
rect 275646 230256 275652 230308
rect 275704 230296 275710 230308
rect 313090 230296 313096 230308
rect 275704 230268 313096 230296
rect 275704 230256 275710 230268
rect 313090 230256 313096 230268
rect 313148 230256 313154 230308
rect 528830 230256 528836 230308
rect 528888 230296 528894 230308
rect 539594 230296 539600 230308
rect 528888 230268 539600 230296
rect 528888 230256 528894 230268
rect 539594 230256 539600 230268
rect 539652 230256 539658 230308
rect 674564 230240 674616 230246
rect 388438 230188 388444 230240
rect 388496 230228 388502 230240
rect 391658 230228 391664 230240
rect 388496 230200 391664 230228
rect 388496 230188 388502 230200
rect 391658 230188 391664 230200
rect 391716 230188 391722 230240
rect 444466 230188 444472 230240
rect 444524 230228 444530 230240
rect 447686 230228 447692 230240
rect 444524 230200 447692 230228
rect 444524 230188 444530 230200
rect 447686 230188 447692 230200
rect 447744 230188 447750 230240
rect 451550 230188 451556 230240
rect 451608 230228 451614 230240
rect 453298 230228 453304 230240
rect 451608 230200 453304 230228
rect 451608 230188 451614 230200
rect 453298 230188 453304 230200
rect 453356 230188 453362 230240
rect 453482 230188 453488 230240
rect 453540 230228 453546 230240
rect 455782 230228 455788 230240
rect 453540 230200 455788 230228
rect 453540 230188 453546 230200
rect 455782 230188 455788 230200
rect 455840 230188 455846 230240
rect 468294 230188 468300 230240
rect 468352 230228 468358 230240
rect 469122 230228 469128 230240
rect 468352 230200 469128 230228
rect 468352 230188 468358 230200
rect 469122 230188 469128 230200
rect 469180 230188 469186 230240
rect 490190 230188 490196 230240
rect 490248 230228 490254 230240
rect 493686 230228 493692 230240
rect 490248 230200 493692 230228
rect 490248 230188 490254 230200
rect 493686 230188 493692 230200
rect 493744 230188 493750 230240
rect 674564 230182 674616 230188
rect 95234 230120 95240 230172
rect 95292 230160 95298 230172
rect 157288 230160 157294 230172
rect 95292 230132 157294 230160
rect 95292 230120 95298 230132
rect 157288 230120 157294 230132
rect 157346 230120 157352 230172
rect 157426 230120 157432 230172
rect 157484 230160 157490 230172
rect 161106 230160 161112 230172
rect 157484 230132 161112 230160
rect 157484 230120 157490 230132
rect 161106 230120 161112 230132
rect 161164 230120 161170 230172
rect 176746 230120 176752 230172
rect 176804 230160 176810 230172
rect 235810 230160 235816 230172
rect 176804 230132 235816 230160
rect 176804 230120 176810 230132
rect 235810 230120 235816 230132
rect 235868 230120 235874 230172
rect 264238 230120 264244 230172
rect 264296 230160 264302 230172
rect 302786 230160 302792 230172
rect 264296 230132 302792 230160
rect 264296 230120 264302 230132
rect 302786 230120 302792 230132
rect 302844 230120 302850 230172
rect 302970 230120 302976 230172
rect 303028 230160 303034 230172
rect 329834 230160 329840 230172
rect 303028 230132 329840 230160
rect 303028 230120 303034 230132
rect 329834 230120 329840 230132
rect 329892 230120 329898 230172
rect 334250 230120 334256 230172
rect 334308 230160 334314 230172
rect 355594 230160 355600 230172
rect 334308 230132 355600 230160
rect 334308 230120 334314 230132
rect 355594 230120 355600 230132
rect 355652 230120 355658 230172
rect 521102 230120 521108 230172
rect 521160 230160 521166 230172
rect 529198 230160 529204 230172
rect 521160 230132 529204 230160
rect 521160 230120 521166 230132
rect 529198 230120 529204 230132
rect 529256 230120 529262 230172
rect 532694 230120 532700 230172
rect 532752 230160 532758 230172
rect 547138 230160 547144 230172
rect 532752 230132 547144 230160
rect 532752 230120 532758 230132
rect 547138 230120 547144 230132
rect 547196 230120 547202 230172
rect 454126 230052 454132 230104
rect 454184 230092 454190 230104
rect 455322 230092 455328 230104
rect 454184 230064 455328 230092
rect 454184 230052 454190 230064
rect 455322 230052 455328 230064
rect 455380 230052 455386 230104
rect 491478 230052 491484 230104
rect 491536 230092 491542 230104
rect 492490 230092 492496 230104
rect 491536 230064 492496 230092
rect 491536 230052 491542 230064
rect 492490 230052 492496 230064
rect 492548 230052 492554 230104
rect 126882 229984 126888 230036
rect 126940 230024 126946 230036
rect 195054 230024 195060 230036
rect 126940 229996 195060 230024
rect 126940 229984 126946 229996
rect 195054 229984 195060 229996
rect 195112 229984 195118 230036
rect 195422 229984 195428 230036
rect 195480 230024 195486 230036
rect 214742 230024 214748 230036
rect 195480 229996 214748 230024
rect 195480 229984 195486 229996
rect 214742 229984 214748 229996
rect 214800 229984 214806 230036
rect 219986 229984 219992 230036
rect 220044 230024 220050 230036
rect 230658 230024 230664 230036
rect 220044 229996 230664 230024
rect 220044 229984 220050 229996
rect 230658 229984 230664 229996
rect 230716 229984 230722 230036
rect 242526 229984 242532 230036
rect 242584 230024 242590 230036
rect 287330 230024 287336 230036
rect 242584 229996 287336 230024
rect 242584 229984 242590 229996
rect 287330 229984 287336 229996
rect 287388 229984 287394 230036
rect 287514 229984 287520 230036
rect 287572 230024 287578 230036
rect 307938 230024 307944 230036
rect 287572 229996 307944 230024
rect 287572 229984 287578 229996
rect 307938 229984 307944 229996
rect 307996 229984 308002 230036
rect 312630 229984 312636 230036
rect 312688 230024 312694 230036
rect 340138 230024 340144 230036
rect 312688 229996 340144 230024
rect 312688 229984 312694 229996
rect 340138 229984 340144 229996
rect 340196 229984 340202 230036
rect 354950 229984 354956 230036
rect 355008 230024 355014 230036
rect 371050 230024 371056 230036
rect 355008 229996 371056 230024
rect 355008 229984 355014 229996
rect 371050 229984 371056 229996
rect 371108 229984 371114 230036
rect 476666 229984 476672 230036
rect 476724 230024 476730 230036
rect 481634 230024 481640 230036
rect 476724 229996 481640 230024
rect 476724 229984 476730 229996
rect 481634 229984 481640 229996
rect 481692 229984 481698 230036
rect 515306 229984 515312 230036
rect 515364 230024 515370 230036
rect 524598 230024 524604 230036
rect 515364 229996 524604 230024
rect 515364 229984 515370 229996
rect 524598 229984 524604 229996
rect 524656 229984 524662 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 549254 230024 549260 230036
rect 534684 229996 549260 230024
rect 534684 229984 534690 229996
rect 549254 229984 549260 229996
rect 549312 229984 549318 230036
rect 674452 229968 674504 229974
rect 674452 229910 674504 229916
rect 86218 229848 86224 229900
rect 86276 229888 86282 229900
rect 156690 229888 156696 229900
rect 86276 229860 156696 229888
rect 86276 229848 86282 229860
rect 156690 229848 156696 229860
rect 156748 229848 156754 229900
rect 158530 229888 158536 229900
rect 157168 229860 158536 229888
rect 68278 229712 68284 229764
rect 68336 229752 68342 229764
rect 142614 229752 142620 229764
rect 68336 229724 142620 229752
rect 68336 229712 68342 229724
rect 142614 229712 142620 229724
rect 142672 229712 142678 229764
rect 147766 229752 147772 229764
rect 147646 229724 147772 229752
rect 147646 229684 147674 229724
rect 147766 229712 147772 229724
rect 147824 229712 147830 229764
rect 157168 229752 157196 229860
rect 158530 229848 158536 229860
rect 158588 229848 158594 229900
rect 163958 229848 163964 229900
rect 164016 229888 164022 229900
rect 225506 229888 225512 229900
rect 164016 229860 225512 229888
rect 164016 229848 164022 229860
rect 225506 229848 225512 229860
rect 225564 229848 225570 229900
rect 230474 229848 230480 229900
rect 230532 229888 230538 229900
rect 277026 229888 277032 229900
rect 230532 229860 277032 229888
rect 230532 229848 230538 229860
rect 277026 229848 277032 229860
rect 277084 229848 277090 229900
rect 282546 229848 282552 229900
rect 282604 229888 282610 229900
rect 318242 229888 318248 229900
rect 282604 229860 318248 229888
rect 282604 229848 282610 229860
rect 318242 229848 318248 229860
rect 318300 229848 318306 229900
rect 324222 229848 324228 229900
rect 324280 229888 324286 229900
rect 350442 229888 350448 229900
rect 324280 229860 350448 229888
rect 324280 229848 324286 229860
rect 350442 229848 350448 229860
rect 350500 229848 350506 229900
rect 366726 229848 366732 229900
rect 366784 229888 366790 229900
rect 383930 229888 383936 229900
rect 366784 229860 383936 229888
rect 366784 229848 366790 229860
rect 383930 229848 383936 229860
rect 383988 229848 383994 229900
rect 457346 229848 457352 229900
rect 457404 229888 457410 229900
rect 464062 229888 464068 229900
rect 457404 229860 464068 229888
rect 457404 229848 457410 229860
rect 464062 229848 464068 229860
rect 464120 229848 464126 229900
rect 469582 229848 469588 229900
rect 469640 229888 469646 229900
rect 469640 229860 474228 229888
rect 469640 229848 469646 229860
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 147968 229724 157196 229752
rect 142816 229656 147674 229684
rect 82078 229576 82084 229628
rect 82136 229616 82142 229628
rect 142816 229616 142844 229656
rect 82136 229588 142844 229616
rect 82136 229576 82142 229588
rect 147122 229508 147128 229560
rect 147180 229548 147186 229560
rect 147968 229548 147996 229724
rect 157288 229712 157294 229764
rect 157346 229752 157352 229764
rect 166258 229752 166264 229764
rect 157346 229724 166264 229752
rect 157346 229712 157352 229724
rect 166258 229712 166264 229724
rect 166316 229712 166322 229764
rect 171042 229712 171048 229764
rect 171100 229752 171106 229764
rect 219986 229752 219992 229764
rect 171100 229724 219992 229752
rect 171100 229712 171106 229724
rect 219986 229712 219992 229724
rect 220044 229712 220050 229764
rect 246114 229752 246120 229764
rect 224926 229724 246120 229752
rect 148134 229576 148140 229628
rect 148192 229616 148198 229628
rect 155954 229616 155960 229628
rect 148192 229588 155960 229616
rect 148192 229576 148198 229588
rect 155954 229576 155960 229588
rect 156012 229576 156018 229628
rect 157334 229576 157340 229628
rect 157392 229616 157398 229628
rect 157392 229588 214604 229616
rect 157392 229576 157398 229588
rect 147180 229520 147996 229548
rect 156800 229520 157012 229548
rect 147180 229508 147186 229520
rect 102134 229440 102140 229492
rect 102192 229480 102198 229492
rect 143994 229480 144000 229492
rect 102192 229452 144000 229480
rect 102192 229440 102198 229452
rect 143994 229440 144000 229452
rect 144052 229440 144058 229492
rect 144178 229440 144184 229492
rect 144236 229480 144242 229492
rect 146938 229480 146944 229492
rect 144236 229452 146944 229480
rect 144236 229440 144242 229452
rect 146938 229440 146944 229452
rect 146996 229440 147002 229492
rect 156800 229480 156828 229520
rect 148060 229452 156828 229480
rect 156984 229480 157012 229520
rect 210050 229480 210056 229492
rect 156984 229452 210056 229480
rect 111058 229304 111064 229356
rect 111116 229344 111122 229356
rect 147582 229344 147588 229356
rect 111116 229316 147588 229344
rect 111116 229304 111122 229316
rect 147582 229304 147588 229316
rect 147640 229304 147646 229356
rect 147766 229304 147772 229356
rect 147824 229344 147830 229356
rect 148060 229344 148088 229452
rect 210050 229440 210056 229452
rect 210108 229440 210114 229492
rect 214576 229480 214604 229588
rect 214742 229576 214748 229628
rect 214800 229616 214806 229628
rect 224926 229616 224954 229724
rect 246114 229712 246120 229724
rect 246172 229712 246178 229764
rect 256510 229712 256516 229764
rect 256568 229752 256574 229764
rect 297634 229752 297640 229764
rect 256568 229724 297640 229752
rect 256568 229712 256574 229724
rect 297634 229712 297640 229724
rect 297692 229712 297698 229764
rect 318058 229712 318064 229764
rect 318116 229752 318122 229764
rect 318116 229724 335354 229752
rect 318116 229712 318122 229724
rect 266722 229616 266728 229628
rect 214800 229588 224954 229616
rect 229066 229588 266728 229616
rect 214800 229576 214806 229588
rect 220354 229480 220360 229492
rect 214576 229452 220360 229480
rect 220354 229440 220360 229452
rect 220412 229440 220418 229492
rect 220722 229440 220728 229492
rect 220780 229480 220786 229492
rect 229066 229480 229094 229588
rect 266722 229576 266728 229588
rect 266780 229576 266786 229628
rect 296990 229576 296996 229628
rect 297048 229616 297054 229628
rect 323394 229616 323400 229628
rect 297048 229588 323400 229616
rect 297048 229576 297054 229588
rect 323394 229576 323400 229588
rect 323452 229576 323458 229628
rect 335326 229616 335354 229724
rect 345014 229712 345020 229764
rect 345072 229752 345078 229764
rect 360746 229752 360752 229764
rect 345072 229724 360752 229752
rect 345072 229712 345078 229724
rect 360746 229712 360752 229724
rect 360804 229712 360810 229764
rect 361206 229712 361212 229764
rect 361264 229752 361270 229764
rect 378778 229752 378784 229764
rect 361264 229724 378784 229752
rect 361264 229712 361270 229724
rect 378778 229712 378784 229724
rect 378836 229712 378842 229764
rect 391198 229712 391204 229764
rect 391256 229752 391262 229764
rect 398742 229752 398748 229764
rect 391256 229724 398748 229752
rect 391256 229712 391262 229724
rect 398742 229712 398748 229724
rect 398800 229712 398806 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 410886 229712 410892 229764
rect 410944 229752 410950 229764
rect 417418 229752 417424 229764
rect 410944 229724 417424 229752
rect 410944 229712 410950 229724
rect 417418 229712 417424 229724
rect 417476 229712 417482 229764
rect 467006 229712 467012 229764
rect 467064 229752 467070 229764
rect 473998 229752 474004 229764
rect 467064 229724 474004 229752
rect 467064 229712 467070 229724
rect 473998 229712 474004 229724
rect 474056 229712 474062 229764
rect 474200 229684 474228 229860
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 489914 229888 489920 229900
rect 481876 229860 489920 229888
rect 481876 229848 481882 229860
rect 489914 229848 489920 229860
rect 489972 229848 489978 229900
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 506566 229888 506572 229900
rect 496044 229860 506572 229888
rect 496044 229848 496050 229860
rect 506566 229848 506572 229860
rect 506624 229848 506630 229900
rect 510798 229848 510804 229900
rect 510856 229888 510862 229900
rect 511902 229888 511908 229900
rect 510856 229860 511908 229888
rect 510856 229848 510862 229860
rect 511902 229848 511908 229860
rect 511960 229848 511966 229900
rect 517238 229848 517244 229900
rect 517296 229888 517302 229900
rect 525978 229888 525984 229900
rect 517296 229860 525984 229888
rect 517296 229848 517302 229860
rect 525978 229848 525984 229860
rect 526036 229848 526042 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 559558 229888 559564 229900
rect 536616 229860 559564 229888
rect 536616 229848 536622 229860
rect 559558 229848 559564 229860
rect 559616 229848 559622 229900
rect 476022 229780 476028 229832
rect 476080 229820 476086 229832
rect 478598 229820 478604 229832
rect 476080 229792 478604 229820
rect 476080 229780 476086 229792
rect 478598 229780 478604 229792
rect 478656 229780 478662 229832
rect 673454 229780 673460 229832
rect 673512 229820 673518 229832
rect 673512 229792 674360 229820
rect 673512 229780 673518 229792
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 488074 229752 488080 229764
rect 479300 229724 488080 229752
rect 479300 229712 479306 229724
rect 488074 229712 488080 229724
rect 488132 229712 488138 229764
rect 492122 229712 492128 229764
rect 492180 229752 492186 229764
rect 505186 229752 505192 229764
rect 492180 229724 505192 229752
rect 492180 229712 492186 229724
rect 505186 229712 505192 229724
rect 505244 229712 505250 229764
rect 507578 229712 507584 229764
rect 507636 229752 507642 229764
rect 516778 229752 516784 229764
rect 507636 229724 516784 229752
rect 507636 229712 507642 229724
rect 516778 229712 516784 229724
rect 516836 229712 516842 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534810 229752 534816 229764
rect 523092 229724 534816 229752
rect 523092 229712 523098 229724
rect 534810 229712 534816 229724
rect 534868 229712 534874 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 566458 229752 566464 229764
rect 538548 229724 566464 229752
rect 538548 229712 538554 229724
rect 566458 229712 566464 229724
rect 566516 229712 566522 229764
rect 476758 229684 476764 229696
rect 474200 229656 476764 229684
rect 476758 229644 476764 229656
rect 476816 229644 476822 229696
rect 345290 229616 345296 229628
rect 335326 229588 345296 229616
rect 345290 229576 345296 229588
rect 345348 229576 345354 229628
rect 463786 229576 463792 229628
rect 463844 229616 463850 229628
rect 465718 229616 465724 229628
rect 463844 229588 465724 229616
rect 463844 229576 463850 229588
rect 465718 229576 465724 229588
rect 465776 229576 465782 229628
rect 509510 229576 509516 229628
rect 509568 229616 509574 229628
rect 515398 229616 515404 229628
rect 509568 229588 515404 229616
rect 509568 229576 509574 229588
rect 515398 229576 515404 229588
rect 515456 229576 515462 229628
rect 530118 229576 530124 229628
rect 530176 229616 530182 229628
rect 531130 229616 531136 229628
rect 530176 229588 531136 229616
rect 530176 229576 530182 229588
rect 531130 229576 531136 229588
rect 531188 229576 531194 229628
rect 538306 229616 538312 229628
rect 538186 229588 538312 229616
rect 384298 229508 384304 229560
rect 384356 229548 384362 229560
rect 389082 229548 389088 229560
rect 384356 229520 389088 229548
rect 384356 229508 384362 229520
rect 389082 229508 389088 229520
rect 389140 229508 389146 229560
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 451918 229548 451924 229560
rect 449032 229520 451924 229548
rect 449032 229508 449038 229520
rect 451918 229508 451924 229520
rect 451976 229508 451982 229560
rect 220780 229452 229094 229480
rect 220780 229440 220786 229452
rect 231118 229440 231124 229492
rect 231176 229480 231182 229492
rect 271874 229480 271880 229492
rect 231176 229452 271880 229480
rect 231176 229440 231182 229452
rect 271874 229440 271880 229452
rect 271932 229440 271938 229492
rect 465442 229440 465448 229492
rect 465500 229480 465506 229492
rect 467466 229480 467472 229492
rect 465500 229452 467472 229480
rect 465500 229440 465506 229452
rect 467466 229440 467472 229452
rect 467524 229440 467530 229492
rect 488258 229440 488264 229492
rect 488316 229480 488322 229492
rect 490374 229480 490380 229492
rect 488316 229452 490380 229480
rect 488316 229440 488322 229452
rect 490374 229440 490380 229452
rect 490432 229440 490438 229492
rect 530762 229440 530768 229492
rect 530820 229480 530826 229492
rect 538186 229480 538214 229588
rect 538306 229576 538312 229588
rect 538364 229576 538370 229628
rect 673914 229576 673920 229628
rect 673972 229616 673978 229628
rect 673972 229588 674268 229616
rect 673972 229576 673978 229588
rect 530820 229452 538214 229480
rect 530820 229440 530826 229452
rect 450906 229372 450912 229424
rect 450964 229412 450970 229424
rect 453022 229412 453028 229424
rect 450964 229384 453028 229412
rect 450964 229372 450970 229384
rect 453022 229372 453028 229384
rect 453080 229372 453086 229424
rect 674104 229356 674156 229362
rect 147824 229316 148088 229344
rect 147824 229304 147830 229316
rect 151170 229304 151176 229356
rect 151228 229344 151234 229356
rect 151228 229316 153608 229344
rect 151228 229304 151234 229316
rect 123478 229168 123484 229220
rect 123536 229208 123542 229220
rect 153378 229208 153384 229220
rect 123536 229180 153384 229208
rect 123536 229168 123542 229180
rect 153378 229168 153384 229180
rect 153436 229168 153442 229220
rect 153580 229208 153608 229316
rect 153838 229304 153844 229356
rect 153896 229344 153902 229356
rect 156506 229344 156512 229356
rect 153896 229316 156512 229344
rect 153896 229304 153902 229316
rect 156506 229304 156512 229316
rect 156564 229304 156570 229356
rect 157058 229304 157064 229356
rect 157116 229344 157122 229356
rect 215202 229344 215208 229356
rect 157116 229316 215208 229344
rect 157116 229304 157122 229316
rect 215202 229304 215208 229316
rect 215260 229304 215266 229356
rect 246482 229304 246488 229356
rect 246540 229344 246546 229356
rect 282178 229344 282184 229356
rect 246540 229316 282184 229344
rect 246540 229304 246546 229316
rect 282178 229304 282184 229316
rect 282236 229304 282242 229356
rect 413830 229304 413836 229356
rect 413888 229344 413894 229356
rect 419994 229344 420000 229356
rect 413888 229316 420000 229344
rect 413888 229304 413894 229316
rect 419994 229304 420000 229316
rect 420052 229304 420058 229356
rect 674104 229298 674156 229304
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451734 229276 451740 229288
rect 450320 229248 451740 229276
rect 450320 229236 450326 229248
rect 451734 229236 451740 229248
rect 451792 229236 451798 229288
rect 495342 229236 495348 229288
rect 495400 229276 495406 229288
rect 500218 229276 500224 229288
rect 495400 229248 500224 229276
rect 495400 229236 495406 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 505646 229236 505652 229288
rect 505704 229276 505710 229288
rect 510614 229276 510620 229288
rect 505704 229248 510620 229276
rect 505704 229236 505710 229248
rect 510614 229236 510620 229248
rect 510672 229236 510678 229288
rect 513374 229236 513380 229288
rect 513432 229276 513438 229288
rect 519354 229276 519360 229288
rect 513432 229248 519360 229276
rect 513432 229236 513438 229248
rect 519354 229236 519360 229248
rect 519412 229236 519418 229288
rect 161750 229208 161756 229220
rect 153580 229180 161756 229208
rect 161750 229168 161756 229180
rect 161808 229168 161814 229220
rect 184658 229168 184664 229220
rect 184716 229208 184722 229220
rect 240962 229208 240968 229220
rect 184716 229180 240968 229208
rect 184716 229168 184722 229180
rect 240962 229168 240968 229180
rect 241020 229168 241026 229220
rect 167104 229112 167500 229140
rect 100662 229032 100668 229084
rect 100720 229072 100726 229084
rect 100720 229044 103514 229072
rect 100720 229032 100726 229044
rect 103486 228936 103514 229044
rect 106182 229032 106188 229084
rect 106240 229072 106246 229084
rect 142982 229072 142988 229084
rect 106240 229044 142988 229072
rect 106240 229032 106246 229044
rect 142982 229032 142988 229044
rect 143040 229032 143046 229084
rect 143442 229032 143448 229084
rect 143500 229072 143506 229084
rect 146202 229072 146208 229084
rect 143500 229044 146208 229072
rect 143500 229032 143506 229044
rect 146202 229032 146208 229044
rect 146260 229032 146266 229084
rect 146386 229032 146392 229084
rect 146444 229072 146450 229084
rect 167104 229072 167132 229112
rect 146444 229044 167132 229072
rect 167472 229072 167500 229112
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 503714 229100 503720 229152
rect 503772 229140 503778 229152
rect 509878 229140 509884 229152
rect 503772 229112 509884 229140
rect 503772 229100 503778 229112
rect 509878 229100 509884 229112
rect 509936 229100 509942 229152
rect 519170 229100 519176 229152
rect 519228 229140 519234 229152
rect 519228 229112 521654 229140
rect 519228 229100 519234 229112
rect 205542 229072 205548 229084
rect 167472 229044 205548 229072
rect 146444 229032 146450 229044
rect 205542 229032 205548 229044
rect 205600 229032 205606 229084
rect 206002 229032 206008 229084
rect 206060 229072 206066 229084
rect 214374 229072 214380 229084
rect 206060 229044 214380 229072
rect 206060 229032 206066 229044
rect 214374 229032 214380 229044
rect 214432 229032 214438 229084
rect 214742 229032 214748 229084
rect 214800 229072 214806 229084
rect 257062 229072 257068 229084
rect 214800 229044 257068 229072
rect 214800 229032 214806 229044
rect 257062 229032 257068 229044
rect 257120 229032 257126 229084
rect 257522 229032 257528 229084
rect 257580 229072 257586 229084
rect 296346 229072 296352 229084
rect 257580 229044 296352 229072
rect 257580 229032 257586 229044
rect 296346 229032 296352 229044
rect 296404 229032 296410 229084
rect 302142 229032 302148 229084
rect 302200 229072 302206 229084
rect 331122 229072 331128 229084
rect 302200 229044 331128 229072
rect 302200 229032 302206 229044
rect 331122 229032 331128 229044
rect 331180 229032 331186 229084
rect 521626 229004 521654 229112
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 529934 229140 529940 229152
rect 525024 229112 529940 229140
rect 525024 229100 525030 229112
rect 529934 229100 529940 229112
rect 529992 229100 529998 229152
rect 660942 229100 660948 229152
rect 661000 229140 661006 229152
rect 665450 229140 665456 229152
rect 661000 229112 665456 229140
rect 661000 229100 661006 229112
rect 665450 229100 665456 229112
rect 665508 229100 665514 229152
rect 673472 229112 674038 229140
rect 521626 228976 528554 229004
rect 169294 228936 169300 228948
rect 103486 228908 169300 228936
rect 169294 228896 169300 228908
rect 169352 228896 169358 228948
rect 172330 228896 172336 228948
rect 172388 228936 172394 228948
rect 179690 228936 179696 228948
rect 172388 228908 179696 228936
rect 172388 228896 172394 228908
rect 179690 228896 179696 228908
rect 179748 228896 179754 228948
rect 180058 228896 180064 228948
rect 180116 228936 180122 228948
rect 180116 228908 220124 228936
rect 180116 228896 180122 228908
rect 93762 228760 93768 228812
rect 93820 228800 93826 228812
rect 166810 228800 166816 228812
rect 93820 228772 166816 228800
rect 93820 228760 93826 228772
rect 166810 228760 166816 228772
rect 166868 228760 166874 228812
rect 172146 228760 172152 228812
rect 172204 228800 172210 228812
rect 174630 228800 174636 228812
rect 172204 228772 174636 228800
rect 172204 228760 172210 228772
rect 174630 228760 174636 228772
rect 174688 228760 174694 228812
rect 174814 228760 174820 228812
rect 174872 228800 174878 228812
rect 219802 228800 219808 228812
rect 174872 228772 219808 228800
rect 174872 228760 174878 228772
rect 219802 228760 219808 228772
rect 219860 228760 219866 228812
rect 220096 228800 220124 228908
rect 220354 228896 220360 228948
rect 220412 228936 220418 228948
rect 246758 228936 246764 228948
rect 220412 228908 246764 228936
rect 220412 228896 220418 228908
rect 246758 228896 246764 228908
rect 246816 228896 246822 228948
rect 257706 228896 257712 228948
rect 257764 228936 257770 228948
rect 299566 228936 299572 228948
rect 257764 228908 299572 228936
rect 257764 228896 257770 228908
rect 299566 228896 299572 228908
rect 299624 228896 299630 228948
rect 300670 228896 300676 228948
rect 300728 228936 300734 228948
rect 330478 228936 330484 228948
rect 300728 228908 330484 228936
rect 300728 228896 300734 228908
rect 330478 228896 330484 228908
rect 330536 228896 330542 228948
rect 502426 228896 502432 228948
rect 502484 228936 502490 228948
rect 521010 228936 521016 228948
rect 502484 228908 521016 228936
rect 502484 228896 502490 228908
rect 521010 228896 521016 228908
rect 521068 228896 521074 228948
rect 528526 228936 528554 228976
rect 673472 228948 673500 229112
rect 542814 228936 542820 228948
rect 528526 228908 542820 228936
rect 542814 228896 542820 228908
rect 542872 228896 542878 228948
rect 673454 228896 673460 228948
rect 673512 228896 673518 228948
rect 226150 228800 226156 228812
rect 220096 228772 226156 228800
rect 226150 228760 226156 228772
rect 226208 228760 226214 228812
rect 238570 228760 238576 228812
rect 238628 228800 238634 228812
rect 282822 228800 282828 228812
rect 238628 228772 282828 228800
rect 238628 228760 238634 228772
rect 282822 228760 282828 228772
rect 282880 228760 282886 228812
rect 296622 228760 296628 228812
rect 296680 228800 296686 228812
rect 329190 228800 329196 228812
rect 296680 228772 329196 228800
rect 296680 228760 296686 228772
rect 329190 228760 329196 228772
rect 329248 228760 329254 228812
rect 336458 228760 336464 228812
rect 336516 228800 336522 228812
rect 358814 228800 358820 228812
rect 336516 228772 358820 228800
rect 336516 228760 336522 228772
rect 358814 228760 358820 228772
rect 358872 228760 358878 228812
rect 359918 228760 359924 228812
rect 359976 228800 359982 228812
rect 376846 228800 376852 228812
rect 359976 228772 376852 228800
rect 359976 228760 359982 228772
rect 376846 228760 376852 228772
rect 376904 228760 376910 228812
rect 478874 228760 478880 228812
rect 478932 228800 478938 228812
rect 490190 228800 490196 228812
rect 478932 228772 490196 228800
rect 478932 228760 478938 228772
rect 490190 228760 490196 228772
rect 490248 228760 490254 228812
rect 518526 228760 518532 228812
rect 518584 228800 518590 228812
rect 541618 228800 541624 228812
rect 518584 228772 541624 228800
rect 518584 228760 518590 228772
rect 541618 228760 541624 228772
rect 541676 228760 541682 228812
rect 67542 228624 67548 228676
rect 67600 228664 67606 228676
rect 67600 228636 142844 228664
rect 67600 228624 67606 228636
rect 61654 228488 61660 228540
rect 61712 228528 61718 228540
rect 142614 228528 142620 228540
rect 61712 228500 142620 228528
rect 61712 228488 61718 228500
rect 142614 228488 142620 228500
rect 142672 228488 142678 228540
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 141142 228392 141148 228404
rect 57296 228364 141148 228392
rect 57296 228352 57302 228364
rect 141142 228352 141148 228364
rect 141200 228352 141206 228404
rect 142816 228392 142844 228636
rect 142982 228624 142988 228676
rect 143040 228664 143046 228676
rect 152458 228664 152464 228676
rect 143040 228636 152464 228664
rect 143040 228624 143046 228636
rect 152458 228624 152464 228636
rect 152516 228624 152522 228676
rect 153102 228624 153108 228676
rect 153160 228664 153166 228676
rect 153160 228636 209774 228664
rect 153160 228624 153166 228636
rect 142982 228488 142988 228540
rect 143040 228528 143046 228540
rect 145926 228528 145932 228540
rect 143040 228500 145932 228528
rect 143040 228488 143046 228500
rect 145926 228488 145932 228500
rect 145984 228488 145990 228540
rect 146110 228488 146116 228540
rect 146168 228528 146174 228540
rect 202414 228528 202420 228540
rect 146168 228500 202420 228528
rect 146168 228488 146174 228500
rect 202414 228488 202420 228500
rect 202472 228488 202478 228540
rect 209746 228528 209774 228636
rect 214374 228624 214380 228676
rect 214432 228664 214438 228676
rect 220354 228664 220360 228676
rect 214432 228636 220360 228664
rect 214432 228624 214438 228636
rect 220354 228624 220360 228636
rect 220412 228624 220418 228676
rect 220538 228624 220544 228676
rect 220596 228664 220602 228676
rect 264790 228664 264796 228676
rect 220596 228636 264796 228664
rect 220596 228624 220602 228636
rect 264790 228624 264796 228636
rect 264848 228624 264854 228676
rect 285490 228624 285496 228676
rect 285548 228664 285554 228676
rect 318886 228664 318892 228676
rect 285548 228636 318892 228664
rect 285548 228624 285554 228636
rect 318886 228624 318892 228636
rect 318944 228624 318950 228676
rect 325510 228624 325516 228676
rect 325568 228664 325574 228676
rect 349154 228664 349160 228676
rect 325568 228636 349160 228664
rect 325568 228624 325574 228636
rect 349154 228624 349160 228636
rect 349212 228624 349218 228676
rect 350166 228624 350172 228676
rect 350224 228664 350230 228676
rect 369118 228664 369124 228676
rect 350224 228636 369124 228664
rect 350224 228624 350230 228636
rect 369118 228624 369124 228636
rect 369176 228624 369182 228676
rect 377766 228624 377772 228676
rect 377824 228664 377830 228676
rect 390370 228664 390376 228676
rect 377824 228636 390376 228664
rect 377824 228624 377830 228636
rect 390370 228624 390376 228636
rect 390428 228624 390434 228676
rect 498562 228624 498568 228676
rect 498620 228664 498626 228676
rect 515766 228664 515772 228676
rect 498620 228636 515772 228664
rect 498620 228624 498626 228636
rect 515766 228624 515772 228636
rect 515824 228624 515830 228676
rect 517882 228624 517888 228676
rect 517940 228664 517946 228676
rect 539410 228664 539416 228676
rect 517940 228636 539416 228664
rect 517940 228624 517946 228636
rect 539410 228624 539416 228636
rect 539468 228624 539474 228676
rect 539594 228624 539600 228676
rect 539652 228664 539658 228676
rect 555970 228664 555976 228676
rect 539652 228636 555976 228664
rect 539652 228624 539658 228636
rect 555970 228624 555976 228636
rect 556028 228624 556034 228676
rect 215846 228528 215852 228540
rect 209746 228500 215852 228528
rect 215846 228488 215852 228500
rect 215904 228488 215910 228540
rect 216214 228488 216220 228540
rect 216272 228528 216278 228540
rect 219618 228528 219624 228540
rect 216272 228500 219624 228528
rect 216272 228488 216278 228500
rect 219618 228488 219624 228500
rect 219676 228488 219682 228540
rect 219986 228488 219992 228540
rect 220044 228528 220050 228540
rect 260282 228528 260288 228540
rect 220044 228500 260288 228528
rect 220044 228488 220050 228500
rect 260282 228488 260288 228500
rect 260340 228488 260346 228540
rect 268930 228488 268936 228540
rect 268988 228528 268994 228540
rect 306006 228528 306012 228540
rect 268988 228500 306012 228528
rect 268988 228488 268994 228500
rect 306006 228488 306012 228500
rect 306064 228488 306070 228540
rect 313918 228488 313924 228540
rect 313976 228528 313982 228540
rect 320818 228528 320824 228540
rect 313976 228500 320824 228528
rect 313976 228488 313982 228500
rect 320818 228488 320824 228500
rect 320876 228488 320882 228540
rect 326890 228488 326896 228540
rect 326948 228528 326954 228540
rect 351086 228528 351092 228540
rect 326948 228500 351092 228528
rect 326948 228488 326954 228500
rect 351086 228488 351092 228500
rect 351144 228488 351150 228540
rect 354582 228488 354588 228540
rect 354640 228528 354646 228540
rect 372338 228528 372344 228540
rect 354640 228500 372344 228528
rect 354640 228488 354646 228500
rect 372338 228488 372344 228500
rect 372396 228488 372402 228540
rect 373442 228488 373448 228540
rect 373500 228528 373506 228540
rect 387150 228528 387156 228540
rect 373500 228500 387156 228528
rect 373500 228488 373506 228500
rect 387150 228488 387156 228500
rect 387208 228488 387214 228540
rect 390462 228488 390468 228540
rect 390520 228528 390526 228540
rect 400030 228528 400036 228540
rect 390520 228500 400036 228528
rect 390520 228488 390526 228500
rect 400030 228488 400036 228500
rect 400088 228488 400094 228540
rect 407758 228528 407764 228540
rect 400232 228500 407764 228528
rect 148870 228392 148876 228404
rect 142816 228364 148876 228392
rect 148870 228352 148876 228364
rect 148928 228352 148934 228404
rect 152458 228352 152464 228404
rect 152516 228392 152522 228404
rect 166810 228392 166816 228404
rect 152516 228364 166816 228392
rect 152516 228352 152522 228364
rect 166810 228352 166816 228364
rect 166868 228352 166874 228404
rect 166948 228352 166954 228404
rect 167006 228392 167012 228404
rect 214558 228392 214564 228404
rect 167006 228364 214564 228392
rect 167006 228352 167012 228364
rect 214558 228352 214564 228364
rect 214616 228352 214622 228404
rect 217502 228352 217508 228404
rect 217560 228392 217566 228404
rect 221458 228392 221464 228404
rect 217560 228364 221464 228392
rect 217560 228352 217566 228364
rect 221458 228352 221464 228364
rect 221516 228352 221522 228404
rect 224586 228352 224592 228404
rect 224644 228392 224650 228404
rect 273806 228392 273812 228404
rect 224644 228364 273812 228392
rect 224644 228352 224650 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 274266 228352 274272 228404
rect 274324 228392 274330 228404
rect 312446 228392 312452 228404
rect 274324 228364 312452 228392
rect 274324 228352 274330 228364
rect 312446 228352 312452 228364
rect 312504 228352 312510 228404
rect 320082 228352 320088 228404
rect 320140 228392 320146 228404
rect 346854 228392 346860 228404
rect 320140 228364 346860 228392
rect 320140 228352 320146 228364
rect 346854 228352 346860 228364
rect 346912 228352 346918 228404
rect 347038 228352 347044 228404
rect 347096 228392 347102 228404
rect 365898 228392 365904 228404
rect 347096 228364 365904 228392
rect 347096 228352 347102 228364
rect 365898 228352 365904 228364
rect 365956 228352 365962 228404
rect 371142 228352 371148 228404
rect 371200 228392 371206 228404
rect 385218 228392 385224 228404
rect 371200 228364 385224 228392
rect 371200 228352 371206 228364
rect 385218 228352 385224 228364
rect 385276 228352 385282 228404
rect 386230 228352 386236 228404
rect 386288 228392 386294 228404
rect 397454 228392 397460 228404
rect 386288 228364 397460 228392
rect 386288 228352 386294 228364
rect 397454 228352 397460 228364
rect 397512 228352 397518 228404
rect 112806 228216 112812 228268
rect 112864 228256 112870 228268
rect 184934 228256 184940 228268
rect 112864 228228 184940 228256
rect 112864 228216 112870 228228
rect 184934 228216 184940 228228
rect 184992 228216 184998 228268
rect 189718 228216 189724 228268
rect 189776 228256 189782 228268
rect 239030 228256 239036 228268
rect 189776 228228 239036 228256
rect 189776 228216 189782 228228
rect 239030 228216 239036 228228
rect 239088 228216 239094 228268
rect 254946 228216 254952 228268
rect 255004 228256 255010 228268
rect 295702 228256 295708 228268
rect 255004 228228 295708 228256
rect 255004 228216 255010 228228
rect 295702 228216 295708 228228
rect 295760 228216 295766 228268
rect 400232 228256 400260 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 409782 228488 409788 228540
rect 409840 228528 409846 228540
rect 415486 228528 415492 228540
rect 409840 228500 415492 228528
rect 409840 228488 409846 228500
rect 415486 228488 415492 228500
rect 415544 228488 415550 228540
rect 485682 228488 485688 228540
rect 485740 228528 485746 228540
rect 498286 228528 498292 228540
rect 485740 228500 498292 228528
rect 485740 228488 485746 228500
rect 498286 228488 498292 228500
rect 498344 228488 498350 228540
rect 499850 228488 499856 228540
rect 499908 228528 499914 228540
rect 517698 228528 517704 228540
rect 499908 228500 517704 228528
rect 499908 228488 499914 228500
rect 517698 228488 517704 228500
rect 517756 228488 517762 228540
rect 527542 228488 527548 228540
rect 527600 228528 527606 228540
rect 553302 228528 553308 228540
rect 527600 228500 553308 228528
rect 527600 228488 527606 228500
rect 553302 228488 553308 228500
rect 553360 228488 553366 228540
rect 555418 228488 555424 228540
rect 555476 228528 555482 228540
rect 571334 228528 571340 228540
rect 555476 228500 571340 228528
rect 555476 228488 555482 228500
rect 571334 228488 571340 228500
rect 571392 228488 571398 228540
rect 402790 228352 402796 228404
rect 402848 228392 402854 228404
rect 411622 228392 411628 228404
rect 402848 228364 411628 228392
rect 402848 228352 402854 228364
rect 411622 228352 411628 228364
rect 411680 228352 411686 228404
rect 474458 228352 474464 228404
rect 474516 228392 474522 228404
rect 484578 228392 484584 228404
rect 474516 228364 484584 228392
rect 474516 228352 474522 228364
rect 484578 228352 484584 228364
rect 484636 228352 484642 228404
rect 485038 228352 485044 228404
rect 485096 228392 485102 228404
rect 498562 228392 498568 228404
rect 485096 228364 498568 228392
rect 485096 228352 485102 228364
rect 498562 228352 498568 228364
rect 498620 228352 498626 228404
rect 506566 228352 506572 228404
rect 506624 228392 506630 228404
rect 506624 228364 509234 228392
rect 506624 228352 506630 228364
rect 400140 228228 400260 228256
rect 509206 228256 509234 228364
rect 512086 228352 512092 228404
rect 512144 228392 512150 228404
rect 533522 228392 533528 228404
rect 512144 228364 533528 228392
rect 512144 228352 512150 228364
rect 533522 228352 533528 228364
rect 533580 228352 533586 228404
rect 537202 228352 537208 228404
rect 537260 228392 537266 228404
rect 565630 228392 565636 228404
rect 537260 228364 565636 228392
rect 537260 228352 537266 228364
rect 565630 228352 565636 228364
rect 565688 228352 565694 228404
rect 663518 228352 663524 228404
rect 663576 228392 663582 228404
rect 672074 228392 672080 228404
rect 663576 228364 672080 228392
rect 663576 228352 663582 228364
rect 672074 228352 672080 228364
rect 672132 228352 672138 228404
rect 512730 228256 512736 228268
rect 509206 228228 512736 228256
rect 400140 228132 400168 228228
rect 512730 228216 512736 228228
rect 512788 228216 512794 228268
rect 539410 228216 539416 228268
rect 539468 228256 539474 228268
rect 540882 228256 540888 228268
rect 539468 228228 540888 228256
rect 539468 228216 539474 228228
rect 540882 228216 540888 228228
rect 540940 228216 540946 228268
rect 119982 228080 119988 228132
rect 120040 228120 120046 228132
rect 190086 228120 190092 228132
rect 120040 228092 190092 228120
rect 120040 228080 120046 228092
rect 190086 228080 190092 228092
rect 190144 228080 190150 228132
rect 192938 228080 192944 228132
rect 192996 228120 193002 228132
rect 192996 228092 200114 228120
rect 192996 228080 193002 228092
rect 126698 227944 126704 227996
rect 126756 227984 126762 227996
rect 195238 227984 195244 227996
rect 126756 227956 195244 227984
rect 126756 227944 126762 227956
rect 195238 227944 195244 227956
rect 195296 227944 195302 227996
rect 200086 227984 200114 228092
rect 202414 228080 202420 228132
rect 202472 228120 202478 228132
rect 210694 228120 210700 228132
rect 202472 228092 210700 228120
rect 202472 228080 202478 228092
rect 210694 228080 210700 228092
rect 210752 228080 210758 228132
rect 213914 228080 213920 228132
rect 213972 228120 213978 228132
rect 214374 228120 214380 228132
rect 213972 228092 214380 228120
rect 213972 228080 213978 228092
rect 214374 228080 214380 228092
rect 214432 228080 214438 228132
rect 214558 228080 214564 228132
rect 214616 228120 214622 228132
rect 214616 228092 215294 228120
rect 214616 228080 214622 228092
rect 206002 227984 206008 227996
rect 200086 227956 206008 227984
rect 206002 227944 206008 227956
rect 206060 227944 206066 227996
rect 214742 227984 214748 227996
rect 209746 227956 214748 227984
rect 88242 227808 88248 227860
rect 88300 227848 88306 227860
rect 95234 227848 95240 227860
rect 88300 227820 95240 227848
rect 88300 227808 88306 227820
rect 95234 227808 95240 227820
rect 95292 227808 95298 227860
rect 133506 227808 133512 227860
rect 133564 227848 133570 227860
rect 200390 227848 200396 227860
rect 133564 227820 200396 227848
rect 133564 227808 133570 227820
rect 200390 227808 200396 227820
rect 200448 227808 200454 227860
rect 203518 227808 203524 227860
rect 203576 227848 203582 227860
rect 203576 227820 205128 227848
rect 203576 227808 203582 227820
rect 42426 227672 42432 227724
rect 42484 227712 42490 227724
rect 43254 227712 43260 227724
rect 42484 227684 43260 227712
rect 42484 227672 42490 227684
rect 43254 227672 43260 227684
rect 43312 227672 43318 227724
rect 64782 227672 64788 227724
rect 64840 227712 64846 227724
rect 111058 227712 111064 227724
rect 64840 227684 111064 227712
rect 64840 227672 64846 227684
rect 111058 227672 111064 227684
rect 111116 227672 111122 227724
rect 117222 227672 117228 227724
rect 117280 227712 117286 227724
rect 187510 227712 187516 227724
rect 117280 227684 187516 227712
rect 117280 227672 117286 227684
rect 187510 227672 187516 227684
rect 187568 227672 187574 227724
rect 187694 227672 187700 227724
rect 187752 227712 187758 227724
rect 187752 227684 193076 227712
rect 187752 227672 187758 227684
rect 110138 227536 110144 227588
rect 110196 227576 110202 227588
rect 182358 227576 182364 227588
rect 110196 227548 182364 227576
rect 110196 227536 110202 227548
rect 182358 227536 182364 227548
rect 182416 227536 182422 227588
rect 185394 227536 185400 227588
rect 185452 227576 185458 227588
rect 192662 227576 192668 227588
rect 185452 227548 192668 227576
rect 185452 227536 185458 227548
rect 192662 227536 192668 227548
rect 192720 227536 192726 227588
rect 193048 227576 193076 227684
rect 200022 227672 200028 227724
rect 200080 227712 200086 227724
rect 204898 227712 204904 227724
rect 200080 227684 204904 227712
rect 200080 227672 200086 227684
rect 204898 227672 204904 227684
rect 204956 227672 204962 227724
rect 205100 227712 205128 227820
rect 205450 227808 205456 227860
rect 205508 227848 205514 227860
rect 209746 227848 209774 227956
rect 214742 227944 214748 227956
rect 214800 227944 214806 227996
rect 215266 227984 215294 228092
rect 219802 228080 219808 228132
rect 219860 228120 219866 228132
rect 231302 228120 231308 228132
rect 219860 228092 231308 228120
rect 219860 228080 219866 228092
rect 231302 228080 231308 228092
rect 231360 228080 231366 228132
rect 233878 228080 233884 228132
rect 233936 228120 233942 228132
rect 272518 228120 272524 228132
rect 233936 228092 272524 228120
rect 233936 228080 233942 228092
rect 272518 228080 272524 228092
rect 272576 228080 272582 228132
rect 400122 228080 400128 228132
rect 400180 228080 400186 228132
rect 415026 228012 415032 228064
rect 415084 228052 415090 228064
rect 421926 228052 421932 228064
rect 415084 228024 421932 228052
rect 415084 228012 415090 228024
rect 421926 228012 421932 228024
rect 421984 228012 421990 228064
rect 220998 227984 221004 227996
rect 215266 227956 221004 227984
rect 220998 227944 221004 227956
rect 221056 227944 221062 227996
rect 221458 227944 221464 227996
rect 221516 227984 221522 227996
rect 251266 227984 251272 227996
rect 221516 227956 251272 227984
rect 221516 227944 221522 227956
rect 251266 227944 251272 227956
rect 251324 227944 251330 227996
rect 416682 227876 416688 227928
rect 416740 227916 416746 227928
rect 420638 227916 420644 227928
rect 416740 227888 420644 227916
rect 416740 227876 416746 227888
rect 420638 227876 420644 227888
rect 420696 227876 420702 227928
rect 447042 227876 447048 227928
rect 447100 227916 447106 227928
rect 450538 227916 450544 227928
rect 447100 227888 450544 227916
rect 447100 227876 447106 227888
rect 450538 227876 450544 227888
rect 450596 227876 450602 227928
rect 205508 227820 209774 227848
rect 205508 227808 205514 227820
rect 210970 227808 210976 227860
rect 211028 227848 211034 227860
rect 219986 227848 219992 227860
rect 211028 227820 219992 227848
rect 211028 227808 211034 227820
rect 219986 227808 219992 227820
rect 220044 227808 220050 227860
rect 226150 227808 226156 227860
rect 226208 227848 226214 227860
rect 233878 227848 233884 227860
rect 226208 227820 233884 227848
rect 226208 227808 226214 227820
rect 233878 227808 233884 227820
rect 233936 227808 233942 227860
rect 239306 227808 239312 227860
rect 239364 227848 239370 227860
rect 243538 227848 243544 227860
rect 239364 227820 243544 227848
rect 239364 227808 239370 227820
rect 243538 227808 243544 227820
rect 243596 227808 243602 227860
rect 246298 227808 246304 227860
rect 246356 227848 246362 227860
rect 248690 227848 248696 227860
rect 246356 227820 248696 227848
rect 246356 227808 246362 227820
rect 248690 227808 248696 227820
rect 248748 227808 248754 227860
rect 249058 227808 249064 227860
rect 249116 227848 249122 227860
rect 253842 227848 253848 227860
rect 249116 227820 253848 227848
rect 249116 227808 249122 227820
rect 253842 227808 253848 227820
rect 253900 227808 253906 227860
rect 331030 227740 331036 227792
rect 331088 227780 331094 227792
rect 334250 227780 334256 227792
rect 331088 227752 334256 227780
rect 331088 227740 331094 227752
rect 334250 227740 334256 227752
rect 334308 227740 334314 227792
rect 351086 227740 351092 227792
rect 351144 227780 351150 227792
rect 353018 227780 353024 227792
rect 351144 227752 353024 227780
rect 351144 227740 351150 227752
rect 353018 227740 353024 227752
rect 353076 227740 353082 227792
rect 371786 227740 371792 227792
rect 371844 227780 371850 227792
rect 373626 227780 373632 227792
rect 371844 227752 373632 227780
rect 371844 227740 371850 227752
rect 373626 227740 373632 227752
rect 373684 227740 373690 227792
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 420638 227740 420644 227792
rect 420696 227780 420702 227792
rect 423858 227780 423864 227792
rect 420696 227752 423864 227780
rect 420696 227740 420702 227752
rect 423858 227740 423864 227752
rect 423916 227740 423922 227792
rect 471514 227740 471520 227792
rect 471572 227780 471578 227792
rect 479518 227780 479524 227792
rect 471572 227752 479524 227780
rect 471572 227740 471578 227752
rect 479518 227740 479524 227752
rect 479576 227740 479582 227792
rect 489914 227740 489920 227792
rect 489972 227780 489978 227792
rect 494514 227780 494520 227792
rect 489972 227752 494520 227780
rect 489972 227740 489978 227752
rect 494514 227740 494520 227752
rect 494572 227740 494578 227792
rect 660482 227740 660488 227792
rect 660540 227780 660546 227792
rect 665174 227780 665180 227792
rect 660540 227752 665180 227780
rect 660540 227740 660546 227752
rect 665174 227740 665180 227752
rect 665232 227740 665238 227792
rect 668946 227740 668952 227792
rect 669004 227780 669010 227792
rect 672718 227780 672724 227792
rect 669004 227752 672724 227780
rect 669004 227740 669010 227752
rect 672718 227740 672724 227752
rect 672776 227740 672782 227792
rect 217778 227712 217784 227724
rect 205100 227684 217784 227712
rect 217778 227672 217784 227684
rect 217836 227672 217842 227724
rect 219802 227672 219808 227724
rect 219860 227712 219866 227724
rect 228726 227712 228732 227724
rect 219860 227684 228732 227712
rect 219860 227672 219866 227684
rect 228726 227672 228732 227684
rect 228784 227672 228790 227724
rect 228910 227672 228916 227724
rect 228968 227712 228974 227724
rect 268010 227712 268016 227724
rect 228968 227684 268016 227712
rect 228968 227672 228974 227684
rect 268010 227672 268016 227684
rect 268068 227672 268074 227724
rect 291010 227672 291016 227724
rect 291068 227712 291074 227724
rect 322106 227712 322112 227724
rect 291068 227684 322112 227712
rect 291068 227672 291074 227684
rect 322106 227672 322112 227684
rect 322164 227672 322170 227724
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 214742 227576 214748 227588
rect 193048 227548 214748 227576
rect 214742 227536 214748 227548
rect 214800 227536 214806 227588
rect 214926 227536 214932 227588
rect 214984 227576 214990 227588
rect 262214 227576 262220 227588
rect 214984 227548 262220 227576
rect 214984 227536 214990 227548
rect 262214 227536 262220 227548
rect 262272 227536 262278 227588
rect 281350 227536 281356 227588
rect 281408 227576 281414 227588
rect 317598 227576 317604 227588
rect 281408 227548 317604 227576
rect 281408 227536 281414 227548
rect 317598 227536 317604 227548
rect 317656 227536 317662 227588
rect 322106 227536 322112 227588
rect 322164 227576 322170 227588
rect 332410 227576 332416 227588
rect 322164 227548 332416 227576
rect 322164 227536 322170 227548
rect 332410 227536 332416 227548
rect 332468 227536 332474 227588
rect 337746 227536 337752 227588
rect 337804 227576 337810 227588
rect 345014 227576 345020 227588
rect 337804 227548 345020 227576
rect 337804 227536 337810 227548
rect 345014 227536 345020 227548
rect 345072 227536 345078 227588
rect 524598 227536 524604 227588
rect 524656 227576 524662 227588
rect 537478 227576 537484 227588
rect 524656 227548 537484 227576
rect 524656 227536 524662 227548
rect 537478 227536 537484 227548
rect 537536 227536 537542 227588
rect 60642 227400 60648 227452
rect 60700 227440 60706 227452
rect 102134 227440 102140 227452
rect 60700 227412 102140 227440
rect 60700 227400 60706 227412
rect 102134 227400 102140 227412
rect 102192 227400 102198 227452
rect 103422 227400 103428 227452
rect 103480 227440 103486 227452
rect 171226 227440 171232 227452
rect 103480 227412 171232 227440
rect 103480 227400 103486 227412
rect 171226 227400 171232 227412
rect 171284 227400 171290 227452
rect 172146 227400 172152 227452
rect 172204 227440 172210 227452
rect 177206 227440 177212 227452
rect 172204 227412 177212 227440
rect 172204 227400 172210 227412
rect 177206 227400 177212 227412
rect 177264 227400 177270 227452
rect 181346 227400 181352 227452
rect 181404 227440 181410 227452
rect 181404 227412 185900 227440
rect 181404 227400 181410 227412
rect 96430 227264 96436 227316
rect 96488 227304 96494 227316
rect 169478 227304 169484 227316
rect 96488 227276 157196 227304
rect 96488 227264 96494 227276
rect 157168 227236 157196 227276
rect 157444 227276 169484 227304
rect 157168 227208 157288 227236
rect 89622 227128 89628 227180
rect 89680 227168 89686 227180
rect 156690 227168 156696 227180
rect 89680 227140 156696 227168
rect 89680 227128 89686 227140
rect 156690 227128 156696 227140
rect 156748 227128 156754 227180
rect 157260 227168 157288 227208
rect 157444 227168 157472 227276
rect 169478 227264 169484 227276
rect 169536 227264 169542 227316
rect 185578 227304 185584 227316
rect 171336 227276 185584 227304
rect 157260 227140 157472 227168
rect 159634 227128 159640 227180
rect 159692 227168 159698 227180
rect 171336 227168 171364 227276
rect 185578 227264 185584 227276
rect 185636 227264 185642 227316
rect 185872 227304 185900 227412
rect 186130 227400 186136 227452
rect 186188 227440 186194 227452
rect 187694 227440 187700 227452
rect 186188 227412 187700 227440
rect 186188 227400 186194 227412
rect 187694 227400 187700 227412
rect 187752 227400 187758 227452
rect 189902 227400 189908 227452
rect 189960 227440 189966 227452
rect 204714 227440 204720 227452
rect 189960 227412 204720 227440
rect 189960 227400 189966 227412
rect 204714 227400 204720 227412
rect 204772 227400 204778 227452
rect 204898 227400 204904 227452
rect 204956 227440 204962 227452
rect 251910 227440 251916 227452
rect 204956 227412 251916 227440
rect 204956 227400 204962 227412
rect 251910 227400 251916 227412
rect 251968 227400 251974 227452
rect 264790 227400 264796 227452
rect 264848 227440 264854 227452
rect 304718 227440 304724 227452
rect 264848 227412 304724 227440
rect 264848 227400 264854 227412
rect 304718 227400 304724 227412
rect 304776 227400 304782 227452
rect 315482 227400 315488 227452
rect 315540 227440 315546 227452
rect 341426 227440 341432 227452
rect 315540 227412 341432 227440
rect 315540 227400 315546 227412
rect 341426 227400 341432 227412
rect 341484 227400 341490 227452
rect 352558 227400 352564 227452
rect 352616 227440 352622 227452
rect 363322 227440 363328 227452
rect 352616 227412 363328 227440
rect 352616 227400 352622 227412
rect 363322 227400 363328 227412
rect 363380 227400 363386 227452
rect 494698 227400 494704 227452
rect 494756 227440 494762 227452
rect 511074 227440 511080 227452
rect 494756 227412 511080 227440
rect 494756 227400 494762 227412
rect 511074 227400 511080 227412
rect 511132 227400 511138 227452
rect 514018 227400 514024 227452
rect 514076 227440 514082 227452
rect 535730 227440 535736 227452
rect 514076 227412 535736 227440
rect 514076 227400 514082 227412
rect 535730 227400 535736 227412
rect 535788 227400 535794 227452
rect 536098 227400 536104 227452
rect 536156 227440 536162 227452
rect 552658 227440 552664 227452
rect 536156 227412 552664 227440
rect 536156 227400 536162 227412
rect 552658 227400 552664 227412
rect 552716 227400 552722 227452
rect 219526 227304 219532 227316
rect 185872 227276 219532 227304
rect 219526 227264 219532 227276
rect 219584 227264 219590 227316
rect 219986 227264 219992 227316
rect 220044 227304 220050 227316
rect 241606 227304 241612 227316
rect 220044 227276 241612 227304
rect 220044 227264 220050 227276
rect 241606 227264 241612 227276
rect 241664 227264 241670 227316
rect 249242 227264 249248 227316
rect 249300 227304 249306 227316
rect 290550 227304 290556 227316
rect 249300 227276 290556 227304
rect 249300 227264 249306 227276
rect 290550 227264 290556 227276
rect 290608 227264 290614 227316
rect 293770 227264 293776 227316
rect 293828 227304 293834 227316
rect 325326 227304 325332 227316
rect 293828 227276 325332 227304
rect 293828 227264 293834 227276
rect 325326 227264 325332 227276
rect 325384 227264 325390 227316
rect 333882 227264 333888 227316
rect 333940 227304 333946 227316
rect 356238 227304 356244 227316
rect 333940 227276 356244 227304
rect 333940 227264 333946 227276
rect 356238 227264 356244 227276
rect 356296 227264 356302 227316
rect 357250 227264 357256 227316
rect 357308 227304 357314 227316
rect 374270 227304 374276 227316
rect 357308 227276 374276 227304
rect 357308 227264 357314 227276
rect 374270 227264 374276 227276
rect 374328 227264 374334 227316
rect 382090 227264 382096 227316
rect 382148 227304 382154 227316
rect 392946 227304 392952 227316
rect 382148 227276 392952 227304
rect 382148 227264 382154 227276
rect 392946 227264 392952 227276
rect 393004 227264 393010 227316
rect 402606 227304 402612 227316
rect 393286 227276 402612 227304
rect 159692 227140 171364 227168
rect 159692 227128 159698 227140
rect 171594 227128 171600 227180
rect 171652 227168 171658 227180
rect 219802 227168 219808 227180
rect 171652 227140 219808 227168
rect 171652 227128 171658 227140
rect 219802 227128 219808 227140
rect 219860 227128 219866 227180
rect 233694 227168 233700 227180
rect 220096 227140 233700 227168
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142154 227032 142160 227044
rect 56560 227004 142160 227032
rect 56560 226992 56566 227004
rect 142154 226992 142160 227004
rect 142212 226992 142218 227044
rect 143258 226992 143264 227044
rect 143316 227032 143322 227044
rect 204070 227032 204076 227044
rect 143316 227004 204076 227032
rect 143316 226992 143322 227004
rect 204070 226992 204076 227004
rect 204128 226992 204134 227044
rect 214098 227032 214104 227044
rect 204916 227004 214104 227032
rect 122742 226856 122748 226908
rect 122800 226896 122806 226908
rect 185394 226896 185400 226908
rect 122800 226868 185400 226896
rect 122800 226856 122806 226868
rect 185394 226856 185400 226868
rect 185452 226856 185458 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 204916 226896 204944 227004
rect 214098 226992 214104 227004
rect 214156 226992 214162 227044
rect 220096 227032 220124 227140
rect 233694 227128 233700 227140
rect 233752 227128 233758 227180
rect 241146 227128 241152 227180
rect 241204 227168 241210 227180
rect 286686 227168 286692 227180
rect 241204 227140 286692 227168
rect 241204 227128 241210 227140
rect 286686 227128 286692 227140
rect 286744 227128 286750 227180
rect 306190 227128 306196 227180
rect 306248 227168 306254 227180
rect 336918 227168 336924 227180
rect 306248 227140 336924 227168
rect 306248 227128 306254 227140
rect 336918 227128 336924 227140
rect 336976 227128 336982 227180
rect 340690 227128 340696 227180
rect 340748 227168 340754 227180
rect 361390 227168 361396 227180
rect 340748 227140 361396 227168
rect 340748 227128 340754 227140
rect 361390 227128 361396 227140
rect 361448 227128 361454 227180
rect 363506 227128 363512 227180
rect 363564 227168 363570 227180
rect 368474 227168 368480 227180
rect 363564 227140 368480 227168
rect 363564 227128 363570 227140
rect 368474 227128 368480 227140
rect 368532 227128 368538 227180
rect 376662 227128 376668 227180
rect 376720 227168 376726 227180
rect 389726 227168 389732 227180
rect 376720 227140 389732 227168
rect 376720 227128 376726 227140
rect 389726 227128 389732 227140
rect 389784 227128 389790 227180
rect 393130 227128 393136 227180
rect 393188 227168 393194 227180
rect 393286 227168 393314 227276
rect 402606 227264 402612 227276
rect 402664 227264 402670 227316
rect 510614 227264 510620 227316
rect 510672 227304 510678 227316
rect 524414 227304 524420 227316
rect 510672 227276 524420 227304
rect 510672 227264 510678 227276
rect 524414 227264 524420 227276
rect 524472 227264 524478 227316
rect 526254 227264 526260 227316
rect 526312 227304 526318 227316
rect 551554 227304 551560 227316
rect 526312 227276 551560 227304
rect 526312 227264 526318 227276
rect 551554 227264 551560 227276
rect 551612 227264 551618 227316
rect 393188 227140 393314 227168
rect 393188 227128 393194 227140
rect 402238 227128 402244 227180
rect 402296 227168 402302 227180
rect 408402 227168 408408 227180
rect 402296 227140 408408 227168
rect 402296 227128 402302 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 478598 227128 478604 227180
rect 478656 227168 478662 227180
rect 486786 227168 486792 227180
rect 478656 227140 486792 227168
rect 478656 227128 478662 227140
rect 486786 227128 486792 227140
rect 486844 227128 486850 227180
rect 490374 227128 490380 227180
rect 490432 227168 490438 227180
rect 502978 227168 502984 227180
rect 490432 227140 502984 227168
rect 490432 227128 490438 227140
rect 502978 227128 502984 227140
rect 503036 227128 503042 227180
rect 505002 227128 505008 227180
rect 505060 227168 505066 227180
rect 523034 227168 523040 227180
rect 505060 227140 523040 227168
rect 505060 227128 505066 227140
rect 523034 227128 523040 227140
rect 523092 227128 523098 227180
rect 523678 227128 523684 227180
rect 523736 227168 523742 227180
rect 548334 227168 548340 227180
rect 523736 227140 548340 227168
rect 523736 227128 523742 227140
rect 548334 227128 548340 227140
rect 548392 227128 548398 227180
rect 556798 227128 556804 227180
rect 556856 227168 556862 227180
rect 570598 227168 570604 227180
rect 556856 227140 570604 227168
rect 556856 227128 556862 227140
rect 570598 227128 570604 227140
rect 570656 227128 570662 227180
rect 668578 227128 668584 227180
rect 668636 227168 668642 227180
rect 673270 227168 673276 227180
rect 668636 227140 673276 227168
rect 668636 227128 668642 227140
rect 673270 227128 673276 227140
rect 673328 227128 673334 227180
rect 214576 227004 220124 227032
rect 214576 226896 214604 227004
rect 221826 226992 221832 227044
rect 221884 227032 221890 227044
rect 271230 227032 271236 227044
rect 221884 227004 271236 227032
rect 221884 226992 221890 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 308582 227032 308588 227044
rect 271840 227004 308588 227032
rect 271840 226992 271846 227004
rect 308582 226992 308588 227004
rect 308640 226992 308646 227044
rect 310330 226992 310336 227044
rect 310388 227032 310394 227044
rect 338206 227032 338212 227044
rect 310388 227004 338212 227032
rect 310388 226992 310394 227004
rect 338206 226992 338212 227004
rect 338264 226992 338270 227044
rect 338666 226992 338672 227044
rect 338724 227032 338730 227044
rect 360102 227032 360108 227044
rect 338724 227004 360108 227032
rect 338724 226992 338730 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 362770 226992 362776 227044
rect 362828 227032 362834 227044
rect 379054 227032 379060 227044
rect 362828 227004 379060 227032
rect 362828 226992 362834 227004
rect 379054 226992 379060 227004
rect 379112 226992 379118 227044
rect 391750 226992 391756 227044
rect 391808 227032 391814 227044
rect 403526 227032 403532 227044
rect 391808 227004 403532 227032
rect 391808 226992 391814 227004
rect 403526 226992 403532 227004
rect 403584 226992 403590 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 486970 226992 486976 227044
rect 487028 227032 487034 227044
rect 500954 227032 500960 227044
rect 487028 227004 500960 227032
rect 487028 226992 487034 227004
rect 500954 226992 500960 227004
rect 501012 226992 501018 227044
rect 506290 226992 506296 227044
rect 506348 227032 506354 227044
rect 526530 227032 526536 227044
rect 506348 227004 526536 227032
rect 506348 226992 506354 227004
rect 526530 226992 526536 227004
rect 526588 226992 526594 227044
rect 533338 226992 533344 227044
rect 533396 227032 533402 227044
rect 560754 227032 560760 227044
rect 533396 227004 560760 227032
rect 533396 226992 533402 227004
rect 560754 226992 560760 227004
rect 560812 226992 560818 227044
rect 652202 226992 652208 227044
rect 652260 227032 652266 227044
rect 652260 227004 669314 227032
rect 652260 226992 652266 227004
rect 185636 226868 204944 226896
rect 209746 226868 214604 226896
rect 185636 226856 185642 226868
rect 129550 226720 129556 226772
rect 129608 226760 129614 226772
rect 197446 226760 197452 226772
rect 129608 226732 197452 226760
rect 129608 226720 129614 226732
rect 197446 226720 197452 226732
rect 197504 226720 197510 226772
rect 204714 226720 204720 226772
rect 204772 226760 204778 226772
rect 209746 226760 209774 226868
rect 214742 226856 214748 226908
rect 214800 226896 214806 226908
rect 219986 226896 219992 226908
rect 214800 226868 219992 226896
rect 214800 226856 214806 226868
rect 219986 226856 219992 226868
rect 220044 226856 220050 226908
rect 267366 226896 267372 226908
rect 229066 226868 267372 226896
rect 204772 226732 209774 226760
rect 204772 226720 204778 226732
rect 214098 226720 214104 226772
rect 214156 226760 214162 226772
rect 218422 226760 218428 226772
rect 214156 226732 218428 226760
rect 214156 226720 214162 226732
rect 218422 226720 218428 226732
rect 218480 226720 218486 226772
rect 219342 226720 219348 226772
rect 219400 226760 219406 226772
rect 229066 226760 229094 226868
rect 267366 226856 267372 226868
rect 267424 226856 267430 226908
rect 378778 226788 378784 226840
rect 378836 226828 378842 226840
rect 385862 226828 385868 226840
rect 378836 226800 385868 226828
rect 378836 226788 378842 226800
rect 385862 226788 385868 226800
rect 385920 226788 385926 226840
rect 669286 226828 669314 227004
rect 673454 226828 673460 226840
rect 669286 226800 673460 226828
rect 673454 226788 673460 226800
rect 673512 226788 673518 226840
rect 219400 226732 229094 226760
rect 219400 226720 219406 226732
rect 235810 226720 235816 226772
rect 235868 226760 235874 226772
rect 280246 226760 280252 226772
rect 235868 226732 280252 226760
rect 235868 226720 235874 226732
rect 280246 226720 280252 226732
rect 280304 226720 280310 226772
rect 136542 226584 136548 226636
rect 136600 226624 136606 226636
rect 203150 226624 203156 226636
rect 136600 226596 203156 226624
rect 136600 226584 136606 226596
rect 203150 226584 203156 226596
rect 203208 226584 203214 226636
rect 204070 226584 204076 226636
rect 204128 226624 204134 226636
rect 208118 226624 208124 226636
rect 204128 226596 208124 226624
rect 204128 226584 204134 226596
rect 208118 226584 208124 226596
rect 208176 226584 208182 226636
rect 212166 226584 212172 226636
rect 212224 226624 212230 226636
rect 214926 226624 214932 226636
rect 212224 226596 214932 226624
rect 212224 226584 212230 226596
rect 214926 226584 214932 226596
rect 214984 226584 214990 226636
rect 219526 226584 219532 226636
rect 219584 226624 219590 226636
rect 223574 226624 223580 226636
rect 219584 226596 223580 226624
rect 219584 226584 219590 226596
rect 223574 226584 223580 226596
rect 223632 226584 223638 226636
rect 225598 226584 225604 226636
rect 225656 226624 225662 226636
rect 238386 226624 238392 226636
rect 225656 226596 238392 226624
rect 225656 226584 225662 226596
rect 238386 226584 238392 226596
rect 238444 226584 238450 226636
rect 259362 226584 259368 226636
rect 259420 226624 259426 226636
rect 298278 226624 298284 226636
rect 259420 226596 298284 226624
rect 259420 226584 259426 226596
rect 298278 226584 298284 226596
rect 298336 226584 298342 226636
rect 673270 226556 673276 226568
rect 672842 226528 673276 226556
rect 673270 226516 673276 226528
rect 673328 226516 673334 226568
rect 106918 226448 106924 226500
rect 106976 226488 106982 226500
rect 146570 226488 146576 226500
rect 106976 226460 146576 226488
rect 106976 226448 106982 226460
rect 146570 226448 146576 226460
rect 146628 226448 146634 226500
rect 150066 226448 150072 226500
rect 150124 226488 150130 226500
rect 213270 226488 213276 226500
rect 150124 226460 213276 226488
rect 150124 226448 150130 226460
rect 213270 226448 213276 226460
rect 213328 226448 213334 226500
rect 216398 226448 216404 226500
rect 216456 226488 216462 226500
rect 220538 226488 220544 226500
rect 216456 226460 220544 226488
rect 216456 226448 216462 226460
rect 220538 226448 220544 226460
rect 220596 226448 220602 226500
rect 220722 226448 220728 226500
rect 220780 226488 220786 226500
rect 228910 226488 228916 226500
rect 220780 226460 228916 226488
rect 220780 226448 220786 226460
rect 228910 226448 228916 226460
rect 228968 226448 228974 226500
rect 369118 226448 369124 226500
rect 369176 226488 369182 226500
rect 376202 226488 376208 226500
rect 369176 226460 376208 226488
rect 369176 226448 369182 226460
rect 376202 226448 376208 226460
rect 376260 226448 376266 226500
rect 403986 226448 403992 226500
rect 404044 226488 404050 226500
rect 412266 226488 412272 226500
rect 404044 226460 412272 226488
rect 404044 226448 404050 226460
rect 412266 226448 412272 226460
rect 412324 226448 412330 226500
rect 474734 226448 474740 226500
rect 474792 226488 474798 226500
rect 482738 226488 482744 226500
rect 474792 226460 482744 226488
rect 474792 226448 474798 226460
rect 482738 226448 482744 226460
rect 482796 226448 482802 226500
rect 672724 226432 672776 226438
rect 386046 226380 386052 226432
rect 386104 226420 386110 226432
rect 391198 226420 391204 226432
rect 386104 226392 391204 226420
rect 386104 226380 386110 226392
rect 391198 226380 391204 226392
rect 391256 226380 391262 226432
rect 672724 226374 672776 226380
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 408678 226352 408684 226364
rect 407816 226324 408684 226352
rect 407816 226312 407822 226324
rect 408678 226312 408684 226324
rect 408736 226312 408742 226364
rect 481634 226312 481640 226364
rect 481692 226352 481698 226364
rect 487798 226352 487804 226364
rect 481692 226324 487804 226352
rect 481692 226312 481698 226324
rect 487798 226312 487804 226324
rect 487856 226312 487862 226364
rect 488074 226312 488080 226364
rect 488132 226352 488138 226364
rect 490006 226352 490012 226364
rect 488132 226324 490012 226352
rect 488132 226312 488138 226324
rect 490006 226312 490012 226324
rect 490064 226312 490070 226364
rect 122558 226244 122564 226296
rect 122616 226284 122622 226296
rect 193950 226284 193956 226296
rect 122616 226256 193956 226284
rect 122616 226244 122622 226256
rect 193950 226244 193956 226256
rect 194008 226244 194014 226296
rect 194134 226244 194140 226296
rect 194192 226284 194198 226296
rect 204898 226284 204904 226296
rect 194192 226256 204904 226284
rect 194192 226244 194198 226256
rect 204898 226244 204904 226256
rect 204956 226244 204962 226296
rect 205082 226244 205088 226296
rect 205140 226284 205146 226296
rect 254486 226284 254492 226296
rect 205140 226256 254492 226284
rect 205140 226244 205146 226256
rect 254486 226244 254492 226256
rect 254544 226244 254550 226296
rect 260650 226244 260656 226296
rect 260708 226284 260714 226296
rect 298922 226284 298928 226296
rect 260708 226256 298928 226284
rect 260708 226244 260714 226256
rect 298922 226244 298928 226256
rect 298980 226244 298986 226296
rect 308858 226244 308864 226296
rect 308916 226284 308922 226296
rect 336274 226284 336280 226296
rect 308916 226256 336280 226284
rect 308916 226244 308922 226256
rect 336274 226244 336280 226256
rect 336332 226244 336338 226296
rect 388622 226244 388628 226296
rect 388680 226284 388686 226296
rect 394234 226284 394240 226296
rect 388680 226256 394240 226284
rect 388680 226244 388686 226256
rect 394234 226244 394240 226256
rect 394292 226244 394298 226296
rect 539962 226284 539968 226296
rect 528526 226256 539968 226284
rect 72418 226108 72424 226160
rect 72476 226148 72482 226160
rect 141142 226148 141148 226160
rect 72476 226120 141148 226148
rect 72476 226108 72482 226120
rect 141142 226108 141148 226120
rect 141200 226108 141206 226160
rect 141510 226108 141516 226160
rect 141568 226148 141574 226160
rect 145006 226148 145012 226160
rect 141568 226120 145012 226148
rect 141568 226108 141574 226120
rect 145006 226108 145012 226120
rect 145064 226108 145070 226160
rect 145190 226108 145196 226160
rect 145248 226148 145254 226160
rect 146754 226148 146760 226160
rect 145248 226120 146760 226148
rect 145248 226108 145254 226120
rect 146754 226108 146760 226120
rect 146812 226108 146818 226160
rect 148962 226108 148968 226160
rect 149020 226148 149026 226160
rect 213454 226148 213460 226160
rect 149020 226120 213460 226148
rect 149020 226108 149026 226120
rect 213454 226108 213460 226120
rect 213512 226108 213518 226160
rect 213638 226108 213644 226160
rect 213696 226148 213702 226160
rect 219986 226148 219992 226160
rect 213696 226120 219992 226148
rect 213696 226108 213702 226120
rect 219986 226108 219992 226120
rect 220044 226108 220050 226160
rect 222010 226108 222016 226160
rect 222068 226148 222074 226160
rect 269942 226148 269948 226160
rect 222068 226120 269948 226148
rect 222068 226108 222074 226120
rect 269942 226108 269948 226120
rect 270000 226108 270006 226160
rect 270218 226108 270224 226160
rect 270276 226148 270282 226160
rect 287514 226148 287520 226160
rect 270276 226120 287520 226148
rect 270276 226108 270282 226120
rect 287514 226108 287520 226120
rect 287572 226108 287578 226160
rect 288066 226108 288072 226160
rect 288124 226148 288130 226160
rect 322750 226148 322756 226160
rect 288124 226120 322756 226148
rect 288124 226108 288130 226120
rect 322750 226108 322756 226120
rect 322808 226108 322814 226160
rect 525978 226108 525984 226160
rect 526036 226148 526042 226160
rect 528526 226148 528554 226256
rect 539962 226244 539968 226256
rect 540020 226244 540026 226296
rect 563698 226244 563704 226296
rect 563756 226284 563762 226296
rect 568114 226284 568120 226296
rect 563756 226256 568120 226284
rect 563756 226244 563762 226256
rect 568114 226244 568120 226256
rect 568172 226244 568178 226296
rect 672604 226160 672656 226166
rect 538490 226148 538496 226160
rect 526036 226120 528554 226148
rect 538186 226120 538496 226148
rect 526036 226108 526042 226120
rect 83458 225972 83464 226024
rect 83516 226012 83522 226024
rect 163038 226012 163044 226024
rect 83516 225984 163044 226012
rect 83516 225972 83522 225984
rect 163038 225972 163044 225984
rect 163096 225972 163102 226024
rect 196618 225972 196624 226024
rect 196676 226012 196682 226024
rect 236454 226012 236460 226024
rect 196676 225984 236460 226012
rect 196676 225972 196682 225984
rect 236454 225972 236460 225984
rect 236512 225972 236518 226024
rect 252462 225972 252468 226024
rect 252520 226012 252526 226024
rect 293126 226012 293132 226024
rect 252520 225984 293132 226012
rect 252520 225972 252526 225984
rect 293126 225972 293132 225984
rect 293184 225972 293190 226024
rect 299382 225972 299388 226024
rect 299440 226012 299446 226024
rect 328546 226012 328552 226024
rect 299440 225984 328552 226012
rect 299440 225972 299446 225984
rect 328546 225972 328552 225984
rect 328604 225972 328610 226024
rect 335170 225972 335176 226024
rect 335228 226012 335234 226024
rect 356882 226012 356888 226024
rect 335228 225984 356888 226012
rect 335228 225972 335234 225984
rect 356882 225972 356888 225984
rect 356940 225972 356946 226024
rect 361206 225972 361212 226024
rect 361264 226012 361270 226024
rect 377490 226012 377496 226024
rect 361264 225984 377496 226012
rect 361264 225972 361270 225984
rect 377490 225972 377496 225984
rect 377548 225972 377554 226024
rect 498102 225972 498108 226024
rect 498160 226012 498166 226024
rect 514294 226012 514300 226024
rect 498160 225984 514300 226012
rect 498160 225972 498166 225984
rect 514294 225972 514300 225984
rect 514352 225972 514358 226024
rect 516594 225972 516600 226024
rect 516652 226012 516658 226024
rect 538186 226012 538214 226120
rect 538490 226108 538496 226120
rect 538548 226108 538554 226160
rect 672604 226102 672656 226108
rect 672074 226040 672080 226092
rect 672132 226080 672138 226092
rect 672132 226052 672520 226080
rect 672132 226040 672138 226052
rect 516652 225984 538214 226012
rect 516652 225972 516658 225984
rect 538306 225972 538312 226024
rect 538364 226012 538370 226024
rect 557258 226012 557264 226024
rect 538364 225984 557264 226012
rect 538364 225972 538370 225984
rect 557258 225972 557264 225984
rect 557316 225972 557322 226024
rect 76558 225836 76564 225888
rect 76616 225876 76622 225888
rect 158254 225876 158260 225888
rect 76616 225848 158260 225876
rect 76616 225836 76622 225848
rect 158254 225836 158260 225848
rect 158312 225836 158318 225888
rect 169662 225836 169668 225888
rect 169720 225876 169726 225888
rect 171594 225876 171600 225888
rect 169720 225848 171600 225876
rect 169720 225836 169726 225848
rect 171594 225836 171600 225848
rect 171652 225836 171658 225888
rect 171778 225836 171784 225888
rect 171836 225876 171842 225888
rect 204530 225876 204536 225888
rect 171836 225848 204536 225876
rect 171836 225836 171842 225848
rect 204530 225836 204536 225848
rect 204588 225836 204594 225888
rect 204898 225836 204904 225888
rect 204956 225876 204962 225888
rect 213638 225876 213644 225888
rect 204956 225848 213644 225876
rect 204956 225836 204962 225848
rect 213638 225836 213644 225848
rect 213696 225836 213702 225888
rect 219986 225836 219992 225888
rect 220044 225876 220050 225888
rect 244182 225876 244188 225888
rect 220044 225848 244188 225876
rect 220044 225836 220050 225848
rect 244182 225836 244188 225848
rect 244240 225836 244246 225888
rect 261846 225836 261852 225888
rect 261904 225876 261910 225888
rect 300854 225876 300860 225888
rect 261904 225848 300860 225876
rect 261904 225836 261910 225848
rect 300854 225836 300860 225848
rect 300912 225836 300918 225888
rect 312906 225836 312912 225888
rect 312964 225876 312970 225888
rect 341702 225876 341708 225888
rect 312964 225848 341708 225876
rect 312964 225836 312970 225848
rect 341702 225836 341708 225848
rect 341760 225836 341766 225888
rect 341978 225836 341984 225888
rect 342036 225876 342042 225888
rect 365254 225876 365260 225888
rect 342036 225848 365260 225876
rect 342036 225836 342042 225848
rect 365254 225836 365260 225848
rect 365312 225836 365318 225888
rect 375006 225836 375012 225888
rect 375064 225876 375070 225888
rect 387794 225876 387800 225888
rect 375064 225848 387800 225876
rect 375064 225836 375070 225848
rect 387794 225836 387800 225848
rect 387852 225836 387858 225888
rect 394326 225836 394332 225888
rect 394384 225876 394390 225888
rect 403250 225876 403256 225888
rect 394384 225848 403256 225876
rect 394384 225836 394390 225848
rect 403250 225836 403256 225848
rect 403308 225836 403314 225888
rect 501138 225836 501144 225888
rect 501196 225876 501202 225888
rect 519170 225876 519176 225888
rect 501196 225848 519176 225876
rect 501196 225836 501202 225848
rect 519170 225836 519176 225848
rect 519228 225836 519234 225888
rect 521746 225836 521752 225888
rect 521804 225876 521810 225888
rect 545758 225876 545764 225888
rect 521804 225848 545764 225876
rect 521804 225836 521810 225848
rect 545758 225836 545764 225848
rect 545816 225836 545822 225888
rect 672258 225836 672264 225888
rect 672316 225876 672322 225888
rect 672316 225848 672406 225876
rect 672316 225836 672322 225848
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462958 225808 462964 225820
rect 458692 225780 462964 225808
rect 458692 225768 458698 225780
rect 462958 225768 462964 225780
rect 463016 225768 463022 225820
rect 66162 225700 66168 225752
rect 66220 225740 66226 225752
rect 149790 225740 149796 225752
rect 66220 225712 149796 225740
rect 66220 225700 66226 225712
rect 149790 225700 149796 225712
rect 149848 225700 149854 225752
rect 151262 225700 151268 225752
rect 151320 225740 151326 225752
rect 151320 225712 203380 225740
rect 151320 225700 151326 225712
rect 58986 225564 58992 225616
rect 59044 225604 59050 225616
rect 141510 225604 141516 225616
rect 59044 225576 141516 225604
rect 59044 225564 59050 225576
rect 141510 225564 141516 225576
rect 141568 225564 141574 225616
rect 141786 225564 141792 225616
rect 141844 225604 141850 225616
rect 203150 225604 203156 225616
rect 141844 225576 203156 225604
rect 141844 225564 141850 225576
rect 203150 225564 203156 225576
rect 203208 225564 203214 225616
rect 203352 225604 203380 225712
rect 204898 225700 204904 225752
rect 204956 225740 204962 225752
rect 248874 225740 248880 225752
rect 204956 225712 248880 225740
rect 204956 225700 204962 225712
rect 248874 225700 248880 225712
rect 248932 225700 248938 225752
rect 251082 225700 251088 225752
rect 251140 225740 251146 225752
rect 294414 225740 294420 225752
rect 251140 225712 294420 225740
rect 251140 225700 251146 225712
rect 294414 225700 294420 225712
rect 294472 225700 294478 225752
rect 296438 225700 296444 225752
rect 296496 225740 296502 225752
rect 327902 225740 327908 225752
rect 296496 225712 327908 225740
rect 296496 225700 296502 225712
rect 327902 225700 327908 225712
rect 327960 225700 327966 225752
rect 329742 225700 329748 225752
rect 329800 225740 329806 225752
rect 353662 225740 353668 225752
rect 329800 225712 353668 225740
rect 329800 225700 329806 225712
rect 353662 225700 353668 225712
rect 353720 225700 353726 225752
rect 365346 225700 365352 225752
rect 365404 225740 365410 225752
rect 383286 225740 383292 225752
rect 365404 225712 383292 225740
rect 365404 225700 365410 225712
rect 383286 225700 383292 225712
rect 383344 225700 383350 225752
rect 387702 225700 387708 225752
rect 387760 225740 387766 225752
rect 397822 225740 397828 225752
rect 387760 225712 397828 225740
rect 387760 225700 387766 225712
rect 397822 225700 397828 225712
rect 397880 225700 397886 225752
rect 481174 225700 481180 225752
rect 481232 225740 481238 225752
rect 492674 225740 492680 225752
rect 481232 225712 492680 225740
rect 481232 225700 481238 225712
rect 492674 225700 492680 225712
rect 492732 225700 492738 225752
rect 493686 225700 493692 225752
rect 493744 225740 493750 225752
rect 505370 225740 505376 225752
rect 493744 225712 505376 225740
rect 493744 225700 493750 225712
rect 505370 225700 505376 225712
rect 505428 225700 505434 225752
rect 508866 225700 508872 225752
rect 508924 225740 508930 225752
rect 529198 225740 529204 225752
rect 508924 225712 529204 225740
rect 508924 225700 508930 225712
rect 529198 225700 529204 225712
rect 529256 225700 529262 225752
rect 535914 225700 535920 225752
rect 535972 225740 535978 225752
rect 563054 225740 563060 225752
rect 535972 225712 563060 225740
rect 535972 225700 535978 225712
rect 563054 225700 563060 225712
rect 563112 225700 563118 225752
rect 672264 225684 672316 225690
rect 672264 225626 672316 225632
rect 217134 225604 217140 225616
rect 203352 225576 217140 225604
rect 217134 225564 217140 225576
rect 217192 225564 217198 225616
rect 217870 225564 217876 225616
rect 217928 225604 217934 225616
rect 266078 225604 266084 225616
rect 217928 225576 266084 225604
rect 217928 225564 217934 225576
rect 266078 225564 266084 225576
rect 266136 225564 266142 225616
rect 266998 225564 267004 225616
rect 267056 225604 267062 225616
rect 274450 225604 274456 225616
rect 267056 225576 274456 225604
rect 267056 225564 267062 225576
rect 274450 225564 274456 225576
rect 274508 225564 274514 225616
rect 278406 225564 278412 225616
rect 278464 225604 278470 225616
rect 313274 225604 313280 225616
rect 278464 225576 313280 225604
rect 278464 225564 278470 225576
rect 313274 225564 313280 225576
rect 313332 225564 313338 225616
rect 327718 225564 327724 225616
rect 327776 225604 327782 225616
rect 352374 225604 352380 225616
rect 327776 225576 352380 225604
rect 327776 225564 327782 225576
rect 352374 225564 352380 225576
rect 352432 225564 352438 225616
rect 352926 225564 352932 225616
rect 352984 225604 352990 225616
rect 371602 225604 371608 225616
rect 352984 225576 371608 225604
rect 352984 225564 352990 225576
rect 371602 225564 371608 225576
rect 371660 225564 371666 225616
rect 382918 225564 382924 225616
rect 382976 225604 382982 225616
rect 396166 225604 396172 225616
rect 382976 225576 396172 225604
rect 382976 225564 382982 225576
rect 396166 225564 396172 225576
rect 396224 225564 396230 225616
rect 410978 225564 410984 225616
rect 411036 225604 411042 225616
rect 416130 225604 416136 225616
rect 411036 225576 416136 225604
rect 411036 225564 411042 225576
rect 416130 225564 416136 225576
rect 416188 225564 416194 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 488718 225604 488724 225616
rect 477368 225576 488724 225604
rect 477368 225564 477374 225576
rect 488718 225564 488724 225576
rect 488776 225564 488782 225616
rect 489362 225564 489368 225616
rect 489420 225604 489426 225616
rect 503162 225604 503168 225616
rect 489420 225576 503168 225604
rect 489420 225564 489426 225576
rect 503162 225564 503168 225576
rect 503220 225564 503226 225616
rect 510154 225564 510160 225616
rect 510212 225604 510218 225616
rect 530578 225604 530584 225616
rect 510212 225576 530584 225604
rect 510212 225564 510218 225576
rect 530578 225564 530584 225576
rect 530636 225564 530642 225616
rect 531406 225564 531412 225616
rect 531464 225604 531470 225616
rect 558178 225604 558184 225616
rect 531464 225576 558184 225604
rect 531464 225564 531470 225576
rect 558178 225564 558184 225576
rect 558236 225564 558242 225616
rect 125226 225428 125232 225480
rect 125284 225468 125290 225480
rect 196158 225468 196164 225480
rect 125284 225440 196164 225468
rect 125284 225428 125290 225440
rect 196158 225428 196164 225440
rect 196216 225428 196222 225480
rect 197998 225428 198004 225480
rect 198056 225468 198062 225480
rect 204898 225468 204904 225480
rect 198056 225440 204904 225468
rect 198056 225428 198062 225440
rect 204898 225428 204904 225440
rect 204956 225428 204962 225480
rect 209590 225428 209596 225480
rect 209648 225468 209654 225480
rect 259638 225468 259644 225480
rect 209648 225440 259644 225468
rect 209648 225428 209654 225440
rect 259638 225428 259644 225440
rect 259696 225428 259702 225480
rect 297358 225428 297364 225480
rect 297416 225468 297422 225480
rect 310514 225468 310520 225480
rect 297416 225440 310520 225468
rect 297416 225428 297422 225440
rect 310514 225428 310520 225440
rect 310572 225428 310578 225480
rect 671890 225428 671896 225480
rect 671948 225468 671954 225480
rect 671948 225440 672182 225468
rect 671948 225428 671954 225440
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 129366 225292 129372 225344
rect 129424 225332 129430 225344
rect 199102 225332 199108 225344
rect 129424 225304 199108 225332
rect 129424 225292 129430 225304
rect 199102 225292 199108 225304
rect 199160 225292 199166 225344
rect 203150 225292 203156 225344
rect 203208 225332 203214 225344
rect 209406 225332 209412 225344
rect 203208 225304 209412 225332
rect 203208 225292 203214 225304
rect 209406 225292 209412 225304
rect 209464 225292 209470 225344
rect 222930 225332 222936 225344
rect 209746 225304 222936 225332
rect 62022 225156 62028 225208
rect 62080 225196 62086 225208
rect 130378 225196 130384 225208
rect 62080 225168 130384 225196
rect 62080 225156 62086 225168
rect 130378 225156 130384 225168
rect 130436 225156 130442 225208
rect 135070 225156 135076 225208
rect 135128 225196 135134 225208
rect 204254 225196 204260 225208
rect 135128 225168 204260 225196
rect 135128 225156 135134 225168
rect 204254 225156 204260 225168
rect 204312 225156 204318 225208
rect 204530 225156 204536 225208
rect 204588 225196 204594 225208
rect 209746 225196 209774 225304
rect 222930 225292 222936 225304
rect 222988 225292 222994 225344
rect 242894 225292 242900 225344
rect 242952 225332 242958 225344
rect 285030 225332 285036 225344
rect 242952 225304 285036 225332
rect 242952 225292 242958 225304
rect 285030 225292 285036 225304
rect 285088 225292 285094 225344
rect 204588 225168 209774 225196
rect 204588 225156 204594 225168
rect 215202 225156 215208 225208
rect 215260 225196 215266 225208
rect 217870 225196 217876 225208
rect 215260 225168 217876 225196
rect 215260 225156 215266 225168
rect 217870 225156 217876 225168
rect 217928 225156 217934 225208
rect 426434 225156 426440 225208
rect 426492 225196 426498 225208
rect 426986 225196 426992 225208
rect 426492 225168 426992 225196
rect 426492 225156 426498 225168
rect 426986 225156 426992 225168
rect 427044 225156 427050 225208
rect 666462 225156 666468 225208
rect 666520 225196 666526 225208
rect 666520 225168 669314 225196
rect 666520 225156 666526 225168
rect 132402 225020 132408 225072
rect 132460 225060 132466 225072
rect 201678 225060 201684 225072
rect 132460 225032 201684 225060
rect 132460 225020 132466 225032
rect 201678 225020 201684 225032
rect 201736 225020 201742 225072
rect 203886 225020 203892 225072
rect 203944 225060 203950 225072
rect 255130 225060 255136 225072
rect 203944 225032 255136 225060
rect 203944 225020 203950 225032
rect 255130 225020 255136 225032
rect 255188 225020 255194 225072
rect 669286 225060 669314 225168
rect 672034 225140 672086 225146
rect 672034 225082 672086 225088
rect 669286 225032 671968 225060
rect 355226 224952 355232 225004
rect 355284 224992 355290 225004
rect 358170 224992 358176 225004
rect 355284 224964 358176 224992
rect 355284 224952 355290 224964
rect 358170 224952 358176 224964
rect 358228 224952 358234 225004
rect 404170 224952 404176 225004
rect 404228 224992 404234 225004
rect 410610 224992 410616 225004
rect 404228 224964 410616 224992
rect 404228 224952 404234 224964
rect 410610 224952 410616 224964
rect 410668 224952 410674 225004
rect 416498 224952 416504 225004
rect 416556 224992 416562 225004
rect 422202 224992 422208 225004
rect 416556 224964 422208 224992
rect 416556 224952 416562 224964
rect 422202 224952 422208 224964
rect 422260 224952 422266 225004
rect 96246 224884 96252 224936
rect 96304 224924 96310 224936
rect 172974 224924 172980 224936
rect 96304 224896 172980 224924
rect 96304 224884 96310 224896
rect 172974 224884 172980 224896
rect 173032 224884 173038 224936
rect 173176 224896 176700 224924
rect 89438 224748 89444 224800
rect 89496 224788 89502 224800
rect 168190 224788 168196 224800
rect 89496 224760 168196 224788
rect 89496 224748 89502 224760
rect 168190 224748 168196 224760
rect 168248 224748 168254 224800
rect 171962 224748 171968 224800
rect 172020 224788 172026 224800
rect 173176 224788 173204 224896
rect 172020 224760 173204 224788
rect 176672 224788 176700 224896
rect 177482 224884 177488 224936
rect 177540 224924 177546 224936
rect 199746 224924 199752 224936
rect 177540 224896 199752 224924
rect 177540 224884 177546 224896
rect 199746 224884 199752 224896
rect 199804 224884 199810 224936
rect 199930 224884 199936 224936
rect 199988 224924 199994 224936
rect 248046 224924 248052 224936
rect 199988 224896 248052 224924
rect 199988 224884 199994 224896
rect 248046 224884 248052 224896
rect 248104 224884 248110 224936
rect 272518 224884 272524 224936
rect 272576 224924 272582 224936
rect 309870 224924 309876 224936
rect 272576 224896 309876 224924
rect 272576 224884 272582 224896
rect 309870 224884 309876 224896
rect 309928 224884 309934 224936
rect 319806 224884 319812 224936
rect 319864 224924 319870 224936
rect 345934 224924 345940 224936
rect 319864 224896 345940 224924
rect 319864 224884 319870 224896
rect 345934 224884 345940 224896
rect 345992 224884 345998 224936
rect 519354 224884 519360 224936
rect 519412 224924 519418 224936
rect 534994 224924 535000 224936
rect 519412 224896 535000 224924
rect 519412 224884 519418 224896
rect 534994 224884 535000 224896
rect 535052 224924 535058 224936
rect 621014 224924 621020 224936
rect 535052 224896 621020 224924
rect 535052 224884 535058 224896
rect 621014 224884 621020 224896
rect 621072 224884 621078 224936
rect 232590 224788 232596 224800
rect 176672 224760 232596 224788
rect 172020 224748 172026 224760
rect 232590 224748 232596 224760
rect 232648 224748 232654 224800
rect 245470 224748 245476 224800
rect 245528 224788 245534 224800
rect 287698 224788 287704 224800
rect 245528 224760 287704 224788
rect 245528 224748 245534 224760
rect 287698 224748 287704 224760
rect 287756 224748 287762 224800
rect 311526 224748 311532 224800
rect 311584 224788 311590 224800
rect 338850 224788 338856 224800
rect 311584 224760 338856 224788
rect 311584 224748 311590 224760
rect 338850 224748 338856 224760
rect 338908 224748 338914 224800
rect 462498 224748 462504 224800
rect 462556 224788 462562 224800
rect 469306 224788 469312 224800
rect 462556 224760 469312 224788
rect 462556 224748 462562 224760
rect 469306 224748 469312 224760
rect 469364 224748 469370 224800
rect 506934 224748 506940 224800
rect 506992 224788 506998 224800
rect 526346 224788 526352 224800
rect 506992 224760 526352 224788
rect 506992 224748 506998 224760
rect 526346 224748 526352 224760
rect 526404 224748 526410 224800
rect 529934 224748 529940 224800
rect 529992 224788 529998 224800
rect 529992 224760 549024 224788
rect 529992 224748 529998 224760
rect 350350 224680 350356 224732
rect 350408 224720 350414 224732
rect 354950 224720 354956 224732
rect 350408 224692 354956 224720
rect 350408 224680 350414 224692
rect 354950 224680 354956 224692
rect 355008 224680 355014 224732
rect 79962 224612 79968 224664
rect 80020 224652 80026 224664
rect 160462 224652 160468 224664
rect 80020 224624 160468 224652
rect 80020 224612 80026 224624
rect 160462 224612 160468 224624
rect 160520 224612 160526 224664
rect 165154 224612 165160 224664
rect 165212 224652 165218 224664
rect 227438 224652 227444 224664
rect 165212 224624 227444 224652
rect 165212 224612 165218 224624
rect 227438 224612 227444 224624
rect 227496 224612 227502 224664
rect 228726 224612 228732 224664
rect 228784 224652 228790 224664
rect 274910 224652 274916 224664
rect 228784 224624 274916 224652
rect 228784 224612 228790 224624
rect 274910 224612 274916 224624
rect 274968 224612 274974 224664
rect 275094 224612 275100 224664
rect 275152 224652 275158 224664
rect 311158 224652 311164 224664
rect 275152 224624 311164 224652
rect 275152 224612 275158 224624
rect 311158 224612 311164 224624
rect 311216 224612 311222 224664
rect 322842 224612 322848 224664
rect 322900 224652 322906 224664
rect 349798 224652 349804 224664
rect 322900 224624 349804 224652
rect 322900 224612 322906 224624
rect 349798 224612 349804 224624
rect 349856 224612 349862 224664
rect 359458 224612 359464 224664
rect 359516 224652 359522 224664
rect 378134 224652 378140 224664
rect 359516 224624 378140 224652
rect 359516 224612 359522 224624
rect 378134 224612 378140 224624
rect 378192 224612 378198 224664
rect 494054 224612 494060 224664
rect 494112 224652 494118 224664
rect 510154 224652 510160 224664
rect 494112 224624 510160 224652
rect 494112 224612 494118 224624
rect 510154 224612 510160 224624
rect 510212 224612 510218 224664
rect 520458 224612 520464 224664
rect 520516 224652 520522 224664
rect 544378 224652 544384 224664
rect 520516 224624 544384 224652
rect 520516 224612 520522 224624
rect 544378 224612 544384 224624
rect 544436 224612 544442 224664
rect 548996 224652 549024 224760
rect 549254 224748 549260 224800
rect 549312 224788 549318 224800
rect 557074 224788 557080 224800
rect 549312 224760 557080 224788
rect 549312 224748 549318 224760
rect 557074 224748 557080 224760
rect 557132 224748 557138 224800
rect 557258 224748 557264 224800
rect 557316 224788 557322 224800
rect 626534 224788 626540 224800
rect 557316 224760 626540 224788
rect 557316 224748 557322 224760
rect 626534 224748 626540 224760
rect 626592 224748 626598 224800
rect 671820 224732 671872 224738
rect 671820 224674 671872 224680
rect 549990 224652 549996 224664
rect 548996 224624 549996 224652
rect 549990 224612 549996 224624
rect 550048 224652 550054 224664
rect 625246 224652 625252 224664
rect 550048 224624 625252 224652
rect 550048 224612 550054 224624
rect 625246 224612 625252 224624
rect 625304 224612 625310 224664
rect 668026 224612 668032 224664
rect 668084 224652 668090 224664
rect 668084 224624 671738 224652
rect 668084 224612 668090 224624
rect 85482 224476 85488 224528
rect 85540 224516 85546 224528
rect 165614 224516 165620 224528
rect 85540 224488 165620 224516
rect 85540 224476 85546 224488
rect 165614 224476 165620 224488
rect 165672 224476 165678 224528
rect 165982 224476 165988 224528
rect 166040 224516 166046 224528
rect 185394 224516 185400 224528
rect 166040 224488 185400 224516
rect 166040 224476 166046 224488
rect 185394 224476 185400 224488
rect 185452 224476 185458 224528
rect 185578 224476 185584 224528
rect 185636 224516 185642 224528
rect 237742 224516 237748 224528
rect 185636 224488 237748 224516
rect 185636 224476 185642 224488
rect 237742 224476 237748 224488
rect 237800 224476 237806 224528
rect 248322 224476 248328 224528
rect 248380 224516 248386 224528
rect 291838 224516 291844 224528
rect 248380 224488 291844 224516
rect 248380 224476 248386 224488
rect 291838 224476 291844 224488
rect 291896 224476 291902 224528
rect 294874 224476 294880 224528
rect 294932 224516 294938 224528
rect 325970 224516 325976 224528
rect 294932 224488 325976 224516
rect 294932 224476 294938 224488
rect 325970 224476 325976 224488
rect 326028 224476 326034 224528
rect 331858 224476 331864 224528
rect 331916 224516 331922 224528
rect 337562 224516 337568 224528
rect 331916 224488 337568 224516
rect 331916 224476 331922 224488
rect 337562 224476 337568 224488
rect 337620 224476 337626 224528
rect 346302 224476 346308 224528
rect 346360 224516 346366 224528
rect 366542 224516 366548 224528
rect 346360 224488 366548 224516
rect 346360 224476 346366 224488
rect 366542 224476 366548 224488
rect 366600 224476 366606 224528
rect 379238 224476 379244 224528
rect 379296 224516 379302 224528
rect 393590 224516 393596 224528
rect 379296 224488 393596 224516
rect 379296 224476 379302 224488
rect 393590 224476 393596 224488
rect 393648 224476 393654 224528
rect 447502 224476 447508 224528
rect 447560 224516 447566 224528
rect 448054 224516 448060 224528
rect 447560 224488 448060 224516
rect 447560 224476 447566 224488
rect 448054 224476 448060 224488
rect 448112 224476 448118 224528
rect 456058 224476 456064 224528
rect 456116 224516 456122 224528
rect 459738 224516 459744 224528
rect 456116 224488 459744 224516
rect 456116 224476 456122 224488
rect 459738 224476 459744 224488
rect 459796 224476 459802 224528
rect 491294 224476 491300 224528
rect 491352 224516 491358 224528
rect 506014 224516 506020 224528
rect 491352 224488 506020 224516
rect 491352 224476 491358 224488
rect 506014 224476 506020 224488
rect 506072 224476 506078 224528
rect 515950 224476 515956 224528
rect 516008 224516 516014 224528
rect 538950 224516 538956 224528
rect 516008 224488 538956 224516
rect 516008 224476 516014 224488
rect 538950 224476 538956 224488
rect 539008 224476 539014 224528
rect 542446 224476 542452 224528
rect 542504 224516 542510 224528
rect 542814 224516 542820 224528
rect 542504 224488 542820 224516
rect 542504 224476 542510 224488
rect 542814 224476 542820 224488
rect 542872 224516 542878 224528
rect 623222 224516 623228 224528
rect 542872 224488 623228 224516
rect 542872 224476 542878 224488
rect 623222 224476 623228 224488
rect 623280 224476 623286 224528
rect 671246 224408 671252 224460
rect 671304 224448 671310 224460
rect 671304 224420 671622 224448
rect 671304 224408 671310 224420
rect 73706 224340 73712 224392
rect 73764 224380 73770 224392
rect 155310 224380 155316 224392
rect 73764 224352 155316 224380
rect 73764 224340 73770 224352
rect 155310 224340 155316 224352
rect 155368 224340 155374 224392
rect 155862 224340 155868 224392
rect 155920 224380 155926 224392
rect 159634 224380 159640 224392
rect 155920 224352 159640 224380
rect 155920 224340 155926 224352
rect 159634 224340 159640 224352
rect 159692 224340 159698 224392
rect 161658 224340 161664 224392
rect 161716 224380 161722 224392
rect 224862 224380 224868 224392
rect 161716 224352 224868 224380
rect 161716 224340 161722 224352
rect 224862 224340 224868 224352
rect 224920 224340 224926 224392
rect 233142 224340 233148 224392
rect 233200 224380 233206 224392
rect 277670 224380 277676 224392
rect 233200 224352 277676 224380
rect 233200 224340 233206 224352
rect 277670 224340 277676 224352
rect 277728 224340 277734 224392
rect 289630 224340 289636 224392
rect 289688 224380 289694 224392
rect 296990 224380 296996 224392
rect 289688 224352 296996 224380
rect 289688 224340 289694 224352
rect 296990 224340 296996 224352
rect 297048 224340 297054 224392
rect 299106 224340 299112 224392
rect 299164 224380 299170 224392
rect 331398 224380 331404 224392
rect 299164 224352 331404 224380
rect 299164 224340 299170 224352
rect 331398 224340 331404 224352
rect 331456 224340 331462 224392
rect 342162 224340 342168 224392
rect 342220 224380 342226 224392
rect 362034 224380 362040 224392
rect 342220 224352 362040 224380
rect 342220 224340 342226 224352
rect 362034 224340 362040 224352
rect 362092 224340 362098 224392
rect 366726 224340 366732 224392
rect 366784 224380 366790 224392
rect 381630 224380 381636 224392
rect 366784 224352 381636 224380
rect 366784 224340 366790 224352
rect 381630 224340 381636 224352
rect 381688 224340 381694 224392
rect 394510 224340 394516 224392
rect 394568 224380 394574 224392
rect 404538 224380 404544 224392
rect 394568 224352 404544 224380
rect 394568 224340 394574 224352
rect 404538 224340 404544 224352
rect 404596 224340 404602 224392
rect 480530 224340 480536 224392
rect 480588 224380 480594 224392
rect 492858 224380 492864 224392
rect 480588 224352 492864 224380
rect 480588 224340 480594 224352
rect 492858 224340 492864 224352
rect 492916 224340 492922 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516778 224380 516784 224392
rect 499264 224352 516784 224380
rect 499264 224340 499270 224352
rect 516778 224340 516784 224352
rect 516836 224340 516842 224392
rect 525610 224340 525616 224392
rect 525668 224380 525674 224392
rect 550634 224380 550640 224392
rect 525668 224352 550640 224380
rect 525668 224340 525674 224352
rect 550634 224340 550640 224352
rect 550692 224340 550698 224392
rect 625982 224380 625988 224392
rect 558012 224352 625988 224380
rect 554958 224272 554964 224324
rect 555016 224312 555022 224324
rect 555878 224312 555884 224324
rect 555016 224284 555884 224312
rect 555016 224272 555022 224284
rect 555878 224272 555884 224284
rect 555936 224312 555942 224324
rect 558012 224312 558040 224352
rect 625982 224340 625988 224352
rect 626040 224340 626046 224392
rect 555936 224284 558040 224312
rect 555936 224272 555942 224284
rect 68922 224204 68928 224256
rect 68980 224244 68986 224256
rect 152734 224244 152740 224256
rect 68980 224216 152740 224244
rect 68980 224204 68986 224216
rect 152734 224204 152740 224216
rect 152792 224204 152798 224256
rect 168006 224204 168012 224256
rect 168064 224244 168070 224256
rect 230014 224244 230020 224256
rect 168064 224216 230020 224244
rect 168064 224204 168070 224216
rect 230014 224204 230020 224216
rect 230072 224204 230078 224256
rect 231670 224204 231676 224256
rect 231728 224244 231734 224256
rect 278958 224244 278964 224256
rect 231728 224216 278964 224244
rect 231728 224204 231734 224216
rect 278958 224204 278964 224216
rect 279016 224204 279022 224256
rect 286318 224204 286324 224256
rect 286376 224244 286382 224256
rect 289906 224244 289912 224256
rect 286376 224216 289912 224244
rect 286376 224204 286382 224216
rect 289906 224204 289912 224216
rect 289964 224204 289970 224256
rect 290826 224204 290832 224256
rect 290884 224244 290890 224256
rect 324038 224244 324044 224256
rect 290884 224216 324044 224244
rect 290884 224204 290890 224216
rect 324038 224204 324044 224216
rect 324096 224204 324102 224256
rect 339402 224204 339408 224256
rect 339460 224244 339466 224256
rect 362310 224244 362316 224256
rect 339460 224216 362316 224244
rect 339460 224204 339466 224216
rect 362310 224204 362316 224216
rect 362368 224204 362374 224256
rect 372522 224204 372528 224256
rect 372580 224244 372586 224256
rect 387426 224244 387432 224256
rect 372580 224216 387432 224244
rect 372580 224204 372586 224216
rect 387426 224204 387432 224216
rect 387484 224204 387490 224256
rect 390186 224204 390192 224256
rect 390244 224244 390250 224256
rect 401962 224244 401968 224256
rect 390244 224216 401968 224244
rect 390244 224204 390250 224216
rect 401962 224204 401968 224216
rect 402020 224204 402026 224256
rect 405550 224204 405556 224256
rect 405608 224244 405614 224256
rect 414198 224244 414204 224256
rect 405608 224216 414204 224244
rect 405608 224204 405614 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 470226 224204 470232 224256
rect 470284 224244 470290 224256
rect 480346 224244 480352 224256
rect 470284 224216 480352 224244
rect 470284 224204 470290 224216
rect 480346 224204 480352 224216
rect 480404 224204 480410 224256
rect 483750 224204 483756 224256
rect 483808 224244 483814 224256
rect 497458 224244 497464 224256
rect 483808 224216 497464 224244
rect 483808 224204 483814 224216
rect 497458 224204 497464 224216
rect 497516 224204 497522 224256
rect 523494 224244 523500 224256
rect 505066 224216 523500 224244
rect 102042 224068 102048 224120
rect 102100 224108 102106 224120
rect 178494 224108 178500 224120
rect 102100 224080 178500 224108
rect 102100 224068 102106 224080
rect 178494 224068 178500 224080
rect 178552 224068 178558 224120
rect 179322 224068 179328 224120
rect 179380 224108 179386 224120
rect 185578 224108 185584 224120
rect 179380 224080 185584 224108
rect 179380 224068 179386 224080
rect 185578 224068 185584 224080
rect 185636 224068 185642 224120
rect 194778 224068 194784 224120
rect 194836 224108 194842 224120
rect 250622 224108 250628 224120
rect 194836 224080 250628 224108
rect 194836 224068 194842 224080
rect 250622 224068 250628 224080
rect 250680 224068 250686 224120
rect 266262 224068 266268 224120
rect 266320 224108 266326 224120
rect 303430 224108 303436 224120
rect 266320 224080 303436 224108
rect 266320 224068 266326 224080
rect 303430 224068 303436 224080
rect 303488 224068 303494 224120
rect 304258 224068 304264 224120
rect 304316 224108 304322 224120
rect 315298 224108 315304 224120
rect 304316 224080 315304 224108
rect 304316 224068 304322 224080
rect 315298 224068 315304 224080
rect 315356 224068 315362 224120
rect 504358 224068 504364 224120
rect 504416 224108 504422 224120
rect 505066 224108 505094 224216
rect 523494 224204 523500 224216
rect 523552 224204 523558 224256
rect 535270 224204 535276 224256
rect 535328 224244 535334 224256
rect 535328 224216 543734 224244
rect 535328 224204 535334 224216
rect 543706 224176 543734 224216
rect 562318 224204 562324 224256
rect 562376 224244 562382 224256
rect 571426 224244 571432 224256
rect 562376 224216 571432 224244
rect 562376 224204 562382 224216
rect 571426 224204 571432 224216
rect 571484 224204 571490 224256
rect 651282 224204 651288 224256
rect 651340 224244 651346 224256
rect 666462 224244 666468 224256
rect 651340 224216 666468 224244
rect 651340 224204 651346 224216
rect 666462 224204 666468 224216
rect 666520 224204 666526 224256
rect 667842 224204 667848 224256
rect 667900 224244 667906 224256
rect 667900 224216 671508 224244
rect 667900 224204 667906 224216
rect 562134 224176 562140 224188
rect 543706 224148 562140 224176
rect 562134 224136 562140 224148
rect 562192 224136 562198 224188
rect 504416 224080 505094 224108
rect 504416 224068 504422 224080
rect 539962 224000 539968 224052
rect 540020 224040 540026 224052
rect 622578 224040 622584 224052
rect 540020 224012 622584 224040
rect 540020 224000 540026 224012
rect 622578 224000 622584 224012
rect 622636 224000 622642 224052
rect 669038 224000 669044 224052
rect 669096 224040 669102 224052
rect 669096 224012 671398 224040
rect 669096 224000 669102 224012
rect 105998 223932 106004 223984
rect 106056 223972 106062 223984
rect 181070 223972 181076 223984
rect 106056 223944 181076 223972
rect 106056 223932 106062 223944
rect 181070 223932 181076 223944
rect 181128 223932 181134 223984
rect 185394 223932 185400 223984
rect 185452 223972 185458 223984
rect 194594 223972 194600 223984
rect 185452 223944 194600 223972
rect 185452 223932 185458 223944
rect 194594 223932 194600 223944
rect 194652 223932 194658 223984
rect 194962 223932 194968 223984
rect 195020 223972 195026 223984
rect 199838 223972 199844 223984
rect 195020 223944 199844 223972
rect 195020 223932 195026 223944
rect 199838 223932 199844 223944
rect 199896 223932 199902 223984
rect 201402 223932 201408 223984
rect 201460 223972 201466 223984
rect 255774 223972 255780 223984
rect 201460 223944 255780 223972
rect 201460 223932 201466 223944
rect 255774 223932 255780 223944
rect 255832 223932 255838 223984
rect 279418 223864 279424 223916
rect 279476 223904 279482 223916
rect 284754 223904 284760 223916
rect 279476 223876 284760 223904
rect 279476 223864 279482 223876
rect 284754 223864 284760 223876
rect 284812 223864 284818 223916
rect 524414 223864 524420 223916
rect 524472 223904 524478 223916
rect 525058 223904 525064 223916
rect 524472 223876 525064 223904
rect 524472 223864 524478 223876
rect 525058 223864 525064 223876
rect 525116 223904 525122 223916
rect 619634 223904 619640 223916
rect 525116 223876 619640 223904
rect 525116 223864 525122 223876
rect 619634 223864 619640 223876
rect 619692 223864 619698 223916
rect 671252 223848 671304 223854
rect 108666 223796 108672 223848
rect 108724 223836 108730 223848
rect 183646 223836 183652 223848
rect 108724 223808 183652 223836
rect 108724 223796 108730 223808
rect 183646 223796 183652 223808
rect 183704 223796 183710 223848
rect 184382 223796 184388 223848
rect 184440 223836 184446 223848
rect 207474 223836 207480 223848
rect 184440 223808 207480 223836
rect 184440 223796 184446 223808
rect 207474 223796 207480 223808
rect 207532 223796 207538 223848
rect 227530 223796 227536 223848
rect 227588 223836 227594 223848
rect 273162 223836 273168 223848
rect 227588 223808 273168 223836
rect 227588 223796 227594 223808
rect 273162 223796 273168 223808
rect 273220 223796 273226 223848
rect 671252 223790 671304 223796
rect 505186 223728 505192 223780
rect 505244 223768 505250 223780
rect 507670 223768 507676 223780
rect 505244 223740 507676 223768
rect 505244 223728 505250 223740
rect 507670 223728 507676 223740
rect 507728 223728 507734 223780
rect 517698 223728 517704 223780
rect 517756 223768 517762 223780
rect 617058 223768 617064 223780
rect 517756 223740 617064 223768
rect 517756 223728 517762 223740
rect 617058 223728 617064 223740
rect 617116 223728 617122 223780
rect 115290 223660 115296 223712
rect 115348 223700 115354 223712
rect 188798 223700 188804 223712
rect 115348 223672 188804 223700
rect 115348 223660 115354 223672
rect 188798 223660 188804 223672
rect 188856 223660 188862 223712
rect 191558 223660 191564 223712
rect 191616 223700 191622 223712
rect 194962 223700 194968 223712
rect 191616 223672 194968 223700
rect 191616 223660 191622 223672
rect 194962 223660 194968 223672
rect 195020 223660 195026 223712
rect 207658 223660 207664 223712
rect 207716 223700 207722 223712
rect 228082 223700 228088 223712
rect 207716 223672 228088 223700
rect 207716 223660 207722 223672
rect 228082 223660 228088 223672
rect 228140 223660 228146 223712
rect 460566 223660 460572 223712
rect 460624 223700 460630 223712
rect 463142 223700 463148 223712
rect 460624 223672 463148 223700
rect 460624 223660 460630 223672
rect 463142 223660 463148 223672
rect 463200 223660 463206 223712
rect 505370 223592 505376 223644
rect 505428 223632 505434 223644
rect 614942 223632 614948 223644
rect 505428 223604 614948 223632
rect 505428 223592 505434 223604
rect 614942 223592 614948 223604
rect 615000 223592 615006 223644
rect 671160 223576 671212 223582
rect 87966 223524 87972 223576
rect 88024 223564 88030 223576
rect 164970 223564 164976 223576
rect 88024 223536 164976 223564
rect 88024 223524 88030 223536
rect 164970 223524 164976 223536
rect 165028 223524 165034 223576
rect 171778 223524 171784 223576
rect 171836 223564 171842 223576
rect 181714 223564 181720 223576
rect 171836 223536 181720 223564
rect 171836 223524 171842 223536
rect 181714 223524 181720 223536
rect 181772 223524 181778 223576
rect 183186 223524 183192 223576
rect 183244 223564 183250 223576
rect 184658 223564 184664 223576
rect 183244 223536 184664 223564
rect 183244 223524 183250 223536
rect 184658 223524 184664 223536
rect 184716 223524 184722 223576
rect 187326 223524 187332 223576
rect 187384 223564 187390 223576
rect 242250 223564 242256 223576
rect 187384 223536 242256 223564
rect 187384 223524 187390 223536
rect 242250 223524 242256 223536
rect 242308 223524 242314 223576
rect 249426 223524 249432 223576
rect 249484 223564 249490 223576
rect 276290 223564 276296 223576
rect 249484 223536 276296 223564
rect 249484 223524 249490 223536
rect 276290 223524 276296 223536
rect 276348 223524 276354 223576
rect 278590 223524 278596 223576
rect 278648 223564 278654 223576
rect 315022 223564 315028 223576
rect 278648 223536 315028 223564
rect 278648 223524 278654 223536
rect 315022 223524 315028 223536
rect 315080 223524 315086 223576
rect 406746 223524 406752 223576
rect 406804 223564 406810 223576
rect 414842 223564 414848 223576
rect 406804 223536 414848 223564
rect 406804 223524 406810 223536
rect 414842 223524 414848 223536
rect 414900 223524 414906 223576
rect 454862 223524 454868 223576
rect 454920 223564 454926 223576
rect 460474 223564 460480 223576
rect 454920 223536 460480 223564
rect 454920 223524 454926 223536
rect 460474 223524 460480 223536
rect 460532 223524 460538 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 671160 223518 671212 223524
rect 562134 223456 562140 223508
rect 562192 223496 562198 223508
rect 563330 223496 563336 223508
rect 562192 223468 563336 223496
rect 562192 223456 562198 223468
rect 563330 223456 563336 223468
rect 563388 223456 563394 223508
rect 671022 223440 671074 223446
rect 88886 223388 88892 223440
rect 88944 223428 88950 223440
rect 107654 223428 107660 223440
rect 88944 223400 107660 223428
rect 88944 223388 88950 223400
rect 107654 223388 107660 223400
rect 107712 223388 107718 223440
rect 108298 223388 108304 223440
rect 108356 223428 108362 223440
rect 175918 223428 175924 223440
rect 108356 223400 175924 223428
rect 108356 223388 108362 223400
rect 175918 223388 175924 223400
rect 175976 223388 175982 223440
rect 184842 223388 184848 223440
rect 184900 223428 184906 223440
rect 239674 223428 239680 223440
rect 184900 223400 239680 223428
rect 184900 223388 184906 223400
rect 239674 223388 239680 223400
rect 239732 223388 239738 223440
rect 244090 223388 244096 223440
rect 244148 223428 244154 223440
rect 286042 223428 286048 223440
rect 244148 223400 286048 223428
rect 244148 223388 244154 223400
rect 286042 223388 286048 223400
rect 286100 223388 286106 223440
rect 291194 223428 291200 223440
rect 287026 223400 291200 223428
rect 81342 223252 81348 223304
rect 81400 223292 81406 223304
rect 151906 223292 151912 223304
rect 81400 223264 151912 223292
rect 81400 223252 81406 223264
rect 151906 223252 151912 223264
rect 151964 223252 151970 223304
rect 156414 223292 156420 223304
rect 152108 223264 156420 223292
rect 68738 223116 68744 223168
rect 68796 223156 68802 223168
rect 146478 223156 146484 223168
rect 68796 223128 146484 223156
rect 68796 223116 68802 223128
rect 146478 223116 146484 223128
rect 146536 223116 146542 223168
rect 146662 223116 146668 223168
rect 146720 223156 146726 223168
rect 152108 223156 152136 223264
rect 156414 223252 156420 223264
rect 156472 223252 156478 223304
rect 156598 223252 156604 223304
rect 156656 223292 156662 223304
rect 161934 223292 161940 223304
rect 156656 223264 161940 223292
rect 156656 223252 156662 223264
rect 161934 223252 161940 223264
rect 161992 223252 161998 223304
rect 162302 223252 162308 223304
rect 162360 223292 162366 223304
rect 186866 223292 186872 223304
rect 162360 223264 186872 223292
rect 162360 223252 162366 223264
rect 186866 223252 186872 223264
rect 186924 223252 186930 223304
rect 188154 223252 188160 223304
rect 188212 223292 188218 223304
rect 245102 223292 245108 223304
rect 188212 223264 245108 223292
rect 188212 223252 188218 223264
rect 245102 223252 245108 223264
rect 245160 223252 245166 223304
rect 250898 223252 250904 223304
rect 250956 223292 250962 223304
rect 287026 223292 287054 223400
rect 291194 223388 291200 223400
rect 291252 223388 291258 223440
rect 316678 223388 316684 223440
rect 316736 223428 316742 223440
rect 327258 223428 327264 223440
rect 316736 223400 327264 223428
rect 316736 223388 316742 223400
rect 327258 223388 327264 223400
rect 327316 223388 327322 223440
rect 517514 223388 517520 223440
rect 517572 223428 517578 223440
rect 532510 223428 532516 223440
rect 517572 223400 532516 223428
rect 517572 223388 517578 223400
rect 532510 223388 532516 223400
rect 532568 223388 532574 223440
rect 534810 223388 534816 223440
rect 534868 223428 534874 223440
rect 547414 223428 547420 223440
rect 534868 223400 547420 223428
rect 534868 223388 534874 223400
rect 547414 223388 547420 223400
rect 547472 223388 547478 223440
rect 671022 223382 671074 223388
rect 297542 223320 297548 223372
rect 297600 223360 297606 223372
rect 305362 223360 305368 223372
rect 297600 223332 305368 223360
rect 297600 223320 297606 223332
rect 305362 223320 305368 223332
rect 305420 223320 305426 223372
rect 250956 223264 287054 223292
rect 250956 223252 250962 223264
rect 288986 223252 288992 223304
rect 289044 223292 289050 223304
rect 295058 223292 295064 223304
rect 289044 223264 295064 223292
rect 289044 223252 289050 223264
rect 295058 223252 295064 223264
rect 295116 223252 295122 223304
rect 307662 223252 307668 223304
rect 307720 223292 307726 223304
rect 335630 223292 335636 223304
rect 307720 223264 335636 223292
rect 307720 223252 307726 223264
rect 335630 223252 335636 223264
rect 335688 223252 335694 223304
rect 337930 223252 337936 223304
rect 337988 223292 337994 223304
rect 359182 223292 359188 223304
rect 337988 223264 359188 223292
rect 337988 223252 337994 223264
rect 359182 223252 359188 223264
rect 359240 223252 359246 223304
rect 493042 223252 493048 223304
rect 493100 223292 493106 223304
rect 508498 223292 508504 223304
rect 493100 223264 508504 223292
rect 493100 223252 493106 223264
rect 508498 223252 508504 223264
rect 508556 223252 508562 223304
rect 514662 223252 514668 223304
rect 514720 223292 514726 223304
rect 535454 223292 535460 223304
rect 514720 223264 535460 223292
rect 514720 223252 514726 223264
rect 535454 223252 535460 223264
rect 535512 223252 535518 223304
rect 154942 223156 154948 223168
rect 146720 223128 152136 223156
rect 152200 223128 154948 223156
rect 146720 223116 146726 223128
rect 75822 222980 75828 223032
rect 75880 223020 75886 223032
rect 152200 223020 152228 223128
rect 154942 223116 154948 223128
rect 155000 223116 155006 223168
rect 156414 223116 156420 223168
rect 156472 223156 156478 223168
rect 176102 223156 176108 223168
rect 156472 223128 176108 223156
rect 156472 223116 156478 223128
rect 176102 223116 176108 223128
rect 176160 223116 176166 223168
rect 181990 223116 181996 223168
rect 182048 223156 182054 223168
rect 240318 223156 240324 223168
rect 182048 223128 240324 223156
rect 182048 223116 182054 223128
rect 240318 223116 240324 223128
rect 240376 223116 240382 223168
rect 241330 223116 241336 223168
rect 241388 223156 241394 223168
rect 283466 223156 283472 223168
rect 241388 223128 283472 223156
rect 241388 223116 241394 223128
rect 283466 223116 283472 223128
rect 283524 223116 283530 223168
rect 288250 223116 288256 223168
rect 288308 223156 288314 223168
rect 321462 223156 321468 223168
rect 288308 223128 321468 223156
rect 288308 223116 288314 223128
rect 321462 223116 321468 223128
rect 321520 223116 321526 223168
rect 323946 223116 323952 223168
rect 324004 223156 324010 223168
rect 348510 223156 348516 223168
rect 324004 223128 348516 223156
rect 324004 223116 324010 223128
rect 348510 223116 348516 223128
rect 348568 223116 348574 223168
rect 358538 223116 358544 223168
rect 358596 223156 358602 223168
rect 374638 223156 374644 223168
rect 358596 223128 374644 223156
rect 358596 223116 358602 223128
rect 374638 223116 374644 223128
rect 374696 223116 374702 223168
rect 483106 223116 483112 223168
rect 483164 223156 483170 223168
rect 496078 223156 496084 223168
rect 483164 223128 496084 223156
rect 483164 223116 483170 223128
rect 496078 223116 496084 223128
rect 496136 223116 496142 223168
rect 503346 223116 503352 223168
rect 503404 223156 503410 223168
rect 521746 223156 521752 223168
rect 503404 223128 521752 223156
rect 503404 223116 503410 223128
rect 521746 223116 521752 223128
rect 521804 223116 521810 223168
rect 529474 223116 529480 223168
rect 529532 223156 529538 223168
rect 555694 223156 555700 223168
rect 529532 223128 555700 223156
rect 529532 223116 529538 223128
rect 555694 223116 555700 223128
rect 555752 223116 555758 223168
rect 669038 223116 669044 223168
rect 669096 223156 669102 223168
rect 669096 223128 670956 223156
rect 669096 223116 669102 223128
rect 75880 222992 152228 223020
rect 75880 222980 75886 222992
rect 152366 222980 152372 223032
rect 152424 223020 152430 223032
rect 152424 222992 157012 223020
rect 152424 222980 152430 222992
rect 71406 222844 71412 222896
rect 71464 222884 71470 222896
rect 151630 222884 151636 222896
rect 71464 222856 151636 222884
rect 71464 222844 71470 222856
rect 151630 222844 151636 222856
rect 151688 222844 151694 222896
rect 151768 222844 151774 222896
rect 151826 222884 151832 222896
rect 156414 222884 156420 222896
rect 151826 222856 156420 222884
rect 151826 222844 151832 222856
rect 156414 222844 156420 222856
rect 156472 222844 156478 222896
rect 156984 222884 157012 222992
rect 157518 222980 157524 223032
rect 157576 223020 157582 223032
rect 219066 223020 219072 223032
rect 157576 222992 219072 223020
rect 157576 222980 157582 222992
rect 219066 222980 219072 222992
rect 219124 222980 219130 223032
rect 245286 222980 245292 223032
rect 245344 223020 245350 223032
rect 289262 223020 289268 223032
rect 245344 222992 289268 223020
rect 245344 222980 245350 222992
rect 289262 222980 289268 222992
rect 289320 222980 289326 223032
rect 291654 222980 291660 223032
rect 291712 223020 291718 223032
rect 300210 223020 300216 223032
rect 291712 222992 300216 223020
rect 291712 222980 291718 222992
rect 300210 222980 300216 222992
rect 300268 222980 300274 223032
rect 315666 222980 315672 223032
rect 315724 223020 315730 223032
rect 344646 223020 344652 223032
rect 315724 222992 344652 223020
rect 315724 222980 315730 222992
rect 344646 222980 344652 222992
rect 344704 222980 344710 223032
rect 346578 223020 346584 223032
rect 344986 222992 346584 223020
rect 171778 222884 171784 222896
rect 156984 222856 171784 222884
rect 171778 222844 171784 222856
rect 171836 222844 171842 222896
rect 172882 222844 172888 222896
rect 172940 222884 172946 222896
rect 212626 222884 212632 222896
rect 172940 222856 212632 222884
rect 172940 222844 172946 222856
rect 212626 222844 212632 222856
rect 212684 222844 212690 222896
rect 213178 222844 213184 222896
rect 213236 222884 213242 222896
rect 233326 222884 233332 222896
rect 213236 222856 233332 222884
rect 213236 222844 213242 222856
rect 233326 222844 233332 222856
rect 233384 222844 233390 222896
rect 234522 222844 234528 222896
rect 234580 222884 234586 222896
rect 281534 222884 281540 222896
rect 234580 222856 281540 222884
rect 234580 222844 234586 222856
rect 281534 222844 281540 222856
rect 281592 222844 281598 222896
rect 282730 222844 282736 222896
rect 282788 222884 282794 222896
rect 316310 222884 316316 222896
rect 282788 222856 316316 222884
rect 282788 222844 282794 222856
rect 316310 222844 316316 222856
rect 316368 222844 316374 222896
rect 321462 222844 321468 222896
rect 321520 222884 321526 222896
rect 344986 222884 345014 222992
rect 346578 222980 346584 222992
rect 346636 222980 346642 223032
rect 349062 222980 349068 223032
rect 349120 223020 349126 223032
rect 367186 223020 367192 223032
rect 349120 222992 367192 223020
rect 349120 222980 349126 222992
rect 367186 222980 367192 222992
rect 367244 222980 367250 223032
rect 368382 222980 368388 223032
rect 368440 223020 368446 223032
rect 382642 223020 382648 223032
rect 368440 222992 382648 223020
rect 368440 222980 368446 222992
rect 382642 222980 382648 222992
rect 382700 222980 382706 223032
rect 383562 222980 383568 223032
rect 383620 223020 383626 223032
rect 394878 223020 394884 223032
rect 383620 222992 394884 223020
rect 383620 222980 383626 222992
rect 394878 222980 394884 222992
rect 394936 222980 394942 223032
rect 486602 222980 486608 223032
rect 486660 223020 486666 223032
rect 500402 223020 500408 223032
rect 486660 222992 500408 223020
rect 486660 222980 486666 222992
rect 500402 222980 500408 222992
rect 500460 222980 500466 223032
rect 508222 222980 508228 223032
rect 508280 223020 508286 223032
rect 527174 223020 527180 223032
rect 508280 222992 527180 223020
rect 508280 222980 508286 222992
rect 527174 222980 527180 222992
rect 527232 222980 527238 223032
rect 532050 222980 532056 223032
rect 532108 223020 532114 223032
rect 559006 223020 559012 223032
rect 532108 222992 559012 223020
rect 532108 222980 532114 222992
rect 559006 222980 559012 222992
rect 559064 222980 559070 223032
rect 321520 222856 345014 222884
rect 321520 222844 321526 222856
rect 345290 222844 345296 222896
rect 345348 222884 345354 222896
rect 347866 222884 347872 222896
rect 345348 222856 347872 222884
rect 345348 222844 345354 222856
rect 347866 222844 347872 222856
rect 347924 222844 347930 222896
rect 367830 222884 367836 222896
rect 354646 222856 367836 222884
rect 85298 222708 85304 222760
rect 85356 222748 85362 222760
rect 156598 222748 156604 222760
rect 85356 222720 156604 222748
rect 85356 222708 85362 222720
rect 156598 222708 156604 222720
rect 156656 222708 156662 222760
rect 156782 222708 156788 222760
rect 156840 222748 156846 222760
rect 159818 222748 159824 222760
rect 156840 222720 159824 222748
rect 156840 222708 156846 222720
rect 159818 222708 159824 222720
rect 159876 222708 159882 222760
rect 165614 222708 165620 222760
rect 165672 222748 165678 222760
rect 192018 222748 192024 222760
rect 165672 222720 192024 222748
rect 165672 222708 165678 222720
rect 192018 222708 192024 222720
rect 192076 222708 192082 222760
rect 193950 222708 193956 222760
rect 194008 222748 194014 222760
rect 247402 222748 247408 222760
rect 194008 222720 247408 222748
rect 194008 222708 194014 222720
rect 247402 222708 247408 222720
rect 247460 222708 247466 222760
rect 284202 222708 284208 222760
rect 284260 222748 284266 222760
rect 316954 222748 316960 222760
rect 284260 222720 316960 222748
rect 284260 222708 284266 222720
rect 316954 222708 316960 222720
rect 317012 222708 317018 222760
rect 347222 222708 347228 222760
rect 347280 222748 347286 222760
rect 354646 222748 354674 222856
rect 367830 222844 367836 222856
rect 367888 222844 367894 222896
rect 375190 222844 375196 222896
rect 375248 222884 375254 222896
rect 391014 222884 391020 222896
rect 375248 222856 391020 222884
rect 375248 222844 375254 222856
rect 391014 222844 391020 222856
rect 391072 222844 391078 222896
rect 395798 222844 395804 222896
rect 395856 222884 395862 222896
rect 406470 222884 406476 222896
rect 395856 222856 406476 222884
rect 395856 222844 395862 222856
rect 406470 222844 406476 222856
rect 406528 222844 406534 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 479886 222844 479892 222896
rect 479944 222884 479950 222896
rect 492030 222884 492036 222896
rect 479944 222856 492036 222884
rect 479944 222844 479950 222856
rect 492030 222844 492036 222856
rect 492088 222844 492094 222896
rect 500770 222844 500776 222896
rect 500828 222884 500834 222896
rect 517514 222884 517520 222896
rect 500828 222856 517520 222884
rect 500828 222844 500834 222856
rect 517514 222844 517520 222856
rect 517572 222844 517578 222896
rect 519814 222844 519820 222896
rect 519872 222884 519878 222896
rect 543274 222884 543280 222896
rect 519872 222856 543280 222884
rect 519872 222844 519878 222856
rect 543274 222844 543280 222856
rect 543332 222844 543338 222896
rect 554038 222844 554044 222896
rect 554096 222884 554102 222896
rect 632698 222884 632704 222896
rect 554096 222856 632704 222884
rect 554096 222844 554102 222856
rect 632698 222844 632704 222856
rect 632756 222844 632762 222896
rect 347280 222720 354674 222748
rect 347280 222708 347286 222720
rect 558178 222708 558184 222760
rect 558236 222748 558242 222760
rect 620278 222748 620284 222760
rect 558236 222720 596174 222748
rect 558236 222708 558242 222720
rect 78582 222572 78588 222624
rect 78640 222612 78646 222624
rect 88886 222612 88892 222624
rect 78640 222584 88892 222612
rect 78640 222572 78646 222584
rect 88886 222572 88892 222584
rect 88944 222572 88950 222624
rect 99282 222572 99288 222624
rect 99340 222612 99346 222624
rect 99340 222584 103514 222612
rect 99340 222572 99346 222584
rect 103486 222476 103514 222584
rect 107654 222572 107660 222624
rect 107712 222612 107718 222624
rect 126514 222612 126520 222624
rect 107712 222584 126520 222612
rect 107712 222572 107718 222584
rect 126514 222572 126520 222584
rect 126572 222572 126578 222624
rect 191374 222612 191380 222624
rect 127084 222584 191380 222612
rect 108298 222476 108304 222488
rect 103486 222448 108304 222476
rect 108298 222436 108304 222448
rect 108356 222436 108362 222488
rect 118418 222436 118424 222488
rect 118476 222476 118482 222488
rect 127084 222476 127112 222584
rect 191374 222572 191380 222584
rect 191432 222572 191438 222624
rect 197170 222572 197176 222624
rect 197228 222612 197234 222624
rect 249978 222612 249984 222624
rect 197228 222584 249984 222612
rect 197228 222572 197234 222584
rect 249978 222572 249984 222584
rect 250036 222572 250042 222624
rect 482738 222572 482744 222624
rect 482796 222612 482802 222624
rect 593966 222612 593972 222624
rect 482796 222584 593972 222612
rect 482796 222572 482802 222584
rect 593966 222572 593972 222584
rect 594024 222572 594030 222624
rect 596146 222612 596174 222720
rect 605806 222720 620284 222748
rect 605806 222612 605834 222720
rect 620278 222708 620284 222720
rect 620336 222708 620342 222760
rect 627086 222612 627092 222624
rect 596146 222584 605834 222612
rect 619192 222584 627092 222612
rect 146662 222476 146668 222488
rect 118476 222448 127112 222476
rect 132466 222448 146668 222476
rect 118476 222436 118482 222448
rect 126514 222300 126520 222352
rect 126572 222340 126578 222352
rect 132466 222340 132494 222448
rect 146662 222436 146668 222448
rect 146720 222436 146726 222488
rect 206830 222476 206836 222488
rect 146956 222448 206836 222476
rect 126572 222312 132494 222340
rect 126572 222300 126578 222312
rect 139118 222300 139124 222352
rect 139176 222340 139182 222352
rect 146956 222340 146984 222448
rect 206830 222436 206836 222448
rect 206888 222436 206894 222488
rect 207842 222436 207848 222488
rect 207900 222476 207906 222488
rect 258350 222476 258356 222488
rect 207900 222448 258356 222476
rect 207900 222436 207906 222448
rect 258350 222436 258356 222448
rect 258408 222436 258414 222488
rect 502426 222436 502432 222488
rect 502484 222476 502490 222488
rect 558178 222476 558184 222488
rect 502484 222448 558184 222476
rect 502484 222436 502490 222448
rect 558178 222436 558184 222448
rect 558236 222436 558242 222488
rect 558546 222436 558552 222488
rect 558604 222476 558610 222488
rect 559834 222476 559840 222488
rect 558604 222448 559840 222476
rect 558604 222436 558610 222448
rect 559834 222436 559840 222448
rect 559892 222476 559898 222488
rect 619192 222476 619220 222584
rect 627086 222572 627092 222584
rect 627144 222572 627150 222624
rect 559892 222448 619220 222476
rect 559892 222436 559898 222448
rect 620278 222436 620284 222488
rect 620336 222476 620342 222488
rect 630674 222476 630680 222488
rect 620336 222448 630680 222476
rect 620336 222436 620342 222448
rect 630674 222436 630680 222448
rect 630732 222436 630738 222488
rect 490006 222368 490012 222420
rect 490064 222408 490070 222420
rect 490064 222380 499574 222408
rect 490064 222368 490070 222380
rect 139176 222312 146984 222340
rect 139176 222300 139182 222312
rect 147122 222300 147128 222352
rect 147180 222340 147186 222352
rect 211982 222340 211988 222352
rect 147180 222312 211988 222340
rect 147180 222300 147186 222312
rect 211982 222300 211988 222312
rect 212040 222300 212046 222352
rect 237006 222300 237012 222352
rect 237064 222340 237070 222352
rect 280890 222340 280896 222352
rect 237064 222312 280896 222340
rect 237064 222300 237070 222312
rect 280890 222300 280896 222312
rect 280948 222300 280954 222352
rect 484578 222300 484584 222352
rect 484636 222340 484642 222352
rect 499546 222340 499574 222380
rect 629846 222340 629852 222352
rect 484636 222312 489914 222340
rect 499546 222312 629852 222340
rect 484636 222300 484642 222312
rect 489886 222204 489914 222312
rect 629846 222300 629852 222312
rect 629904 222300 629910 222352
rect 502426 222204 502432 222216
rect 489886 222176 502432 222204
rect 502426 222164 502432 222176
rect 502484 222164 502490 222216
rect 532510 222164 532516 222216
rect 532568 222204 532574 222216
rect 621198 222204 621204 222216
rect 532568 222176 621204 222204
rect 532568 222164 532574 222176
rect 621198 222164 621204 222176
rect 621256 222164 621262 222216
rect 111978 222096 111984 222148
rect 112036 222136 112042 222148
rect 185854 222136 185860 222148
rect 112036 222108 185860 222136
rect 112036 222096 112042 222108
rect 185854 222096 185860 222108
rect 185912 222096 185918 222148
rect 200390 222096 200396 222148
rect 200448 222136 200454 222148
rect 252922 222136 252928 222148
rect 200448 222108 252928 222136
rect 200448 222096 200454 222108
rect 252922 222096 252928 222108
rect 252980 222096 252986 222148
rect 258074 222096 258080 222148
rect 258132 222136 258138 222148
rect 263870 222136 263876 222148
rect 258132 222108 263876 222136
rect 258132 222096 258138 222108
rect 263870 222096 263876 222108
rect 263928 222096 263934 222148
rect 270034 222096 270040 222148
rect 270092 222136 270098 222148
rect 306374 222136 306380 222148
rect 270092 222108 306380 222136
rect 270092 222096 270098 222108
rect 306374 222096 306380 222108
rect 306432 222096 306438 222148
rect 310698 222096 310704 222148
rect 310756 222136 310762 222148
rect 312630 222136 312636 222148
rect 310756 222108 312636 222136
rect 310756 222096 310762 222108
rect 312630 222096 312636 222108
rect 312688 222096 312694 222148
rect 331398 222096 331404 222148
rect 331456 222136 331462 222148
rect 353938 222136 353944 222148
rect 331456 222108 353944 222136
rect 331456 222096 331462 222108
rect 353938 222096 353944 222108
rect 353996 222096 354002 222148
rect 452562 222096 452568 222148
rect 452620 222136 452626 222148
rect 455598 222136 455604 222148
rect 452620 222108 455604 222136
rect 452620 222096 452626 222108
rect 455598 222096 455604 222108
rect 455656 222096 455662 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 527174 222028 527180 222080
rect 527232 222068 527238 222080
rect 528186 222068 528192 222080
rect 527232 222040 528192 222068
rect 527232 222028 527238 222040
rect 528186 222028 528192 222040
rect 528244 222068 528250 222080
rect 528244 222040 550634 222068
rect 528244 222028 528250 222040
rect 91278 221960 91284 222012
rect 91336 222000 91342 222012
rect 167178 222000 167184 222012
rect 91336 221972 167184 222000
rect 91336 221960 91342 221972
rect 167178 221960 167184 221972
rect 167236 221960 167242 222012
rect 167454 221960 167460 222012
rect 167512 222000 167518 222012
rect 172698 222000 172704 222012
rect 167512 221972 172704 222000
rect 167512 221960 167518 221972
rect 172698 221960 172704 221972
rect 172756 221960 172762 222012
rect 226518 222000 226524 222012
rect 172900 221972 226524 222000
rect 94590 221824 94596 221876
rect 94648 221864 94654 221876
rect 169846 221864 169852 221876
rect 94648 221836 169852 221864
rect 94648 221824 94654 221836
rect 169846 221824 169852 221836
rect 169904 221824 169910 221876
rect 97718 221688 97724 221740
rect 97776 221728 97782 221740
rect 167454 221728 167460 221740
rect 97776 221700 167460 221728
rect 97776 221688 97782 221700
rect 167454 221688 167460 221700
rect 167512 221688 167518 221740
rect 167638 221688 167644 221740
rect 167696 221728 167702 221740
rect 167696 221700 168052 221728
rect 167696 221688 167702 221700
rect 73890 221552 73896 221604
rect 73948 221592 73954 221604
rect 82078 221592 82084 221604
rect 73948 221564 82084 221592
rect 73948 221552 73954 221564
rect 82078 221552 82084 221564
rect 82136 221552 82142 221604
rect 86310 221552 86316 221604
rect 86368 221592 86374 221604
rect 161934 221592 161940 221604
rect 86368 221564 161940 221592
rect 86368 221552 86374 221564
rect 161934 221552 161940 221564
rect 161992 221552 161998 221604
rect 162118 221552 162124 221604
rect 162176 221592 162182 221604
rect 167822 221592 167828 221604
rect 162176 221564 167828 221592
rect 162176 221552 162182 221564
rect 167822 221552 167828 221564
rect 167880 221552 167886 221604
rect 168024 221592 168052 221700
rect 168190 221688 168196 221740
rect 168248 221728 168254 221740
rect 172900 221728 172928 221972
rect 226518 221960 226524 221972
rect 226576 221960 226582 222012
rect 232130 221960 232136 222012
rect 232188 222000 232194 222012
rect 234706 222000 234712 222012
rect 232188 221972 234712 222000
rect 232188 221960 232194 221972
rect 234706 221960 234712 221972
rect 234764 221960 234770 222012
rect 261018 221960 261024 222012
rect 261076 222000 261082 222012
rect 301682 222000 301688 222012
rect 261076 221972 301688 222000
rect 261076 221960 261082 221972
rect 301682 221960 301688 221972
rect 301740 221960 301746 222012
rect 313182 221960 313188 222012
rect 313240 222000 313246 222012
rect 340414 222000 340420 222012
rect 313240 221972 340420 222000
rect 313240 221960 313246 221972
rect 340414 221960 340420 221972
rect 340472 221960 340478 222012
rect 550606 222000 550634 222040
rect 553946 222028 553952 222080
rect 554004 222068 554010 222080
rect 596910 222068 596916 222080
rect 554004 222040 596916 222068
rect 554004 222028 554010 222040
rect 596910 222028 596916 222040
rect 596968 222028 596974 222080
rect 552934 222000 552940 222012
rect 550606 221972 552940 222000
rect 552934 221960 552940 221972
rect 552992 221960 552998 222012
rect 553228 221972 553532 222000
rect 424962 221892 424968 221944
rect 425020 221932 425026 221944
rect 429194 221932 429200 221944
rect 425020 221904 429200 221932
rect 425020 221892 425026 221904
rect 429194 221892 429200 221904
rect 429252 221892 429258 221944
rect 544010 221932 544016 221944
rect 543706 221904 544016 221932
rect 174078 221824 174084 221876
rect 174136 221864 174142 221876
rect 231946 221864 231952 221876
rect 174136 221836 231952 221864
rect 174136 221824 174142 221836
rect 231946 221824 231952 221836
rect 232004 221824 232010 221876
rect 233694 221824 233700 221876
rect 233752 221864 233758 221876
rect 277946 221864 277952 221876
rect 233752 221836 277952 221864
rect 233752 221824 233758 221836
rect 277946 221824 277952 221836
rect 278004 221824 278010 221876
rect 280062 221824 280068 221876
rect 280120 221864 280126 221876
rect 313734 221864 313740 221876
rect 280120 221836 313740 221864
rect 280120 221824 280126 221836
rect 313734 221824 313740 221836
rect 313792 221824 313798 221876
rect 318242 221824 318248 221876
rect 318300 221864 318306 221876
rect 343818 221864 343824 221876
rect 318300 221836 343824 221864
rect 318300 221824 318306 221836
rect 343818 221824 343824 221836
rect 343876 221824 343882 221876
rect 353294 221824 353300 221876
rect 353352 221864 353358 221876
rect 372706 221864 372712 221876
rect 353352 221836 372712 221864
rect 353352 221824 353358 221836
rect 372706 221824 372712 221836
rect 372764 221824 372770 221876
rect 380342 221864 380348 221876
rect 373966 221836 380348 221864
rect 168248 221700 172928 221728
rect 168248 221688 168254 221700
rect 174906 221688 174912 221740
rect 174964 221728 174970 221740
rect 174964 221700 185348 221728
rect 174964 221688 174970 221700
rect 185320 221660 185348 221700
rect 185762 221688 185768 221740
rect 185820 221728 185826 221740
rect 243078 221728 243084 221740
rect 185820 221700 243084 221728
rect 185820 221688 185826 221700
rect 243078 221688 243084 221700
rect 243136 221688 243142 221740
rect 263134 221728 263140 221740
rect 243556 221700 263140 221728
rect 185320 221632 185440 221660
rect 182634 221592 182640 221604
rect 168024 221564 182640 221592
rect 182634 221552 182640 221564
rect 182692 221552 182698 221604
rect 185412 221592 185440 221632
rect 232130 221592 232136 221604
rect 185412 221564 232136 221592
rect 232130 221552 232136 221564
rect 232188 221552 232194 221604
rect 243556 221592 243584 221700
rect 263134 221688 263140 221700
rect 263192 221688 263198 221740
rect 263502 221688 263508 221740
rect 263560 221728 263566 221740
rect 301038 221728 301044 221740
rect 263560 221700 301044 221728
rect 263560 221688 263566 221700
rect 301038 221688 301044 221700
rect 301096 221688 301102 221740
rect 303246 221688 303252 221740
rect 303304 221728 303310 221740
rect 332594 221728 332600 221740
rect 303304 221700 332600 221728
rect 303304 221688 303310 221700
rect 332594 221688 332600 221700
rect 332652 221688 332658 221740
rect 344646 221688 344652 221740
rect 344704 221728 344710 221740
rect 364518 221728 364524 221740
rect 344704 221700 364524 221728
rect 344704 221688 344710 221700
rect 364518 221688 364524 221700
rect 364576 221688 364582 221740
rect 370958 221688 370964 221740
rect 371016 221728 371022 221740
rect 373966 221728 373994 221836
rect 380342 221824 380348 221836
rect 380400 221824 380406 221876
rect 492490 221824 492496 221876
rect 492548 221864 492554 221876
rect 506842 221864 506848 221876
rect 492548 221836 506848 221864
rect 492548 221824 492554 221836
rect 506842 221824 506848 221836
rect 506900 221824 506906 221876
rect 522666 221824 522672 221876
rect 522724 221864 522730 221876
rect 543706 221864 543734 221904
rect 544010 221892 544016 221904
rect 544068 221892 544074 221944
rect 522724 221836 543734 221864
rect 522724 221824 522730 221836
rect 544194 221824 544200 221876
rect 544252 221864 544258 221876
rect 553228 221864 553256 221972
rect 553504 221932 553532 221972
rect 597094 221960 597100 222012
rect 597152 222000 597158 222012
rect 605006 222000 605012 222012
rect 597152 221972 605012 222000
rect 597152 221960 597158 221972
rect 605006 221960 605012 221972
rect 605064 221960 605070 222012
rect 553504 221904 563008 221932
rect 544252 221836 553256 221864
rect 562980 221864 563008 221904
rect 597278 221864 597284 221876
rect 562980 221836 597284 221864
rect 544252 221824 544258 221836
rect 597278 221824 597284 221836
rect 597336 221824 597342 221876
rect 597462 221824 597468 221876
rect 597520 221864 597526 221876
rect 603166 221864 603172 221876
rect 597520 221836 603172 221864
rect 597520 221824 597526 221836
rect 603166 221824 603172 221836
rect 603224 221824 603230 221876
rect 520182 221796 520188 221808
rect 514726 221768 520188 221796
rect 371016 221700 373994 221728
rect 371016 221688 371022 221700
rect 380066 221688 380072 221740
rect 380124 221728 380130 221740
rect 386506 221728 386512 221740
rect 380124 221700 386512 221728
rect 380124 221688 380130 221700
rect 386506 221688 386512 221700
rect 386564 221688 386570 221740
rect 484762 221688 484768 221740
rect 484820 221728 484826 221740
rect 497826 221728 497832 221740
rect 484820 221700 497832 221728
rect 484820 221688 484826 221700
rect 497826 221688 497832 221700
rect 497884 221688 497890 221740
rect 501322 221688 501328 221740
rect 501380 221728 501386 221740
rect 514726 221728 514754 221768
rect 520182 221756 520188 221768
rect 520240 221756 520246 221808
rect 560754 221796 560760 221808
rect 558242 221768 560760 221796
rect 501380 221700 514754 221728
rect 501380 221688 501386 221700
rect 524230 221688 524236 221740
rect 524288 221728 524294 221740
rect 543688 221728 543694 221740
rect 524288 221700 543694 221728
rect 524288 221688 524294 221700
rect 543688 221688 543694 221700
rect 543746 221688 543752 221740
rect 543826 221688 543832 221740
rect 543884 221728 543890 221740
rect 558086 221728 558092 221740
rect 543884 221700 558092 221728
rect 543884 221688 543890 221700
rect 558086 221688 558092 221700
rect 558144 221688 558150 221740
rect 233896 221564 243584 221592
rect 59354 221416 59360 221468
rect 59412 221456 59418 221468
rect 141326 221456 141332 221468
rect 59412 221428 141332 221456
rect 59412 221416 59418 221428
rect 141326 221416 141332 221428
rect 141384 221416 141390 221468
rect 147582 221416 147588 221468
rect 147640 221456 147646 221468
rect 204898 221456 204904 221468
rect 147640 221428 204904 221456
rect 147640 221416 147646 221428
rect 204898 221416 204904 221428
rect 204956 221416 204962 221468
rect 205082 221416 205088 221468
rect 205140 221456 205146 221468
rect 220170 221456 220176 221468
rect 205140 221428 220176 221456
rect 205140 221416 205146 221428
rect 220170 221416 220176 221428
rect 220228 221416 220234 221468
rect 220998 221416 221004 221468
rect 221056 221456 221062 221468
rect 233896 221456 233924 221564
rect 243722 221552 243728 221604
rect 243780 221592 243786 221604
rect 283742 221592 283748 221604
rect 243780 221564 283748 221592
rect 243780 221552 243786 221564
rect 283742 221552 283748 221564
rect 283800 221552 283806 221604
rect 302418 221552 302424 221604
rect 302476 221592 302482 221604
rect 334066 221592 334072 221604
rect 302476 221564 334072 221592
rect 302476 221552 302482 221564
rect 334066 221552 334072 221564
rect 334124 221552 334130 221604
rect 348786 221552 348792 221604
rect 348844 221592 348850 221604
rect 370038 221592 370044 221604
rect 348844 221564 370044 221592
rect 348844 221552 348850 221564
rect 370038 221552 370044 221564
rect 370096 221552 370102 221604
rect 373718 221552 373724 221604
rect 373776 221592 373782 221604
rect 384298 221592 384304 221604
rect 373776 221564 384304 221592
rect 373776 221552 373782 221564
rect 384298 221552 384304 221564
rect 384356 221552 384362 221604
rect 391014 221552 391020 221604
rect 391072 221592 391078 221604
rect 400398 221592 400404 221604
rect 391072 221564 400404 221592
rect 391072 221552 391078 221564
rect 400398 221552 400404 221564
rect 400456 221552 400462 221604
rect 401318 221552 401324 221604
rect 401376 221592 401382 221604
rect 405826 221592 405832 221604
rect 401376 221564 405832 221592
rect 401376 221552 401382 221564
rect 405826 221552 405832 221564
rect 405884 221552 405890 221604
rect 475838 221552 475844 221604
rect 475896 221592 475902 221604
rect 486142 221592 486148 221604
rect 475896 221564 486148 221592
rect 475896 221552 475902 221564
rect 486142 221552 486148 221564
rect 486200 221552 486206 221604
rect 496262 221552 496268 221604
rect 496320 221592 496326 221604
rect 513374 221592 513380 221604
rect 496320 221564 513380 221592
rect 496320 221552 496326 221564
rect 513374 221552 513380 221564
rect 513432 221552 513438 221604
rect 516962 221552 516968 221604
rect 517020 221592 517026 221604
rect 527542 221592 527548 221604
rect 517020 221564 527548 221592
rect 517020 221552 517026 221564
rect 527542 221552 527548 221564
rect 527600 221552 527606 221604
rect 533982 221552 533988 221604
rect 534040 221592 534046 221604
rect 558242 221592 558270 221768
rect 560754 221756 560760 221768
rect 560812 221756 560818 221808
rect 560938 221756 560944 221808
rect 560996 221796 561002 221808
rect 562686 221796 562692 221808
rect 560996 221768 562692 221796
rect 560996 221756 561002 221768
rect 562686 221756 562692 221768
rect 562744 221756 562750 221808
rect 562870 221688 562876 221740
rect 562928 221728 562934 221740
rect 563008 221728 563014 221740
rect 562928 221700 563014 221728
rect 562928 221688 562934 221700
rect 563008 221688 563014 221700
rect 563066 221688 563072 221740
rect 563146 221688 563152 221740
rect 563204 221728 563210 221740
rect 609422 221728 609428 221740
rect 563204 221700 609428 221728
rect 563204 221688 563210 221700
rect 609422 221688 609428 221700
rect 609480 221688 609486 221740
rect 534040 221564 558270 221592
rect 534040 221552 534046 221564
rect 558638 221552 558644 221604
rect 558696 221592 558702 221604
rect 605926 221592 605932 221604
rect 558696 221564 605932 221592
rect 558696 221552 558702 221564
rect 605926 221552 605932 221564
rect 605984 221552 605990 221604
rect 221056 221428 233924 221456
rect 221056 221416 221062 221428
rect 234062 221416 234068 221468
rect 234120 221456 234126 221468
rect 276106 221456 276112 221468
rect 234120 221428 276112 221456
rect 234120 221416 234126 221428
rect 276106 221416 276112 221428
rect 276164 221416 276170 221468
rect 284018 221416 284024 221468
rect 284076 221456 284082 221468
rect 320358 221456 320364 221468
rect 284076 221428 320364 221456
rect 284076 221416 284082 221428
rect 320358 221416 320364 221428
rect 320416 221416 320422 221468
rect 332594 221416 332600 221468
rect 332652 221456 332658 221468
rect 357526 221456 357532 221468
rect 332652 221428 357532 221456
rect 332652 221416 332658 221428
rect 357526 221416 357532 221428
rect 357584 221416 357590 221468
rect 369486 221416 369492 221468
rect 369544 221456 369550 221468
rect 384114 221456 384120 221468
rect 369544 221428 384120 221456
rect 369544 221416 369550 221428
rect 384114 221416 384120 221428
rect 384172 221416 384178 221468
rect 384390 221416 384396 221468
rect 384448 221456 384454 221468
rect 395154 221456 395160 221468
rect 384448 221428 395160 221456
rect 384448 221416 384454 221428
rect 395154 221416 395160 221428
rect 395212 221416 395218 221468
rect 396810 221416 396816 221468
rect 396868 221456 396874 221468
rect 407298 221456 407304 221468
rect 396868 221428 407304 221456
rect 396868 221416 396874 221428
rect 407298 221416 407304 221428
rect 407356 221416 407362 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 468938 221416 468944 221468
rect 468996 221456 469002 221468
rect 476206 221456 476212 221468
rect 468996 221428 476212 221456
rect 468996 221416 469002 221428
rect 476206 221416 476212 221428
rect 476264 221416 476270 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 538766 221456 538772 221468
rect 483808 221428 538772 221456
rect 483808 221416 483814 221428
rect 538766 221416 538772 221428
rect 538824 221416 538830 221468
rect 538950 221416 538956 221468
rect 539008 221456 539014 221468
rect 543090 221456 543096 221468
rect 539008 221428 543096 221456
rect 539008 221416 539014 221428
rect 543090 221416 543096 221428
rect 543148 221416 543154 221468
rect 544010 221416 544016 221468
rect 544068 221456 544074 221468
rect 597094 221456 597100 221468
rect 544068 221428 597100 221456
rect 544068 221416 544074 221428
rect 597094 221416 597100 221428
rect 597152 221416 597158 221468
rect 543274 221348 543280 221400
rect 543332 221388 543338 221400
rect 543826 221388 543832 221400
rect 543332 221360 543832 221388
rect 543332 221348 543338 221360
rect 543826 221348 543832 221360
rect 543884 221348 543890 221400
rect 597278 221348 597284 221400
rect 597336 221388 597342 221400
rect 606110 221388 606116 221400
rect 597336 221360 606116 221388
rect 597336 221348 597342 221360
rect 606110 221348 606116 221360
rect 606168 221348 606174 221400
rect 104526 221280 104532 221332
rect 104584 221320 104590 221332
rect 176470 221320 176476 221332
rect 104584 221292 176476 221320
rect 104584 221280 104590 221292
rect 176470 221280 176476 221292
rect 176528 221280 176534 221332
rect 176626 221292 185532 221320
rect 111150 221144 111156 221196
rect 111208 221184 111214 221196
rect 167638 221184 167644 221196
rect 111208 221156 167644 221184
rect 111208 221144 111214 221156
rect 167638 221144 167644 221156
rect 167696 221144 167702 221196
rect 167822 221144 167828 221196
rect 167880 221184 167886 221196
rect 176626 221184 176654 221292
rect 185504 221252 185532 221292
rect 185854 221280 185860 221332
rect 185912 221320 185918 221332
rect 234246 221320 234252 221332
rect 185912 221292 234252 221320
rect 185912 221280 185918 221292
rect 234246 221280 234252 221292
rect 234304 221280 234310 221332
rect 237834 221280 237840 221332
rect 237892 221320 237898 221332
rect 243722 221320 243728 221332
rect 237892 221292 243728 221320
rect 237892 221280 237898 221292
rect 243722 221280 243728 221292
rect 243780 221280 243786 221332
rect 266814 221280 266820 221332
rect 266872 221320 266878 221332
rect 303798 221320 303804 221332
rect 266872 221292 303804 221320
rect 266872 221280 266878 221292
rect 303798 221280 303804 221292
rect 303856 221280 303862 221332
rect 185504 221224 185716 221252
rect 167880 221156 176654 221184
rect 167880 221144 167886 221156
rect 177298 221144 177304 221196
rect 177356 221184 177362 221196
rect 185302 221184 185308 221196
rect 177356 221156 185308 221184
rect 177356 221144 177362 221156
rect 185302 221144 185308 221156
rect 185360 221144 185366 221196
rect 185688 221184 185716 221224
rect 523494 221212 523500 221264
rect 523552 221252 523558 221264
rect 601694 221252 601700 221264
rect 523552 221224 601700 221252
rect 523552 221212 523558 221224
rect 601694 221212 601700 221224
rect 601752 221212 601758 221264
rect 185688 221156 200114 221184
rect 124398 221008 124404 221060
rect 124456 221048 124462 221060
rect 193306 221048 193312 221060
rect 124456 221020 193312 221048
rect 124456 221008 124462 221020
rect 193306 221008 193312 221020
rect 193364 221008 193370 221060
rect 200086 221048 200114 221156
rect 204898 221144 204904 221196
rect 204956 221184 204962 221196
rect 211338 221184 211344 221196
rect 204956 221156 211344 221184
rect 204956 221144 204962 221156
rect 211338 221144 211344 221156
rect 211396 221144 211402 221196
rect 211522 221144 211528 221196
rect 211580 221184 211586 221196
rect 260834 221184 260840 221196
rect 211580 221156 260840 221184
rect 211580 221144 211586 221156
rect 260834 221144 260840 221156
rect 260892 221144 260898 221196
rect 517514 221076 517520 221128
rect 517572 221116 517578 221128
rect 518434 221116 518440 221128
rect 517572 221088 518440 221116
rect 517572 221076 517578 221088
rect 518434 221076 518440 221088
rect 518492 221116 518498 221128
rect 600590 221116 600596 221128
rect 518492 221088 600596 221116
rect 518492 221076 518498 221088
rect 600590 221076 600596 221088
rect 600648 221076 600654 221128
rect 205082 221048 205088 221060
rect 200086 221020 205088 221048
rect 205082 221008 205088 221020
rect 205140 221008 205146 221060
rect 218146 221008 218152 221060
rect 218204 221048 218210 221060
rect 220998 221048 221004 221060
rect 218204 221020 221004 221048
rect 218204 221008 218210 221020
rect 220998 221008 221004 221020
rect 221056 221008 221062 221060
rect 223482 221008 223488 221060
rect 223540 221048 223546 221060
rect 268194 221048 268200 221060
rect 223540 221020 268200 221048
rect 223540 221008 223546 221020
rect 268194 221008 268200 221020
rect 268252 221008 268258 221060
rect 82998 220940 83004 220992
rect 83056 220980 83062 220992
rect 83056 220952 93854 220980
rect 83056 220940 83062 220952
rect 93826 220912 93854 220952
rect 521010 220940 521016 220992
rect 521068 220980 521074 220992
rect 601326 220980 601332 220992
rect 521068 220952 601332 220980
rect 521068 220940 521074 220952
rect 601326 220940 601332 220952
rect 601384 220940 601390 220992
rect 151078 220912 151084 220924
rect 93826 220884 151084 220912
rect 151078 220872 151084 220884
rect 151136 220872 151142 220924
rect 155034 220872 155040 220924
rect 155092 220912 155098 220924
rect 162118 220912 162124 220924
rect 155092 220884 162124 220912
rect 155092 220872 155098 220884
rect 162118 220872 162124 220884
rect 162176 220872 162182 220924
rect 163774 220872 163780 220924
rect 163832 220912 163838 220924
rect 163832 220884 166626 220912
rect 163832 220872 163838 220884
rect 80514 220804 80520 220856
rect 80572 220844 80578 220856
rect 86126 220844 86132 220856
rect 80572 220816 86132 220844
rect 80572 220804 80578 220816
rect 86126 220804 86132 220816
rect 86184 220804 86190 220856
rect 166598 220844 166626 220884
rect 167086 220872 167092 220924
rect 167144 220912 167150 220924
rect 222286 220912 222292 220924
rect 167144 220884 222292 220912
rect 167144 220872 167150 220884
rect 222286 220872 222292 220884
rect 222344 220872 222350 220924
rect 227898 220872 227904 220924
rect 227956 220912 227962 220924
rect 234062 220912 234068 220924
rect 227956 220884 234068 220912
rect 227956 220872 227962 220884
rect 234062 220872 234068 220884
rect 234120 220872 234126 220924
rect 253842 220872 253848 220924
rect 253900 220912 253906 220924
rect 258626 220912 258632 220924
rect 253900 220884 258632 220912
rect 253900 220872 253906 220884
rect 258626 220872 258632 220884
rect 258684 220872 258690 220924
rect 166598 220816 166672 220844
rect 101214 220736 101220 220788
rect 101272 220776 101278 220788
rect 166442 220776 166448 220788
rect 101272 220748 166448 220776
rect 101272 220736 101278 220748
rect 166442 220736 166448 220748
rect 166500 220736 166506 220788
rect 166644 220776 166672 220816
rect 418338 220804 418344 220856
rect 418396 220844 418402 220856
rect 424042 220844 424048 220856
rect 418396 220816 424048 220844
rect 418396 220804 418402 220816
rect 424042 220804 424048 220816
rect 424100 220804 424106 220856
rect 456702 220804 456708 220856
rect 456760 220844 456766 220856
rect 462130 220844 462136 220856
rect 456760 220816 462136 220844
rect 456760 220804 456766 220816
rect 462130 220804 462136 220816
rect 462188 220804 462194 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 471330 220844 471336 220856
rect 466144 220816 471336 220844
rect 466144 220804 466150 220816
rect 471330 220804 471336 220816
rect 471388 220804 471394 220856
rect 515766 220804 515772 220856
rect 515824 220844 515830 220856
rect 600314 220844 600320 220856
rect 515824 220816 600320 220844
rect 515824 220804 515830 220816
rect 600314 220804 600320 220816
rect 600372 220804 600378 220856
rect 166644 220748 166764 220776
rect 76374 220600 76380 220652
rect 76432 220640 76438 220652
rect 156138 220640 156144 220652
rect 76432 220612 156144 220640
rect 76432 220600 76438 220612
rect 156138 220600 156144 220612
rect 156196 220600 156202 220652
rect 156598 220600 156604 220652
rect 156656 220640 156662 220652
rect 166442 220640 166448 220652
rect 156656 220612 166448 220640
rect 156656 220600 156662 220612
rect 166442 220600 166448 220612
rect 166500 220600 166506 220652
rect 166736 220640 166764 220748
rect 167178 220736 167184 220788
rect 167236 220776 167242 220788
rect 176470 220776 176476 220788
rect 167236 220748 176476 220776
rect 167236 220736 167242 220748
rect 176470 220736 176476 220748
rect 176528 220736 176534 220788
rect 176608 220736 176614 220788
rect 176666 220776 176672 220788
rect 180518 220776 180524 220788
rect 176666 220748 180524 220776
rect 176666 220736 176672 220748
rect 180518 220736 180524 220748
rect 180576 220736 180582 220788
rect 180702 220736 180708 220788
rect 180760 220776 180766 220788
rect 236730 220776 236736 220788
rect 180760 220748 236736 220776
rect 180760 220736 180766 220748
rect 236730 220736 236736 220748
rect 236788 220736 236794 220788
rect 254394 220736 254400 220788
rect 254452 220776 254458 220788
rect 296806 220776 296812 220788
rect 254452 220748 296812 220776
rect 254452 220736 254458 220748
rect 296806 220736 296812 220748
rect 296864 220736 296870 220788
rect 340046 220736 340052 220788
rect 340104 220776 340110 220788
rect 342346 220776 342352 220788
rect 340104 220748 342352 220776
rect 340104 220736 340110 220748
rect 342346 220736 342352 220748
rect 342404 220736 342410 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418154 220776 418160 220788
rect 414256 220748 418160 220776
rect 414256 220736 414262 220748
rect 418154 220736 418160 220748
rect 418212 220736 418218 220788
rect 431954 220736 431960 220788
rect 432012 220776 432018 220788
rect 434806 220776 434812 220788
rect 432012 220748 434812 220776
rect 432012 220736 432018 220748
rect 434806 220736 434812 220748
rect 434864 220736 434870 220788
rect 473998 220736 474004 220788
rect 474056 220776 474062 220788
rect 475378 220776 475384 220788
rect 474056 220748 475384 220776
rect 474056 220736 474062 220748
rect 475378 220736 475384 220748
rect 475436 220736 475442 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 500218 220736 500224 220788
rect 500276 220776 500282 220788
rect 511810 220776 511816 220788
rect 500276 220748 511816 220776
rect 500276 220736 500282 220748
rect 511810 220736 511816 220748
rect 511868 220736 511874 220788
rect 601510 220776 601516 220788
rect 600884 220748 601516 220776
rect 455322 220668 455328 220720
rect 455380 220708 455386 220720
rect 458818 220708 458824 220720
rect 455380 220680 458824 220708
rect 455380 220668 455386 220680
rect 458818 220668 458824 220680
rect 458876 220668 458882 220720
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469582 220708 469588 220720
rect 465776 220680 469588 220708
rect 465776 220668 465782 220680
rect 469582 220668 469588 220680
rect 469640 220668 469646 220720
rect 543826 220668 543832 220720
rect 543884 220708 543890 220720
rect 549070 220708 549076 220720
rect 543884 220680 549076 220708
rect 543884 220668 543890 220680
rect 549070 220668 549076 220680
rect 549128 220668 549134 220720
rect 550634 220668 550640 220720
rect 550692 220708 550698 220720
rect 550818 220708 550824 220720
rect 550692 220680 550824 220708
rect 550692 220668 550698 220680
rect 550818 220668 550824 220680
rect 550876 220708 550882 220720
rect 550876 220680 560294 220708
rect 550876 220668 550882 220680
rect 221274 220640 221280 220652
rect 166736 220612 221280 220640
rect 221274 220600 221280 220612
rect 221332 220600 221338 220652
rect 223758 220640 223764 220652
rect 221568 220612 223764 220640
rect 79686 220464 79692 220516
rect 79744 220504 79750 220516
rect 151722 220504 151728 220516
rect 79744 220476 151728 220504
rect 79744 220464 79750 220476
rect 151722 220464 151728 220476
rect 151780 220464 151786 220516
rect 151906 220464 151912 220516
rect 151964 220504 151970 220516
rect 153562 220504 153568 220516
rect 151964 220476 153568 220504
rect 151964 220464 151970 220476
rect 153562 220464 153568 220476
rect 153620 220464 153626 220516
rect 154206 220464 154212 220516
rect 154264 220504 154270 220516
rect 156782 220504 156788 220516
rect 154264 220476 156788 220504
rect 154264 220464 154270 220476
rect 156782 220464 156788 220476
rect 156840 220464 156846 220516
rect 156966 220464 156972 220516
rect 157024 220504 157030 220516
rect 158898 220504 158904 220516
rect 157024 220476 158904 220504
rect 157024 220464 157030 220476
rect 158898 220464 158904 220476
rect 158956 220464 158962 220516
rect 160830 220464 160836 220516
rect 160888 220504 160894 220516
rect 163774 220504 163780 220516
rect 160888 220476 163780 220504
rect 160888 220464 160894 220476
rect 163774 220464 163780 220476
rect 163832 220464 163838 220516
rect 164142 220464 164148 220516
rect 164200 220504 164206 220516
rect 166902 220504 166908 220516
rect 164200 220476 166908 220504
rect 164200 220464 164206 220476
rect 166902 220464 166908 220476
rect 166960 220464 166966 220516
rect 167086 220464 167092 220516
rect 167144 220504 167150 220516
rect 221568 220504 221596 220612
rect 223758 220600 223764 220612
rect 223816 220600 223822 220652
rect 236178 220600 236184 220652
rect 236236 220640 236242 220652
rect 246482 220640 246488 220652
rect 236236 220612 246488 220640
rect 236236 220600 236242 220612
rect 246482 220600 246488 220612
rect 246540 220600 246546 220652
rect 246942 220600 246948 220652
rect 247000 220640 247006 220652
rect 288618 220640 288624 220652
rect 247000 220612 288624 220640
rect 247000 220600 247006 220612
rect 288618 220600 288624 220612
rect 288676 220600 288682 220652
rect 304902 220600 304908 220652
rect 304960 220640 304966 220652
rect 333238 220640 333244 220652
rect 304960 220612 333244 220640
rect 304960 220600 304966 220612
rect 333238 220600 333244 220612
rect 333296 220600 333302 220652
rect 509878 220600 509884 220652
rect 509936 220640 509942 220652
rect 522574 220640 522580 220652
rect 509936 220612 522580 220640
rect 509936 220600 509942 220612
rect 522574 220600 522580 220612
rect 522632 220600 522638 220652
rect 529014 220600 529020 220652
rect 529072 220640 529078 220652
rect 560266 220640 560294 220680
rect 600884 220640 600912 220748
rect 601510 220736 601516 220748
rect 601568 220736 601574 220788
rect 607306 220640 607312 220652
rect 529072 220612 543734 220640
rect 560266 220612 600912 220640
rect 600976 220612 607312 220640
rect 529072 220600 529078 220612
rect 543706 220572 543734 220612
rect 545022 220572 545028 220584
rect 543706 220544 545028 220572
rect 545022 220532 545028 220544
rect 545080 220532 545086 220584
rect 167144 220476 221596 220504
rect 167144 220464 167150 220476
rect 223758 220464 223764 220516
rect 223816 220504 223822 220516
rect 270586 220504 270592 220516
rect 223816 220476 270592 220504
rect 223816 220464 223822 220476
rect 270586 220464 270592 220476
rect 270644 220464 270650 220516
rect 276750 220464 276756 220516
rect 276808 220504 276814 220516
rect 311342 220504 311348 220516
rect 276808 220476 311348 220504
rect 276808 220464 276814 220476
rect 311342 220464 311348 220476
rect 311400 220464 311406 220516
rect 328086 220464 328092 220516
rect 328144 220504 328150 220516
rect 351270 220504 351276 220516
rect 328144 220476 351276 220504
rect 328144 220464 328150 220476
rect 351270 220464 351276 220476
rect 351328 220464 351334 220516
rect 364518 220464 364524 220516
rect 364576 220504 364582 220516
rect 379698 220504 379704 220516
rect 364576 220476 379704 220504
rect 364576 220464 364582 220476
rect 379698 220464 379704 220476
rect 379756 220464 379762 220516
rect 469122 220464 469128 220516
rect 469180 220504 469186 220516
rect 474550 220504 474556 220516
rect 469180 220476 474556 220504
rect 469180 220464 469186 220476
rect 474550 220464 474556 220476
rect 474608 220464 474614 220516
rect 488442 220464 488448 220516
rect 488500 220504 488506 220516
rect 501874 220504 501880 220516
rect 488500 220476 501880 220504
rect 488500 220464 488506 220476
rect 501874 220464 501880 220476
rect 501932 220464 501938 220516
rect 511626 220464 511632 220516
rect 511684 220504 511690 220516
rect 531682 220504 531688 220516
rect 511684 220476 531688 220504
rect 511684 220464 511690 220476
rect 531682 220464 531688 220476
rect 531740 220464 531746 220516
rect 548334 220464 548340 220516
rect 548392 220504 548398 220516
rect 552842 220504 552848 220516
rect 548392 220476 552848 220504
rect 548392 220464 548398 220476
rect 552842 220464 552848 220476
rect 552900 220464 552906 220516
rect 560570 220464 560576 220516
rect 560628 220504 560634 220516
rect 562870 220504 562876 220516
rect 560628 220476 562876 220504
rect 560628 220464 560634 220476
rect 562870 220464 562876 220476
rect 562928 220464 562934 220516
rect 600976 220504 601004 220612
rect 607306 220600 607312 220612
rect 607364 220600 607370 220652
rect 563026 220476 601004 220504
rect 64598 220328 64604 220380
rect 64656 220368 64662 220380
rect 141970 220368 141976 220380
rect 64656 220340 141976 220368
rect 64656 220328 64662 220340
rect 141970 220328 141976 220340
rect 142028 220328 142034 220380
rect 151768 220328 151774 220380
rect 151826 220368 151832 220380
rect 202414 220368 202420 220380
rect 151826 220340 202420 220368
rect 151826 220328 151832 220340
rect 202414 220328 202420 220340
rect 202472 220328 202478 220380
rect 202782 220328 202788 220380
rect 202840 220368 202846 220380
rect 214558 220368 214564 220380
rect 202840 220340 214564 220368
rect 202840 220328 202846 220340
rect 214558 220328 214564 220340
rect 214616 220328 214622 220380
rect 262398 220368 262404 220380
rect 214760 220340 262404 220368
rect 151078 220300 151084 220312
rect 142126 220272 151084 220300
rect 73062 220192 73068 220244
rect 73120 220232 73126 220244
rect 142126 220232 142154 220272
rect 151078 220260 151084 220272
rect 151136 220260 151142 220312
rect 156598 220232 156604 220244
rect 73120 220204 142154 220232
rect 151280 220204 156604 220232
rect 73120 220192 73126 220204
rect 142338 220124 142344 220176
rect 142396 220164 142402 220176
rect 151280 220164 151308 220204
rect 156598 220192 156604 220204
rect 156656 220192 156662 220244
rect 156782 220192 156788 220244
rect 156840 220232 156846 220244
rect 212902 220232 212908 220244
rect 156840 220204 212908 220232
rect 156840 220192 156846 220204
rect 212902 220192 212908 220204
rect 212960 220192 212966 220244
rect 213822 220192 213828 220244
rect 213880 220232 213886 220244
rect 214760 220232 214788 220340
rect 262398 220328 262404 220340
rect 262456 220328 262462 220380
rect 262674 220328 262680 220380
rect 262732 220368 262738 220380
rect 264238 220368 264244 220380
rect 262732 220340 264244 220368
rect 262732 220328 262738 220340
rect 264238 220328 264244 220340
rect 264296 220328 264302 220380
rect 264606 220328 264612 220380
rect 264664 220368 264670 220380
rect 269298 220368 269304 220380
rect 264664 220340 269304 220368
rect 264664 220328 264670 220340
rect 269298 220328 269304 220340
rect 269356 220328 269362 220380
rect 273438 220328 273444 220380
rect 273496 220368 273502 220380
rect 309226 220368 309232 220380
rect 273496 220340 309232 220368
rect 273496 220328 273502 220340
rect 309226 220328 309232 220340
rect 309284 220328 309290 220380
rect 316494 220328 316500 220380
rect 316552 220368 316558 220380
rect 342898 220368 342904 220380
rect 316552 220340 342904 220368
rect 316552 220328 316558 220340
rect 342898 220328 342904 220340
rect 342956 220328 342962 220380
rect 351270 220328 351276 220380
rect 351328 220368 351334 220380
rect 369302 220368 369308 220380
rect 351328 220340 369308 220368
rect 351328 220328 351334 220340
rect 369302 220328 369308 220340
rect 369360 220328 369366 220380
rect 376938 220328 376944 220380
rect 376996 220368 377002 220380
rect 388438 220368 388444 220380
rect 376996 220340 388444 220368
rect 376996 220328 377002 220340
rect 388438 220328 388444 220340
rect 388496 220328 388502 220380
rect 473170 220328 473176 220380
rect 473228 220368 473234 220380
rect 481174 220368 481180 220380
rect 473228 220340 481180 220368
rect 473228 220328 473234 220340
rect 481174 220328 481180 220340
rect 481232 220328 481238 220380
rect 496446 220328 496452 220380
rect 496504 220368 496510 220380
rect 509326 220368 509332 220380
rect 496504 220340 509332 220368
rect 496504 220328 496510 220340
rect 509326 220328 509332 220340
rect 509384 220328 509390 220380
rect 515398 220328 515404 220380
rect 515456 220368 515462 220380
rect 530026 220368 530032 220380
rect 515456 220340 530032 220368
rect 515456 220328 515462 220340
rect 530026 220328 530032 220340
rect 530084 220328 530090 220380
rect 531130 220328 531136 220380
rect 531188 220368 531194 220380
rect 553394 220368 553400 220380
rect 531188 220340 553400 220368
rect 531188 220328 531194 220340
rect 553394 220328 553400 220340
rect 553452 220328 553458 220380
rect 553946 220328 553952 220380
rect 554004 220368 554010 220380
rect 563026 220368 563054 220476
rect 601142 220464 601148 220516
rect 601200 220504 601206 220516
rect 611446 220504 611452 220516
rect 601200 220476 611452 220504
rect 601200 220464 601206 220476
rect 611446 220464 611452 220476
rect 611504 220464 611510 220516
rect 566458 220368 566464 220380
rect 554004 220340 563054 220368
rect 563164 220340 566464 220368
rect 554004 220328 554010 220340
rect 213880 220204 214788 220232
rect 213880 220192 213886 220204
rect 217134 220192 217140 220244
rect 217192 220232 217198 220244
rect 265158 220232 265164 220244
rect 217192 220204 265164 220232
rect 217192 220192 217198 220204
rect 265158 220192 265164 220204
rect 265216 220192 265222 220244
rect 267642 220192 267648 220244
rect 267700 220232 267706 220244
rect 306834 220232 306840 220244
rect 267700 220204 306840 220232
rect 267700 220192 267706 220204
rect 306834 220192 306840 220204
rect 306892 220192 306898 220244
rect 309042 220192 309048 220244
rect 309100 220232 309106 220244
rect 339678 220232 339684 220244
rect 309100 220204 339684 220232
rect 309100 220192 309106 220204
rect 339678 220192 339684 220204
rect 339736 220192 339742 220244
rect 342990 220192 342996 220244
rect 343048 220232 343054 220244
rect 363322 220232 363328 220244
rect 343048 220204 363328 220232
rect 343048 220192 343054 220204
rect 363322 220192 363328 220204
rect 363380 220192 363386 220244
rect 363690 220192 363696 220244
rect 363748 220232 363754 220244
rect 381078 220232 381084 220244
rect 363748 220204 381084 220232
rect 363748 220192 363754 220204
rect 381078 220192 381084 220204
rect 381136 220192 381142 220244
rect 388438 220192 388444 220244
rect 388496 220232 388502 220244
rect 400950 220232 400956 220244
rect 388496 220204 400956 220232
rect 388496 220192 388502 220204
rect 400950 220192 400956 220204
rect 401008 220192 401014 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 472986 220192 472992 220244
rect 473044 220232 473050 220244
rect 482002 220232 482008 220244
rect 473044 220204 482008 220232
rect 473044 220192 473050 220204
rect 482002 220192 482008 220204
rect 482060 220192 482066 220244
rect 482922 220192 482928 220244
rect 482980 220232 482986 220244
rect 495342 220232 495348 220244
rect 482980 220204 495348 220232
rect 482980 220192 482986 220204
rect 495342 220192 495348 220204
rect 495400 220192 495406 220244
rect 497642 220192 497648 220244
rect 497700 220232 497706 220244
rect 515214 220232 515220 220244
rect 497700 220204 515220 220232
rect 497700 220192 497706 220204
rect 515214 220192 515220 220204
rect 515272 220192 515278 220244
rect 528370 220192 528376 220244
rect 528428 220232 528434 220244
rect 553578 220232 553584 220244
rect 528428 220204 553584 220232
rect 528428 220192 528434 220204
rect 553578 220192 553584 220204
rect 553636 220192 553642 220244
rect 563164 220232 563192 220340
rect 566458 220328 566464 220340
rect 566516 220328 566522 220380
rect 566642 220328 566648 220380
rect 566700 220368 566706 220380
rect 567286 220368 567292 220380
rect 566700 220340 567292 220368
rect 566700 220328 566706 220340
rect 567286 220328 567292 220340
rect 567344 220368 567350 220380
rect 568390 220368 568396 220380
rect 567344 220340 568396 220368
rect 567344 220328 567350 220340
rect 568390 220328 568396 220340
rect 568448 220328 568454 220380
rect 568574 220328 568580 220380
rect 568632 220368 568638 220380
rect 569770 220368 569776 220380
rect 568632 220340 569776 220368
rect 568632 220328 568638 220340
rect 569770 220328 569776 220340
rect 569828 220328 569834 220380
rect 569954 220328 569960 220380
rect 570012 220368 570018 220380
rect 572438 220368 572444 220380
rect 570012 220340 572444 220368
rect 570012 220328 570018 220340
rect 572438 220328 572444 220340
rect 572496 220328 572502 220380
rect 572990 220328 572996 220380
rect 573048 220368 573054 220380
rect 610066 220368 610072 220380
rect 573048 220340 610072 220368
rect 573048 220328 573054 220340
rect 610066 220328 610072 220340
rect 610124 220328 610130 220380
rect 563026 220204 563192 220232
rect 563026 220164 563054 220204
rect 563514 220192 563520 220244
rect 563572 220232 563578 220244
rect 572622 220232 572628 220244
rect 563572 220204 572628 220232
rect 563572 220192 563578 220204
rect 572622 220192 572628 220204
rect 572680 220192 572686 220244
rect 572806 220192 572812 220244
rect 572864 220232 572870 220244
rect 610250 220232 610256 220244
rect 572864 220204 610256 220232
rect 572864 220192 572870 220204
rect 610250 220192 610256 220204
rect 610308 220192 610314 220244
rect 142396 220136 151308 220164
rect 558196 220136 563054 220164
rect 142396 220124 142402 220136
rect 69750 220056 69756 220108
rect 69808 220096 69814 220108
rect 142154 220096 142160 220108
rect 69808 220068 142160 220096
rect 69808 220056 69814 220068
rect 142154 220056 142160 220068
rect 142212 220056 142218 220108
rect 151446 220056 151452 220108
rect 151504 220096 151510 220108
rect 214282 220096 214288 220108
rect 151504 220068 214288 220096
rect 151504 220056 151510 220068
rect 214282 220056 214288 220068
rect 214340 220056 214346 220108
rect 214558 220056 214564 220108
rect 214616 220096 214622 220108
rect 229278 220096 229284 220108
rect 214616 220068 229284 220096
rect 214616 220056 214622 220068
rect 229278 220056 229284 220068
rect 229336 220056 229342 220108
rect 230198 220056 230204 220108
rect 230256 220096 230262 220108
rect 275278 220096 275284 220108
rect 230256 220068 275284 220096
rect 230256 220056 230262 220068
rect 275278 220056 275284 220068
rect 275336 220056 275342 220108
rect 292482 220056 292488 220108
rect 292540 220096 292546 220108
rect 326154 220096 326160 220108
rect 292540 220068 326160 220096
rect 292540 220056 292546 220068
rect 326154 220056 326160 220068
rect 326212 220056 326218 220108
rect 328914 220056 328920 220108
rect 328972 220096 328978 220108
rect 354766 220096 354772 220108
rect 328972 220068 354772 220096
rect 328972 220056 328978 220068
rect 354766 220056 354772 220068
rect 354824 220056 354830 220108
rect 355410 220056 355416 220108
rect 355468 220096 355474 220108
rect 375558 220096 375564 220108
rect 355468 220068 375564 220096
rect 355468 220056 355474 220068
rect 375558 220056 375564 220068
rect 375616 220056 375622 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404722 220096 404728 220108
rect 396040 220068 404728 220096
rect 396040 220056 396046 220068
rect 404722 220056 404728 220068
rect 404780 220056 404786 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426710 220096 426716 220108
rect 421708 220068 426716 220096
rect 421708 220056 421714 220068
rect 426710 220056 426716 220068
rect 426768 220056 426774 220108
rect 478322 220056 478328 220108
rect 478380 220096 478386 220108
rect 489454 220096 489460 220108
rect 478380 220068 489460 220096
rect 478380 220056 478386 220068
rect 489454 220056 489460 220068
rect 489512 220056 489518 220108
rect 489638 220056 489644 220108
rect 489696 220096 489702 220108
rect 504358 220096 504364 220108
rect 489696 220068 504364 220096
rect 489696 220056 489702 220068
rect 504358 220056 504364 220068
rect 504416 220056 504422 220108
rect 513098 220056 513104 220108
rect 513156 220096 513162 220108
rect 534166 220096 534172 220108
rect 513156 220068 534172 220096
rect 513156 220056 513162 220068
rect 534166 220056 534172 220068
rect 534224 220056 534230 220108
rect 538122 220056 538128 220108
rect 538180 220096 538186 220108
rect 558196 220096 558224 220136
rect 538180 220068 558224 220096
rect 538180 220056 538186 220068
rect 586514 220056 586520 220108
rect 586572 220096 586578 220108
rect 633434 220096 633440 220108
rect 586572 220068 633440 220096
rect 586572 220056 586578 220068
rect 633434 220056 633440 220068
rect 633492 220056 633498 220108
rect 586330 220028 586336 220040
rect 558288 220000 586336 220028
rect 107838 219920 107844 219972
rect 107896 219960 107902 219972
rect 127618 219960 127624 219972
rect 107896 219932 127624 219960
rect 107896 219920 107902 219932
rect 127618 219920 127624 219932
rect 127676 219920 127682 219972
rect 127802 219920 127808 219972
rect 127860 219960 127866 219972
rect 127860 219932 185348 219960
rect 127860 219920 127866 219932
rect 185320 219892 185348 219932
rect 185762 219920 185768 219972
rect 185820 219960 185826 219972
rect 185820 219932 190316 219960
rect 185820 219920 185826 219932
rect 185320 219864 185440 219892
rect 114462 219784 114468 219836
rect 114520 219824 114526 219836
rect 185118 219824 185124 219836
rect 114520 219796 185124 219824
rect 114520 219784 114526 219796
rect 185118 219784 185124 219796
rect 185176 219784 185182 219836
rect 185412 219824 185440 219864
rect 190086 219824 190092 219836
rect 185412 219796 190092 219824
rect 190086 219784 190092 219796
rect 190144 219784 190150 219836
rect 190288 219824 190316 219932
rect 190638 219920 190644 219972
rect 190696 219960 190702 219972
rect 244458 219960 244464 219972
rect 190696 219932 244464 219960
rect 190696 219920 190702 219932
rect 244458 219920 244464 219932
rect 244516 219920 244522 219972
rect 253566 219920 253572 219972
rect 253624 219960 253630 219972
rect 293310 219960 293316 219972
rect 253624 219932 293316 219960
rect 253624 219920 253630 219932
rect 293310 219920 293316 219932
rect 293368 219920 293374 219972
rect 558288 219960 558316 220000
rect 586330 219988 586336 220000
rect 586388 219988 586394 220040
rect 550606 219932 558316 219960
rect 530026 219852 530032 219904
rect 530084 219892 530090 219904
rect 550606 219892 550634 219932
rect 530084 219864 550634 219892
rect 530084 219852 530090 219864
rect 560202 219852 560208 219904
rect 560260 219892 560266 219904
rect 608686 219892 608692 219904
rect 560260 219864 608692 219892
rect 560260 219852 560266 219864
rect 608686 219852 608692 219864
rect 608744 219852 608750 219904
rect 620462 219892 620468 219904
rect 615466 219864 620468 219892
rect 202782 219824 202788 219836
rect 190288 219796 202788 219824
rect 202782 219784 202788 219796
rect 202840 219784 202846 219836
rect 252738 219824 252744 219836
rect 202984 219796 252744 219824
rect 121086 219648 121092 219700
rect 121144 219688 121150 219700
rect 121144 219660 122834 219688
rect 121144 219648 121150 219660
rect 122806 219552 122834 219660
rect 127618 219648 127624 219700
rect 127676 219688 127682 219700
rect 140774 219688 140780 219700
rect 127676 219660 140780 219688
rect 127676 219648 127682 219660
rect 140774 219648 140780 219660
rect 140832 219648 140838 219700
rect 140958 219648 140964 219700
rect 141016 219688 141022 219700
rect 141016 219660 200988 219688
rect 141016 219648 141022 219660
rect 127802 219552 127808 219564
rect 122806 219524 127808 219552
rect 127802 219512 127808 219524
rect 127860 219512 127866 219564
rect 134334 219512 134340 219564
rect 134392 219552 134398 219564
rect 200758 219552 200764 219564
rect 134392 219524 200764 219552
rect 134392 219512 134398 219524
rect 200758 219512 200764 219524
rect 200816 219512 200822 219564
rect 200960 219552 200988 219660
rect 201126 219648 201132 219700
rect 201184 219688 201190 219700
rect 202984 219688 203012 219796
rect 252738 219784 252744 219796
rect 252796 219784 252802 219836
rect 270770 219784 270776 219836
rect 270828 219824 270834 219836
rect 279142 219824 279148 219836
rect 270828 219796 279148 219824
rect 270828 219784 270834 219796
rect 279142 219784 279148 219796
rect 279200 219784 279206 219836
rect 286686 219784 286692 219836
rect 286744 219824 286750 219836
rect 319070 219824 319076 219836
rect 286744 219796 319076 219824
rect 286744 219784 286750 219796
rect 319070 219784 319076 219796
rect 319128 219784 319134 219836
rect 506014 219716 506020 219768
rect 506072 219756 506078 219768
rect 589274 219756 589280 219768
rect 506072 219728 589280 219756
rect 506072 219716 506078 219728
rect 589274 219716 589280 219728
rect 589332 219716 589338 219768
rect 589642 219716 589648 219768
rect 589700 219756 589706 219768
rect 600774 219756 600780 219768
rect 589700 219728 600780 219756
rect 589700 219716 589706 219728
rect 600774 219716 600780 219728
rect 600832 219716 600838 219768
rect 600958 219716 600964 219768
rect 601016 219756 601022 219768
rect 615466 219756 615494 219864
rect 620462 219852 620468 219864
rect 620520 219852 620526 219904
rect 601016 219728 615494 219756
rect 601016 219716 601022 219728
rect 201184 219660 203012 219688
rect 201184 219648 201190 219660
rect 203150 219648 203156 219700
rect 203208 219688 203214 219700
rect 203208 219660 206048 219688
rect 203208 219648 203214 219660
rect 205818 219552 205824 219564
rect 200960 219524 205824 219552
rect 205818 219512 205824 219524
rect 205876 219512 205882 219564
rect 206020 219552 206048 219660
rect 207198 219648 207204 219700
rect 207256 219688 207262 219700
rect 257246 219688 257252 219700
rect 207256 219660 257252 219688
rect 207256 219648 207262 219660
rect 257246 219648 257252 219660
rect 257304 219648 257310 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 527542 219580 527548 219632
rect 527600 219620 527606 219632
rect 619910 219620 619916 219632
rect 527600 219592 619916 219620
rect 527600 219580 527606 219592
rect 619910 219580 619916 219592
rect 619968 219580 619974 219632
rect 208578 219552 208584 219564
rect 206020 219524 208584 219552
rect 208578 219512 208584 219524
rect 208636 219512 208642 219564
rect 212902 219512 212908 219564
rect 212960 219552 212966 219564
rect 215938 219552 215944 219564
rect 212960 219524 215944 219552
rect 212960 219512 212966 219524
rect 215938 219512 215944 219524
rect 215996 219512 216002 219564
rect 289814 219512 289820 219564
rect 289872 219552 289878 219564
rect 289872 219524 290136 219552
rect 289872 219512 289878 219524
rect 105814 219444 105820 219496
rect 105872 219484 105878 219496
rect 105872 219456 106182 219484
rect 105872 219444 105878 219456
rect 63954 219376 63960 219428
rect 64012 219416 64018 219428
rect 64874 219416 64880 219428
rect 64012 219388 64880 219416
rect 64012 219376 64018 219388
rect 64874 219376 64880 219388
rect 64932 219376 64938 219428
rect 106154 219416 106182 219456
rect 221642 219444 221648 219496
rect 221700 219484 221706 219496
rect 221700 219456 223712 219484
rect 221700 219444 221706 219456
rect 147122 219416 147128 219428
rect 106154 219388 147128 219416
rect 147122 219376 147128 219388
rect 147180 219376 147186 219428
rect 159174 219376 159180 219428
rect 159232 219416 159238 219428
rect 160002 219416 160008 219428
rect 159232 219388 160008 219416
rect 159232 219376 159238 219388
rect 160002 219376 160008 219388
rect 160060 219376 160066 219428
rect 163314 219376 163320 219428
rect 163372 219416 163378 219428
rect 163958 219416 163964 219428
rect 163372 219388 163964 219416
rect 163372 219376 163378 219388
rect 163958 219376 163964 219388
rect 164016 219376 164022 219428
rect 204530 219416 204536 219428
rect 166966 219388 204536 219416
rect 106918 219280 106924 219292
rect 64846 219252 106924 219280
rect 63126 219104 63132 219156
rect 63184 219144 63190 219156
rect 64846 219144 64874 219252
rect 106918 219240 106924 219252
rect 106976 219240 106982 219292
rect 113634 219240 113640 219292
rect 113692 219280 113698 219292
rect 156322 219280 156328 219292
rect 113692 219252 156328 219280
rect 113692 219240 113698 219252
rect 156322 219240 156328 219252
rect 156380 219240 156386 219292
rect 160002 219240 160008 219292
rect 160060 219280 160066 219292
rect 166966 219280 166994 219388
rect 204530 219376 204536 219388
rect 204588 219376 204594 219428
rect 209682 219376 209688 219428
rect 209740 219416 209746 219428
rect 210418 219416 210424 219428
rect 209740 219388 210424 219416
rect 209740 219376 209746 219388
rect 210418 219376 210424 219388
rect 210476 219376 210482 219428
rect 217962 219376 217968 219428
rect 218020 219416 218026 219428
rect 223684 219416 223712 219456
rect 258074 219416 258080 219428
rect 218020 219388 219434 219416
rect 223684 219388 258080 219416
rect 218020 219376 218026 219388
rect 160060 219252 166994 219280
rect 160060 219240 160066 219252
rect 167454 219240 167460 219292
rect 167512 219280 167518 219292
rect 168190 219280 168196 219292
rect 167512 219252 168196 219280
rect 167512 219240 167518 219252
rect 168190 219240 168196 219252
rect 168248 219240 168254 219292
rect 169110 219240 169116 219292
rect 169168 219280 169174 219292
rect 169662 219280 169668 219292
rect 169168 219252 169668 219280
rect 169168 219240 169174 219252
rect 169662 219240 169668 219252
rect 169720 219240 169726 219292
rect 169938 219240 169944 219292
rect 169996 219280 170002 219292
rect 171042 219280 171048 219292
rect 169996 219252 171048 219280
rect 169996 219240 170002 219252
rect 171042 219240 171048 219252
rect 171100 219240 171106 219292
rect 172422 219240 172428 219292
rect 172480 219280 172486 219292
rect 173158 219280 173164 219292
rect 172480 219252 173164 219280
rect 172480 219240 172486 219252
rect 173158 219240 173164 219252
rect 173216 219240 173222 219292
rect 182358 219240 182364 219292
rect 182416 219280 182422 219292
rect 189718 219280 189724 219292
rect 182416 219252 189724 219280
rect 182416 219240 182422 219252
rect 189718 219240 189724 219252
rect 189776 219240 189782 219292
rect 192294 219240 192300 219292
rect 192352 219280 192358 219292
rect 192938 219280 192944 219292
rect 192352 219252 192944 219280
rect 192352 219240 192358 219252
rect 192938 219240 192944 219252
rect 192996 219240 193002 219292
rect 193122 219240 193128 219292
rect 193180 219280 193186 219292
rect 198182 219280 198188 219292
rect 193180 219252 198188 219280
rect 193180 219240 193186 219252
rect 198182 219240 198188 219252
rect 198240 219240 198246 219292
rect 198918 219240 198924 219292
rect 198976 219280 198982 219292
rect 200022 219280 200028 219292
rect 198976 219252 200028 219280
rect 198976 219240 198982 219252
rect 200022 219240 200028 219252
rect 200080 219240 200086 219292
rect 201862 219240 201868 219292
rect 201920 219280 201926 219292
rect 207658 219280 207664 219292
rect 201920 219252 207664 219280
rect 201920 219240 201926 219252
rect 207658 219240 207664 219252
rect 207716 219240 207722 219292
rect 211338 219240 211344 219292
rect 211396 219280 211402 219292
rect 218146 219280 218152 219292
rect 211396 219252 218152 219280
rect 211396 219240 211402 219252
rect 218146 219240 218152 219252
rect 218204 219240 218210 219292
rect 219406 219280 219434 219388
rect 258074 219376 258080 219388
rect 258132 219376 258138 219428
rect 272886 219376 272892 219428
rect 272944 219416 272950 219428
rect 290108 219416 290136 219524
rect 366726 219512 366732 219564
rect 366784 219552 366790 219564
rect 432138 219552 432144 219564
rect 366784 219524 367048 219552
rect 366784 219512 366790 219524
rect 367020 219434 367048 219524
rect 429212 219524 432144 219552
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 297542 219416 297548 219428
rect 272944 219388 290044 219416
rect 290108 219388 297548 219416
rect 272944 219376 272950 219388
rect 223482 219280 223488 219292
rect 219406 219252 223488 219280
rect 223482 219240 223488 219252
rect 223540 219240 223546 219292
rect 239490 219240 239496 219292
rect 239548 219280 239554 219292
rect 272702 219280 272708 219292
rect 239548 219252 272708 219280
rect 239548 219240 239554 219252
rect 272702 219240 272708 219252
rect 272760 219240 272766 219292
rect 289814 219280 289820 219292
rect 277366 219252 289820 219280
rect 63184 219116 64874 219144
rect 63184 219104 63190 219116
rect 70578 219104 70584 219156
rect 70636 219144 70642 219156
rect 117958 219144 117964 219156
rect 70636 219116 117964 219144
rect 70636 219104 70642 219116
rect 117958 219104 117964 219116
rect 118016 219104 118022 219156
rect 132586 219104 132592 219156
rect 132644 219144 132650 219156
rect 177482 219144 177488 219156
rect 132644 219116 177488 219144
rect 132644 219104 132650 219116
rect 177482 219104 177488 219116
rect 177540 219104 177546 219156
rect 179046 219104 179052 219156
rect 179104 219144 179110 219156
rect 196618 219144 196624 219156
rect 179104 219116 196624 219144
rect 179104 219104 179110 219116
rect 196618 219104 196624 219116
rect 196676 219104 196682 219156
rect 199746 219104 199752 219156
rect 199804 219144 199810 219156
rect 243538 219144 243544 219156
rect 199804 219116 243544 219144
rect 199804 219104 199810 219116
rect 243538 219104 243544 219116
rect 243596 219104 243602 219156
rect 272334 219104 272340 219156
rect 272392 219144 272398 219156
rect 277366 219144 277394 219252
rect 289814 219240 289820 219252
rect 289872 219240 289878 219292
rect 290016 219280 290044 219388
rect 297542 219376 297548 219388
rect 297600 219376 297606 219428
rect 304074 219376 304080 219428
rect 304132 219416 304138 219428
rect 308398 219416 308404 219428
rect 304132 219388 308404 219416
rect 304132 219376 304138 219388
rect 308398 219376 308404 219388
rect 308456 219376 308462 219428
rect 320634 219376 320640 219428
rect 320692 219416 320698 219428
rect 320692 219388 335354 219416
rect 320692 219376 320698 219388
rect 290016 219252 291884 219280
rect 272392 219116 277394 219144
rect 272392 219104 272398 219116
rect 279050 219104 279056 219156
rect 279108 219144 279114 219156
rect 286318 219144 286324 219156
rect 279108 219116 286324 219144
rect 279108 219104 279114 219116
rect 286318 219104 286324 219116
rect 286376 219104 286382 219156
rect 291856 219144 291884 219252
rect 292022 219240 292028 219292
rect 292080 219280 292086 219292
rect 313918 219280 313924 219292
rect 292080 219252 313924 219280
rect 292080 219240 292086 219252
rect 313918 219240 313924 219252
rect 313976 219240 313982 219292
rect 335326 219280 335354 219388
rect 341334 219376 341340 219428
rect 341392 219416 341398 219428
rect 342254 219416 342260 219428
rect 341392 219388 342260 219416
rect 341392 219376 341398 219388
rect 342254 219376 342260 219388
rect 342312 219376 342318 219428
rect 343818 219376 343824 219428
rect 343876 219416 343882 219428
rect 347038 219416 347044 219428
rect 343876 219388 347044 219416
rect 343876 219376 343882 219388
rect 347038 219376 347044 219388
rect 347096 219376 347102 219428
rect 366174 219376 366180 219428
rect 366232 219416 366238 219428
rect 366928 219416 367048 219434
rect 366232 219406 367048 219416
rect 366232 219388 366956 219406
rect 366232 219376 366238 219388
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 428274 219376 428280 219428
rect 428332 219416 428338 219428
rect 429212 219416 429240 219524
rect 432138 219512 432144 219524
rect 432196 219512 432202 219564
rect 501138 219512 501144 219564
rect 501196 219552 501202 219564
rect 501196 219524 505094 219552
rect 501196 219512 501202 219524
rect 505066 219484 505094 219524
rect 505066 219456 589274 219484
rect 428332 219388 429240 219416
rect 428332 219376 428338 219388
rect 561674 219308 561680 219360
rect 561732 219348 561738 219360
rect 562318 219348 562324 219360
rect 561732 219320 562324 219348
rect 561732 219308 561738 219320
rect 562318 219308 562324 219320
rect 562376 219348 562382 219360
rect 566918 219348 566924 219360
rect 562376 219320 566924 219348
rect 562376 219308 562382 219320
rect 566918 219308 566924 219320
rect 566976 219308 566982 219360
rect 567102 219308 567108 219360
rect 567160 219348 567166 219360
rect 571886 219348 571892 219360
rect 567160 219320 571892 219348
rect 567160 219308 567166 219320
rect 571886 219308 571892 219320
rect 571944 219308 571950 219360
rect 572254 219308 572260 219360
rect 572312 219348 572318 219360
rect 589246 219348 589274 219456
rect 589458 219444 589464 219496
rect 589516 219484 589522 219496
rect 600958 219484 600964 219496
rect 589516 219456 600964 219484
rect 589516 219444 589522 219456
rect 600958 219444 600964 219456
rect 601016 219444 601022 219496
rect 601510 219444 601516 219496
rect 601568 219484 601574 219496
rect 607490 219484 607496 219496
rect 601568 219456 607496 219484
rect 601568 219444 601574 219456
rect 607490 219444 607496 219456
rect 607548 219444 607554 219496
rect 596818 219348 596824 219360
rect 572312 219320 582374 219348
rect 589246 219320 596824 219348
rect 572312 219308 572318 219320
rect 345290 219280 345296 219292
rect 335326 219252 345296 219280
rect 345290 219240 345296 219252
rect 345348 219240 345354 219292
rect 419166 219240 419172 219292
rect 419224 219280 419230 219292
rect 422662 219280 422668 219292
rect 419224 219252 422668 219280
rect 419224 219240 419230 219252
rect 422662 219240 422668 219252
rect 422720 219240 422726 219292
rect 557810 219240 557816 219292
rect 557868 219280 557874 219292
rect 557868 219252 558316 219280
rect 557868 219240 557874 219252
rect 291856 219116 291976 219144
rect 62298 218968 62304 219020
rect 62356 219008 62362 219020
rect 72418 219008 72424 219020
rect 62356 218980 72424 219008
rect 62356 218968 62362 218980
rect 72418 218968 72424 218980
rect 72476 218968 72482 219020
rect 77202 218968 77208 219020
rect 77260 219008 77266 219020
rect 140038 219008 140044 219020
rect 77260 218980 140044 219008
rect 77260 218968 77266 218980
rect 140038 218968 140044 218980
rect 140096 218968 140102 219020
rect 153838 219008 153844 219020
rect 142126 218980 153844 219008
rect 50706 218832 50712 218884
rect 50764 218872 50770 218884
rect 62758 218872 62764 218884
rect 50764 218844 62764 218872
rect 50764 218832 50770 218844
rect 62758 218832 62764 218844
rect 62816 218832 62822 218884
rect 83826 218832 83832 218884
rect 83884 218872 83890 218884
rect 142126 218872 142154 218980
rect 153838 218968 153844 218980
rect 153896 218968 153902 219020
rect 203518 219008 203524 219020
rect 154040 218980 203524 219008
rect 143718 218872 143724 218884
rect 83884 218844 142154 218872
rect 142448 218844 143724 218872
rect 83884 218832 83890 218844
rect 59814 218696 59820 218748
rect 59872 218736 59878 218748
rect 142448 218736 142476 218844
rect 143718 218832 143724 218844
rect 143776 218832 143782 218884
rect 146754 218832 146760 218884
rect 146812 218872 146818 218884
rect 146812 218844 151814 218872
rect 146812 218832 146818 218844
rect 59872 218708 142476 218736
rect 59872 218696 59878 218708
rect 142614 218696 142620 218748
rect 142672 218736 142678 218748
rect 143258 218736 143264 218748
rect 142672 218708 143264 218736
rect 142672 218696 142678 218708
rect 143258 218696 143264 218708
rect 143316 218696 143322 218748
rect 144270 218696 144276 218748
rect 144328 218736 144334 218748
rect 144822 218736 144828 218748
rect 144328 218708 144828 218736
rect 144328 218696 144334 218708
rect 144822 218696 144828 218708
rect 144880 218696 144886 218748
rect 145098 218696 145104 218748
rect 145156 218736 145162 218748
rect 145926 218736 145932 218748
rect 145156 218708 145932 218736
rect 145156 218696 145162 218708
rect 145926 218696 145932 218708
rect 145984 218696 145990 218748
rect 148410 218696 148416 218748
rect 148468 218736 148474 218748
rect 148962 218736 148968 218748
rect 148468 218708 148968 218736
rect 148468 218696 148474 218708
rect 148962 218696 148968 218708
rect 149020 218696 149026 218748
rect 149238 218696 149244 218748
rect 149296 218736 149302 218748
rect 150066 218736 150072 218748
rect 149296 218708 150072 218736
rect 149296 218696 149302 218708
rect 150066 218696 150072 218708
rect 150124 218696 150130 218748
rect 151786 218736 151814 218844
rect 153378 218832 153384 218884
rect 153436 218872 153442 218884
rect 154040 218872 154068 218980
rect 203518 218968 203524 218980
rect 203576 218968 203582 219020
rect 206370 218968 206376 219020
rect 206428 219008 206434 219020
rect 253842 219008 253848 219020
rect 206428 218980 253848 219008
rect 206428 218968 206434 218980
rect 253842 218968 253848 218980
rect 253900 218968 253906 219020
rect 259178 218968 259184 219020
rect 259236 219008 259242 219020
rect 291654 219008 291660 219020
rect 259236 218980 291660 219008
rect 259236 218968 259242 218980
rect 291654 218968 291660 218980
rect 291712 218968 291718 219020
rect 291948 219008 291976 219116
rect 295794 219104 295800 219156
rect 295852 219144 295858 219156
rect 296714 219144 296720 219156
rect 295852 219116 296720 219144
rect 295852 219104 295858 219116
rect 296714 219104 296720 219116
rect 296772 219104 296778 219156
rect 300486 219104 300492 219156
rect 300544 219144 300550 219156
rect 322106 219144 322112 219156
rect 300544 219116 322112 219144
rect 300544 219104 300550 219116
rect 322106 219104 322112 219116
rect 322164 219104 322170 219156
rect 325326 219104 325332 219156
rect 325384 219144 325390 219156
rect 327718 219144 327724 219156
rect 325384 219116 327724 219144
rect 325384 219104 325390 219116
rect 327718 219104 327724 219116
rect 327776 219104 327782 219156
rect 340506 219104 340512 219156
rect 340564 219144 340570 219156
rect 352558 219144 352564 219156
rect 340564 219116 352564 219144
rect 340564 219104 340570 219116
rect 352558 219104 352564 219116
rect 352616 219104 352622 219156
rect 362034 219104 362040 219156
rect 362092 219144 362098 219156
rect 370958 219144 370964 219156
rect 362092 219116 370964 219144
rect 362092 219104 362098 219116
rect 370958 219104 370964 219116
rect 371016 219104 371022 219156
rect 552658 219104 552664 219156
rect 552716 219144 552722 219156
rect 558288 219144 558316 219252
rect 572088 219184 572714 219212
rect 552716 219116 558224 219144
rect 558288 219116 567332 219144
rect 552716 219104 552722 219116
rect 297358 219008 297364 219020
rect 291948 218980 297364 219008
rect 297358 218968 297364 218980
rect 297416 218968 297422 219020
rect 307386 218968 307392 219020
rect 307444 219008 307450 219020
rect 331858 219008 331864 219020
rect 307444 218980 331864 219008
rect 307444 218968 307450 218980
rect 331858 218968 331864 218980
rect 331916 218968 331922 219020
rect 333698 218968 333704 219020
rect 333756 219008 333762 219020
rect 355226 219008 355232 219020
rect 333756 218980 355232 219008
rect 333756 218968 333762 218980
rect 355226 218968 355232 218980
rect 355284 218968 355290 219020
rect 357066 218968 357072 219020
rect 357124 219008 357130 219020
rect 369118 219008 369124 219020
rect 357124 218980 369124 219008
rect 357124 218968 357130 218980
rect 369118 218968 369124 218980
rect 369176 218968 369182 219020
rect 370314 218968 370320 219020
rect 370372 219008 370378 219020
rect 380066 219008 380072 219020
rect 370372 218980 380072 219008
rect 370372 218968 370378 218980
rect 380066 218968 380072 218980
rect 380124 218968 380130 219020
rect 380250 218968 380256 219020
rect 380308 219008 380314 219020
rect 388622 219008 388628 219020
rect 380308 218980 388628 219008
rect 380308 218968 380314 218980
rect 388622 218968 388628 218980
rect 388680 218968 388686 219020
rect 547414 218968 547420 219020
rect 547472 219008 547478 219020
rect 557626 219008 557632 219020
rect 547472 218980 557632 219008
rect 547472 218968 547478 218980
rect 557626 218968 557632 218980
rect 557684 218968 557690 219020
rect 558196 219008 558224 219116
rect 567102 219008 567108 219020
rect 558196 218980 567108 219008
rect 567102 218968 567108 218980
rect 567160 218968 567166 219020
rect 153436 218844 154068 218872
rect 153436 218832 153442 218844
rect 156322 218832 156328 218884
rect 156380 218872 156386 218884
rect 162302 218872 162308 218884
rect 156380 218844 162308 218872
rect 156380 218832 156386 218844
rect 162302 218832 162308 218844
rect 162360 218832 162366 218884
rect 162486 218832 162492 218884
rect 162544 218872 162550 218884
rect 171594 218872 171600 218884
rect 162544 218844 171600 218872
rect 162544 218832 162550 218844
rect 171594 218832 171600 218844
rect 171652 218832 171658 218884
rect 180058 218872 180064 218884
rect 171796 218844 180064 218872
rect 151786 218708 162164 218736
rect 100386 218560 100392 218612
rect 100444 218600 100450 218612
rect 105814 218600 105820 218612
rect 100444 218572 105820 218600
rect 100444 218560 100450 218572
rect 105814 218560 105820 218572
rect 105872 218560 105878 218612
rect 120258 218560 120264 218612
rect 120316 218600 120322 218612
rect 162136 218600 162164 218708
rect 165798 218696 165804 218748
rect 165856 218736 165862 218748
rect 171796 218736 171824 218844
rect 180058 218832 180064 218844
rect 180116 218832 180122 218884
rect 180766 218844 184796 218872
rect 165856 218708 171824 218736
rect 165856 218696 165862 218708
rect 175734 218696 175740 218748
rect 175792 218736 175798 218748
rect 180766 218736 180794 218844
rect 175792 218708 180794 218736
rect 175792 218696 175798 218708
rect 181162 218696 181168 218748
rect 181220 218736 181226 218748
rect 184382 218736 184388 218748
rect 181220 218708 184388 218736
rect 181220 218696 181226 218708
rect 184382 218696 184388 218708
rect 184440 218696 184446 218748
rect 184768 218736 184796 218844
rect 188982 218832 188988 218884
rect 189040 218872 189046 218884
rect 194134 218872 194140 218884
rect 189040 218844 194140 218872
rect 189040 218832 189046 218844
rect 194134 218832 194140 218844
rect 194192 218832 194198 218884
rect 194318 218832 194324 218884
rect 194376 218872 194382 218884
rect 239306 218872 239312 218884
rect 194376 218844 239312 218872
rect 194376 218832 194382 218844
rect 239306 218832 239312 218844
rect 239364 218832 239370 218884
rect 246114 218832 246120 218884
rect 246172 218872 246178 218884
rect 279050 218872 279056 218884
rect 246172 218844 279056 218872
rect 246172 218832 246178 218844
rect 279050 218832 279056 218844
rect 279108 218832 279114 218884
rect 279234 218832 279240 218884
rect 279292 218872 279298 218884
rect 279292 218844 282316 218872
rect 279292 218832 279298 218844
rect 189626 218736 189632 218748
rect 184768 218708 189632 218736
rect 189626 218696 189632 218708
rect 189684 218696 189690 218748
rect 189810 218696 189816 218748
rect 189868 218736 189874 218748
rect 195422 218736 195428 218748
rect 189868 218708 195428 218736
rect 189868 218696 189874 218708
rect 195422 218696 195428 218708
rect 195480 218696 195486 218748
rect 195606 218696 195612 218748
rect 195664 218736 195670 218748
rect 197998 218736 198004 218748
rect 195664 218708 198004 218736
rect 195664 218696 195670 218708
rect 197998 218696 198004 218708
rect 198056 218696 198062 218748
rect 198182 218696 198188 218748
rect 198240 218736 198246 218748
rect 246298 218736 246304 218748
rect 198240 218708 246304 218736
rect 198240 218696 198246 218708
rect 246298 218696 246304 218708
rect 246356 218696 246362 218748
rect 252738 218696 252744 218748
rect 252796 218736 252802 218748
rect 252796 218708 282224 218736
rect 252796 218696 252802 218708
rect 171042 218600 171048 218612
rect 120316 218572 162072 218600
rect 162136 218572 171048 218600
rect 120316 218560 120322 218572
rect 107010 218424 107016 218476
rect 107068 218464 107074 218476
rect 152366 218464 152372 218476
rect 107068 218436 152372 218464
rect 107068 218424 107074 218436
rect 152366 218424 152372 218436
rect 152424 218424 152430 218476
rect 152550 218424 152556 218476
rect 152608 218464 152614 218476
rect 153102 218464 153108 218476
rect 152608 218436 153108 218464
rect 152608 218424 152614 218436
rect 153102 218424 153108 218436
rect 153160 218424 153166 218476
rect 156690 218424 156696 218476
rect 156748 218464 156754 218476
rect 157242 218464 157248 218476
rect 156748 218436 157248 218464
rect 156748 218424 156754 218436
rect 157242 218424 157248 218436
rect 157300 218424 157306 218476
rect 162044 218464 162072 218572
rect 171042 218560 171048 218572
rect 171100 218560 171106 218612
rect 171594 218560 171600 218612
rect 171652 218600 171658 218612
rect 181346 218600 181352 218612
rect 171652 218572 181352 218600
rect 171652 218560 171658 218572
rect 181346 218560 181352 218572
rect 181404 218560 181410 218612
rect 186498 218560 186504 218612
rect 186556 218600 186562 218612
rect 194318 218600 194324 218612
rect 186556 218572 194324 218600
rect 186556 218560 186562 218572
rect 194318 218560 194324 218572
rect 194376 218560 194382 218612
rect 198090 218560 198096 218612
rect 198148 218600 198154 218612
rect 200390 218600 200396 218612
rect 198148 218572 200396 218600
rect 198148 218560 198154 218572
rect 200390 218560 200396 218572
rect 200448 218560 200454 218612
rect 203058 218560 203064 218612
rect 203116 218600 203122 218612
rect 206186 218600 206192 218612
rect 203116 218572 206192 218600
rect 203116 218560 203122 218572
rect 206186 218560 206192 218572
rect 206244 218560 206250 218612
rect 208026 218560 208032 218612
rect 208084 218600 208090 218612
rect 211522 218600 211528 218612
rect 208084 218572 211528 218600
rect 208084 218560 208090 218572
rect 211522 218560 211528 218572
rect 211580 218560 211586 218612
rect 217318 218600 217324 218612
rect 211724 218572 217324 218600
rect 165614 218464 165620 218476
rect 162044 218436 165620 218464
rect 165614 218424 165620 218436
rect 165672 218424 165678 218476
rect 166626 218424 166632 218476
rect 166684 218464 166690 218476
rect 201862 218464 201868 218476
rect 166684 218436 201868 218464
rect 166684 218424 166690 218436
rect 201862 218424 201868 218436
rect 201920 218424 201926 218476
rect 211724 218464 211752 218572
rect 217318 218560 217324 218572
rect 217376 218560 217382 218612
rect 219618 218560 219624 218612
rect 219676 218600 219682 218612
rect 264606 218600 264612 218612
rect 219676 218572 264612 218600
rect 219676 218560 219682 218572
rect 264606 218560 264612 218572
rect 264664 218560 264670 218612
rect 265986 218560 265992 218612
rect 266044 218600 266050 218612
rect 272334 218600 272340 218612
rect 266044 218572 272340 218600
rect 266044 218560 266050 218572
rect 272334 218560 272340 218572
rect 272392 218560 272398 218612
rect 272702 218560 272708 218612
rect 272760 218600 272766 218612
rect 279418 218600 279424 218612
rect 272760 218572 279424 218600
rect 272760 218560 272766 218572
rect 279418 218560 279424 218572
rect 279476 218560 279482 218612
rect 202064 218436 211752 218464
rect 117958 218288 117964 218340
rect 118016 218328 118022 218340
rect 123478 218328 123484 218340
rect 118016 218300 123484 218328
rect 118016 218288 118022 218300
rect 123478 218288 123484 218300
rect 123536 218288 123542 218340
rect 131850 218288 131856 218340
rect 131908 218328 131914 218340
rect 132402 218328 132408 218340
rect 131908 218300 132408 218328
rect 131908 218288 131914 218300
rect 132402 218288 132408 218300
rect 132460 218288 132466 218340
rect 136818 218288 136824 218340
rect 136876 218328 136882 218340
rect 139486 218328 139492 218340
rect 136876 218300 139492 218328
rect 136876 218288 136882 218300
rect 139486 218288 139492 218300
rect 139544 218288 139550 218340
rect 140130 218288 140136 218340
rect 140188 218328 140194 218340
rect 181162 218328 181168 218340
rect 140188 218300 181168 218328
rect 140188 218288 140194 218300
rect 181162 218288 181168 218300
rect 181220 218288 181226 218340
rect 181530 218288 181536 218340
rect 181588 218328 181594 218340
rect 181990 218328 181996 218340
rect 181588 218300 181996 218328
rect 181588 218288 181594 218300
rect 181990 218288 181996 218300
rect 182048 218288 182054 218340
rect 184014 218288 184020 218340
rect 184072 218328 184078 218340
rect 184934 218328 184940 218340
rect 184072 218300 184940 218328
rect 184072 218288 184078 218300
rect 184934 218288 184940 218300
rect 184992 218288 184998 218340
rect 185670 218288 185676 218340
rect 185728 218328 185734 218340
rect 186130 218328 186136 218340
rect 185728 218300 186136 218328
rect 185728 218288 185734 218300
rect 186130 218288 186136 218300
rect 186188 218288 186194 218340
rect 196434 218288 196440 218340
rect 196492 218328 196498 218340
rect 202064 218328 202092 218436
rect 212994 218424 213000 218476
rect 213052 218464 213058 218476
rect 221642 218464 221648 218476
rect 213052 218436 221648 218464
rect 213052 218424 213058 218436
rect 221642 218424 221648 218436
rect 221700 218424 221706 218476
rect 225966 218424 225972 218476
rect 226024 218464 226030 218476
rect 266998 218464 267004 218476
rect 226024 218436 267004 218464
rect 226024 218424 226030 218436
rect 266998 218424 267004 218436
rect 267056 218424 267062 218476
rect 282196 218464 282224 218708
rect 282288 218600 282316 218844
rect 285858 218832 285864 218884
rect 285916 218872 285922 218884
rect 292022 218872 292028 218884
rect 285916 218844 292028 218872
rect 285916 218832 285922 218844
rect 292022 218832 292028 218844
rect 292080 218832 292086 218884
rect 314010 218832 314016 218884
rect 314068 218872 314074 218884
rect 340046 218872 340052 218884
rect 314068 218844 340052 218872
rect 314068 218832 314074 218844
rect 340046 218832 340052 218844
rect 340104 218832 340110 218884
rect 347038 218832 347044 218884
rect 347096 218872 347102 218884
rect 363506 218872 363512 218884
rect 347096 218844 363512 218872
rect 347096 218832 347102 218844
rect 363506 218832 363512 218844
rect 363564 218832 363570 218884
rect 368658 218832 368664 218884
rect 368716 218872 368722 218884
rect 378778 218872 378784 218884
rect 368716 218844 378784 218872
rect 368716 218832 368722 218844
rect 378778 218832 378784 218844
rect 378836 218832 378842 218884
rect 382734 218832 382740 218884
rect 382792 218872 382798 218884
rect 383562 218872 383568 218884
rect 382792 218844 383568 218872
rect 382792 218832 382798 218844
rect 383562 218832 383568 218844
rect 383620 218832 383626 218884
rect 386874 218832 386880 218884
rect 386932 218872 386938 218884
rect 398098 218872 398104 218884
rect 386932 218844 398104 218872
rect 386932 218832 386938 218844
rect 398098 218832 398104 218844
rect 398156 218832 398162 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412542 218872 412548 218884
rect 411772 218844 412548 218872
rect 411772 218832 411778 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 557994 218872 558000 218884
rect 543706 218844 558000 218872
rect 291654 218696 291660 218748
rect 291712 218736 291718 218748
rect 324590 218736 324596 218748
rect 291712 218708 324596 218736
rect 291712 218696 291718 218708
rect 324590 218696 324596 218708
rect 324648 218696 324654 218748
rect 327258 218696 327264 218748
rect 327316 218736 327322 218748
rect 351086 218736 351092 218748
rect 327316 218708 351092 218736
rect 327316 218696 327322 218708
rect 351086 218696 351092 218708
rect 351144 218696 351150 218748
rect 353754 218696 353760 218748
rect 353812 218736 353818 218748
rect 371786 218736 371792 218748
rect 353812 218708 371792 218736
rect 353812 218696 353818 218708
rect 371786 218696 371792 218708
rect 371844 218696 371850 218748
rect 383562 218696 383568 218748
rect 383620 218736 383626 218748
rect 396258 218736 396264 218748
rect 383620 218708 396264 218736
rect 383620 218696 383626 218708
rect 396258 218696 396264 218708
rect 396316 218696 396322 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 471330 218696 471336 218748
rect 471388 218736 471394 218748
rect 472894 218736 472900 218748
rect 471388 218708 472900 218736
rect 471388 218696 471394 218708
rect 472894 218696 472900 218708
rect 472952 218696 472958 218748
rect 482738 218696 482744 218748
rect 482796 218736 482802 218748
rect 485314 218736 485320 218748
rect 482796 218708 485320 218736
rect 482796 218696 482802 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 542814 218696 542820 218748
rect 542872 218736 542878 218748
rect 542872 218708 543136 218736
rect 542872 218696 542878 218708
rect 304258 218600 304264 218612
rect 282288 218572 304264 218600
rect 304258 218560 304264 218572
rect 304316 218560 304322 218612
rect 398466 218560 398472 218612
rect 398524 218600 398530 218612
rect 407758 218600 407764 218612
rect 398524 218572 407764 218600
rect 398524 218560 398530 218572
rect 407758 218560 407764 218572
rect 407816 218560 407822 218612
rect 429930 218560 429936 218612
rect 429988 218600 429994 218612
rect 432138 218600 432144 218612
rect 429988 218572 432144 218600
rect 429988 218560 429994 218572
rect 432138 218560 432144 218572
rect 432196 218560 432202 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 537478 218560 537484 218612
rect 537536 218600 537542 218612
rect 543108 218600 543136 218708
rect 543706 218600 543734 218844
rect 557994 218832 558000 218844
rect 558052 218832 558058 218884
rect 566734 218872 566740 218884
rect 558196 218844 566740 218872
rect 548518 218696 548524 218748
rect 548576 218736 548582 218748
rect 558196 218736 558224 218844
rect 566734 218832 566740 218844
rect 566792 218832 566798 218884
rect 567304 218872 567332 219116
rect 567470 219104 567476 219156
rect 567528 219144 567534 219156
rect 572088 219144 572116 219184
rect 567528 219116 572116 219144
rect 572686 219144 572714 219184
rect 574278 219144 574284 219156
rect 572686 219116 574284 219144
rect 567528 219104 567534 219116
rect 574278 219104 574284 219116
rect 574336 219104 574342 219156
rect 567654 218968 567660 219020
rect 567712 219008 567718 219020
rect 575474 219008 575480 219020
rect 567712 218980 575480 219008
rect 567712 218968 567718 218980
rect 575474 218968 575480 218980
rect 575532 218968 575538 219020
rect 567304 218844 567976 218872
rect 548576 218708 558224 218736
rect 558288 218708 567884 218736
rect 548576 218696 548582 218708
rect 537536 218572 543044 218600
rect 543108 218572 543734 218600
rect 537536 218560 537542 218572
rect 288986 218464 288992 218476
rect 282196 218436 288992 218464
rect 288986 218424 288992 218436
rect 289044 218424 289050 218476
rect 294138 218424 294144 218476
rect 294196 218464 294202 218476
rect 316678 218464 316684 218476
rect 294196 218436 316684 218464
rect 294196 218424 294202 218436
rect 316678 218424 316684 218436
rect 316736 218424 316742 218476
rect 512730 218424 512736 218476
rect 512788 218464 512794 218476
rect 542814 218464 542820 218476
rect 512788 218436 542820 218464
rect 512788 218424 512794 218436
rect 542814 218424 542820 218436
rect 542872 218424 542878 218476
rect 543016 218464 543044 218572
rect 545022 218560 545028 218612
rect 545080 218600 545086 218612
rect 557810 218600 557816 218612
rect 545080 218572 557816 218600
rect 545080 218560 545086 218572
rect 557810 218560 557816 218572
rect 557868 218560 557874 218612
rect 557994 218560 558000 218612
rect 558052 218600 558058 218612
rect 558288 218600 558316 218708
rect 558052 218572 558316 218600
rect 558052 218560 558058 218572
rect 560202 218560 560208 218612
rect 560260 218600 560266 218612
rect 567470 218600 567476 218612
rect 560260 218572 567476 218600
rect 560260 218560 560266 218572
rect 567470 218560 567476 218572
rect 567528 218560 567534 218612
rect 567654 218464 567660 218476
rect 543016 218436 567660 218464
rect 567654 218424 567660 218436
rect 567712 218424 567718 218476
rect 567856 218464 567884 218708
rect 567948 218600 567976 218844
rect 568298 218832 568304 218884
rect 568356 218872 568362 218884
rect 572070 218872 572076 218884
rect 568356 218844 572076 218872
rect 568356 218832 568362 218844
rect 572070 218832 572076 218844
rect 572128 218832 572134 218884
rect 572530 218832 572536 218884
rect 572588 218832 572594 218884
rect 572714 218832 572720 218884
rect 572772 218872 572778 218884
rect 574462 218872 574468 218884
rect 572772 218844 574468 218872
rect 572772 218832 572778 218844
rect 574462 218832 574468 218844
rect 574520 218832 574526 218884
rect 582346 218872 582374 219320
rect 596818 219308 596824 219320
rect 596876 219308 596882 219360
rect 589274 219172 589280 219224
rect 589332 219212 589338 219224
rect 597922 219212 597928 219224
rect 589332 219184 597928 219212
rect 589332 219172 589338 219184
rect 597922 219172 597928 219184
rect 597980 219172 597986 219224
rect 626350 218872 626356 218884
rect 582346 218844 626356 218872
rect 626350 218832 626356 218844
rect 626408 218832 626414 218884
rect 568482 218696 568488 218748
rect 568540 218736 568546 218748
rect 572254 218736 572260 218748
rect 568540 218708 572260 218736
rect 568540 218696 568546 218708
rect 572254 218696 572260 218708
rect 572312 218696 572318 218748
rect 572548 218736 572576 218832
rect 601878 218736 601884 218748
rect 572548 218708 601884 218736
rect 601878 218696 601884 218708
rect 601936 218696 601942 218748
rect 598750 218600 598756 218612
rect 567948 218572 598756 218600
rect 598750 218560 598756 218572
rect 598808 218560 598814 218612
rect 604454 218464 604460 218476
rect 567856 218436 604460 218464
rect 604454 218424 604460 218436
rect 604512 218424 604518 218476
rect 458174 218356 458180 218408
rect 458232 218396 458238 218408
rect 458232 218368 460934 218396
rect 458232 218356 458238 218368
rect 196492 218300 202092 218328
rect 196492 218288 196498 218300
rect 202230 218288 202236 218340
rect 202288 218328 202294 218340
rect 202782 218328 202788 218340
rect 202288 218300 202788 218328
rect 202288 218288 202294 218300
rect 202782 218288 202788 218300
rect 202840 218288 202846 218340
rect 204714 218288 204720 218340
rect 204772 218328 204778 218340
rect 207842 218328 207848 218340
rect 204772 218300 207848 218328
rect 204772 218288 204778 218300
rect 207842 218288 207848 218300
rect 207900 218288 207906 218340
rect 208854 218288 208860 218340
rect 208912 218328 208918 218340
rect 209498 218328 209504 218340
rect 208912 218300 209504 218328
rect 208912 218288 208918 218300
rect 209498 218288 209504 218300
rect 209556 218288 209562 218340
rect 210326 218288 210332 218340
rect 210384 218328 210390 218340
rect 213178 218328 213184 218340
rect 210384 218300 213184 218328
rect 210384 218288 210390 218300
rect 213178 218288 213184 218300
rect 213236 218288 213242 218340
rect 222930 218288 222936 218340
rect 222988 218328 222994 218340
rect 231026 218328 231032 218340
rect 222988 218300 231032 218328
rect 222988 218288 222994 218300
rect 231026 218288 231032 218300
rect 231084 218288 231090 218340
rect 232866 218288 232872 218340
rect 232924 218328 232930 218340
rect 270770 218328 270776 218340
rect 232924 218300 270776 218328
rect 232924 218288 232930 218300
rect 270770 218288 270776 218300
rect 270828 218288 270834 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429378 218328 429384 218340
rect 426676 218300 429384 218328
rect 426676 218288 426682 218300
rect 429378 218288 429384 218300
rect 429436 218288 429442 218340
rect 434898 218288 434904 218340
rect 434956 218328 434962 218340
rect 436646 218328 436652 218340
rect 434956 218300 436652 218328
rect 434956 218288 434962 218300
rect 436646 218288 436652 218300
rect 436704 218288 436710 218340
rect 450722 218288 450728 218340
rect 450780 218328 450786 218340
rect 453850 218328 453856 218340
rect 450780 218300 453856 218328
rect 450780 218288 450786 218300
rect 453850 218288 453856 218300
rect 453908 218288 453914 218340
rect 460906 218328 460934 218368
rect 461302 218328 461308 218340
rect 460906 218300 461308 218328
rect 461302 218288 461308 218300
rect 461360 218288 461366 218340
rect 500402 218288 500408 218340
rect 500460 218328 500466 218340
rect 609882 218328 609888 218340
rect 500460 218300 609888 218328
rect 500460 218288 500466 218300
rect 609882 218288 609888 218300
rect 609940 218288 609946 218340
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 56502 218192 56508 218204
rect 55732 218164 56508 218192
rect 55732 218152 55738 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 57422 218152 57428 218204
rect 57480 218192 57486 218204
rect 61654 218192 61660 218204
rect 57480 218164 61660 218192
rect 57480 218152 57486 218164
rect 61654 218152 61660 218164
rect 61712 218152 61718 218204
rect 67266 218152 67272 218204
rect 67324 218192 67330 218204
rect 68278 218192 68284 218204
rect 67324 218164 68284 218192
rect 67324 218152 67330 218164
rect 68278 218152 68284 218164
rect 68336 218152 68342 218204
rect 75546 218152 75552 218204
rect 75604 218192 75610 218204
rect 76558 218192 76564 218204
rect 75604 218164 76564 218192
rect 75604 218152 75610 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 123570 218152 123576 218204
rect 123628 218192 123634 218204
rect 165982 218192 165988 218204
rect 123628 218164 165988 218192
rect 123628 218152 123634 218164
rect 165982 218152 165988 218164
rect 166040 218152 166046 218204
rect 171410 218192 171416 218204
rect 166966 218164 171416 218192
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59354 218056 59360 218068
rect 58216 218028 59360 218056
rect 58216 218016 58222 218028
rect 59354 218016 59360 218028
rect 59412 218016 59418 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62022 218056 62028 218068
rect 61528 218028 62028 218056
rect 61528 218016 61534 218028
rect 62022 218016 62028 218028
rect 62080 218016 62086 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 66438 218016 66444 218068
rect 66496 218056 66502 218068
rect 67542 218056 67548 218068
rect 66496 218028 67548 218056
rect 66496 218016 66502 218028
rect 67542 218016 67548 218028
rect 67600 218016 67606 218068
rect 68094 218016 68100 218068
rect 68152 218056 68158 218068
rect 68738 218056 68744 218068
rect 68152 218028 68744 218056
rect 68152 218016 68158 218028
rect 68738 218016 68744 218028
rect 68796 218016 68802 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 83458 218056 83464 218068
rect 82228 218028 83464 218056
rect 82228 218016 82234 218028
rect 83458 218016 83464 218028
rect 83516 218016 83522 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85298 218056 85304 218068
rect 84712 218028 85304 218056
rect 84712 218016 84718 218028
rect 85298 218016 85304 218028
rect 85356 218016 85362 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 90450 218016 90456 218068
rect 90508 218056 90514 218068
rect 91738 218056 91744 218068
rect 90508 218028 91744 218056
rect 90508 218016 90514 218028
rect 91738 218016 91744 218028
rect 91796 218016 91802 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93762 218056 93768 218068
rect 92992 218028 93768 218056
rect 92992 218016 92998 218028
rect 93762 218016 93768 218028
rect 93820 218016 93826 218068
rect 95418 218016 95424 218068
rect 95476 218056 95482 218068
rect 96246 218056 96252 218068
rect 95476 218028 96252 218056
rect 95476 218016 95482 218028
rect 96246 218016 96252 218028
rect 96304 218016 96310 218068
rect 97074 218016 97080 218068
rect 97132 218056 97138 218068
rect 97994 218056 98000 218068
rect 97132 218028 98000 218056
rect 97132 218016 97138 218028
rect 97994 218016 98000 218028
rect 98052 218016 98058 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 102870 218016 102876 218068
rect 102928 218056 102934 218068
rect 103422 218056 103428 218068
rect 102928 218028 103428 218056
rect 102928 218016 102934 218028
rect 103422 218016 103428 218028
rect 103480 218016 103486 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 105998 218056 106004 218068
rect 105412 218028 106004 218056
rect 105412 218016 105418 218028
rect 105998 218016 106004 218028
rect 106056 218016 106062 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110138 218056 110144 218068
rect 109552 218028 110144 218056
rect 109552 218016 109558 218028
rect 110138 218016 110144 218028
rect 110196 218016 110202 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 117222 218056 117228 218068
rect 116176 218028 117228 218056
rect 116176 218016 116182 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 117774 218016 117780 218068
rect 117832 218056 117838 218068
rect 118694 218056 118700 218068
rect 117832 218028 118700 218056
rect 117832 218016 117838 218028
rect 118694 218016 118700 218028
rect 118752 218016 118758 218068
rect 119430 218016 119436 218068
rect 119488 218056 119494 218068
rect 119982 218056 119988 218068
rect 119488 218028 119988 218056
rect 119488 218016 119494 218028
rect 119982 218016 119988 218028
rect 120040 218016 120046 218068
rect 121914 218016 121920 218068
rect 121972 218056 121978 218068
rect 122558 218056 122564 218068
rect 121972 218028 122564 218056
rect 121972 218016 121978 218028
rect 122558 218016 122564 218028
rect 122616 218016 122622 218068
rect 126054 218016 126060 218068
rect 126112 218056 126118 218068
rect 126698 218056 126704 218068
rect 126112 218028 126704 218056
rect 126112 218016 126118 218028
rect 126698 218016 126704 218028
rect 126756 218016 126762 218068
rect 127710 218016 127716 218068
rect 127768 218056 127774 218068
rect 128262 218056 128268 218068
rect 127768 218028 128268 218056
rect 127768 218016 127774 218028
rect 128262 218016 128268 218028
rect 128320 218016 128326 218068
rect 128538 218016 128544 218068
rect 128596 218056 128602 218068
rect 129366 218056 129372 218068
rect 128596 218028 129372 218056
rect 128596 218016 128602 218028
rect 129366 218016 129372 218028
rect 129424 218016 129430 218068
rect 130194 218016 130200 218068
rect 130252 218056 130258 218068
rect 132494 218056 132500 218068
rect 130252 218028 132500 218056
rect 130252 218016 130258 218028
rect 132494 218016 132500 218028
rect 132552 218016 132558 218068
rect 132678 218016 132684 218068
rect 132736 218056 132742 218068
rect 133506 218056 133512 218068
rect 132736 218028 133512 218056
rect 132736 218016 132742 218028
rect 133506 218016 133512 218028
rect 133564 218016 133570 218068
rect 135990 218016 135996 218068
rect 136048 218056 136054 218068
rect 136542 218056 136548 218068
rect 136048 218028 136548 218056
rect 136048 218016 136054 218028
rect 136542 218016 136548 218028
rect 136600 218016 136606 218068
rect 138474 218016 138480 218068
rect 138532 218056 138538 218068
rect 139118 218056 139124 218068
rect 138532 218028 139124 218056
rect 138532 218016 138538 218028
rect 139118 218016 139124 218028
rect 139176 218016 139182 218068
rect 139486 218016 139492 218068
rect 139544 218056 139550 218068
rect 166966 218056 166994 218164
rect 171410 218152 171416 218164
rect 171468 218152 171474 218204
rect 173250 218152 173256 218204
rect 173308 218192 173314 218204
rect 173308 218164 179552 218192
rect 173308 218152 173314 218164
rect 139544 218028 166994 218056
rect 139544 218016 139550 218028
rect 170766 218016 170772 218068
rect 170824 218056 170830 218068
rect 176470 218056 176476 218068
rect 170824 218028 176476 218056
rect 170824 218016 170830 218028
rect 176470 218016 176476 218028
rect 176528 218016 176534 218068
rect 178218 218016 178224 218068
rect 178276 218056 178282 218068
rect 179322 218056 179328 218068
rect 178276 218028 179328 218056
rect 178276 218016 178282 218028
rect 179322 218016 179328 218028
rect 179380 218016 179386 218068
rect 179524 218056 179552 218164
rect 179874 218152 179880 218204
rect 179932 218192 179938 218204
rect 225598 218192 225604 218204
rect 179932 218164 225604 218192
rect 179932 218152 179938 218164
rect 225598 218152 225604 218164
rect 225656 218152 225662 218204
rect 241974 218152 241980 218204
rect 242032 218192 242038 218204
rect 242894 218192 242900 218204
rect 242032 218164 242900 218192
rect 242032 218152 242038 218164
rect 242894 218152 242900 218164
rect 242952 218152 242958 218204
rect 243538 218152 243544 218204
rect 243596 218192 243602 218204
rect 249058 218192 249064 218204
rect 243596 218164 249064 218192
rect 243596 218152 243602 218164
rect 249058 218152 249064 218164
rect 249116 218152 249122 218204
rect 297450 218152 297456 218204
rect 297508 218192 297514 218204
rect 302878 218192 302884 218204
rect 297508 218164 302884 218192
rect 297508 218152 297514 218164
rect 302878 218152 302884 218164
rect 302936 218152 302942 218204
rect 335538 218152 335544 218204
rect 335596 218192 335602 218204
rect 338666 218192 338672 218204
rect 335596 218164 338672 218192
rect 335596 218152 335602 218164
rect 338666 218152 338672 218164
rect 338724 218152 338730 218204
rect 358722 218152 358728 218204
rect 358780 218192 358786 218204
rect 359458 218192 359464 218204
rect 358780 218164 359464 218192
rect 358780 218152 358786 218164
rect 359458 218152 359464 218164
rect 359516 218152 359522 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 400950 218152 400956 218204
rect 401008 218192 401014 218204
rect 402238 218192 402244 218204
rect 401008 218164 402244 218192
rect 401008 218152 401014 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 427906 218192 427912 218204
rect 425848 218164 427912 218192
rect 425848 218152 425854 218164
rect 427906 218152 427912 218164
rect 427964 218152 427970 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 502978 218152 502984 218204
rect 503036 218192 503042 218204
rect 548518 218192 548524 218204
rect 503036 218164 548524 218192
rect 503036 218152 503042 218164
rect 548518 218152 548524 218164
rect 548576 218152 548582 218204
rect 553394 218152 553400 218204
rect 553452 218192 553458 218204
rect 556522 218192 556528 218204
rect 553452 218164 556528 218192
rect 553452 218152 553458 218164
rect 556522 218152 556528 218164
rect 556580 218152 556586 218204
rect 557626 218152 557632 218204
rect 557684 218192 557690 218204
rect 560202 218192 560208 218204
rect 557684 218164 560208 218192
rect 557684 218152 557690 218164
rect 560202 218152 560208 218164
rect 560260 218152 560266 218204
rect 562134 218152 562140 218204
rect 562192 218192 562198 218204
rect 563054 218192 563060 218204
rect 562192 218164 563060 218192
rect 562192 218152 562198 218164
rect 563054 218152 563060 218164
rect 563112 218152 563118 218204
rect 572438 218152 572444 218204
rect 572496 218192 572502 218204
rect 614482 218192 614488 218204
rect 572496 218164 614488 218192
rect 572496 218152 572502 218164
rect 614482 218152 614488 218164
rect 614540 218152 614546 218204
rect 563348 218096 572300 218124
rect 210326 218056 210332 218068
rect 179524 218028 210332 218056
rect 210326 218016 210332 218028
rect 210384 218016 210390 218068
rect 210510 218016 210516 218068
rect 210568 218056 210574 218068
rect 210970 218056 210976 218068
rect 210568 218028 210976 218056
rect 210568 218016 210574 218028
rect 210970 218016 210976 218028
rect 211028 218016 211034 218068
rect 214650 218016 214656 218068
rect 214708 218056 214714 218068
rect 215202 218056 215208 218068
rect 214708 218028 215208 218056
rect 214708 218016 214714 218028
rect 215202 218016 215208 218028
rect 215260 218016 215266 218068
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216122 218056 216128 218068
rect 215536 218028 216128 218056
rect 215536 218016 215542 218028
rect 216122 218016 216128 218028
rect 216180 218016 216186 218068
rect 218790 218016 218796 218068
rect 218848 218056 218854 218068
rect 219342 218056 219348 218068
rect 218848 218028 219348 218056
rect 218848 218016 218854 218028
rect 219342 218016 219348 218028
rect 219400 218016 219406 218068
rect 221274 218016 221280 218068
rect 221332 218056 221338 218068
rect 221826 218056 221832 218068
rect 221332 218028 221832 218056
rect 221332 218016 221338 218028
rect 221826 218016 221832 218028
rect 221884 218016 221890 218068
rect 225414 218016 225420 218068
rect 225472 218056 225478 218068
rect 226150 218056 226156 218068
rect 225472 218028 226156 218056
rect 225472 218016 225478 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 227070 218016 227076 218068
rect 227128 218056 227134 218068
rect 227530 218056 227536 218068
rect 227128 218028 227536 218056
rect 227128 218016 227134 218028
rect 227530 218016 227536 218028
rect 227588 218016 227594 218068
rect 229554 218016 229560 218068
rect 229612 218056 229618 218068
rect 230474 218056 230480 218068
rect 229612 218028 230480 218056
rect 229612 218016 229618 218028
rect 230474 218016 230480 218028
rect 230532 218016 230538 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235810 218056 235816 218068
rect 235408 218028 235816 218056
rect 235408 218016 235414 218028
rect 235810 218016 235816 218028
rect 235868 218016 235874 218068
rect 240318 218016 240324 218068
rect 240376 218056 240382 218068
rect 241330 218056 241336 218068
rect 240376 218028 241336 218056
rect 240376 218016 240382 218028
rect 241330 218016 241336 218028
rect 241388 218016 241394 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244090 218056 244096 218068
rect 243688 218028 244096 218056
rect 243688 218016 243694 218028
rect 244090 218016 244096 218028
rect 244148 218016 244154 218068
rect 244458 218016 244464 218068
rect 244516 218056 244522 218068
rect 245286 218056 245292 218068
rect 244516 218028 245292 218056
rect 244516 218016 244522 218028
rect 245286 218016 245292 218028
rect 245344 218016 245350 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248322 218056 248328 218068
rect 247828 218028 248328 218056
rect 247828 218016 247834 218028
rect 248322 218016 248328 218028
rect 248380 218016 248386 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249242 218056 249248 218068
rect 248656 218028 249248 218056
rect 248656 218016 248662 218028
rect 249242 218016 249248 218028
rect 249300 218016 249306 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 250898 218056 250904 218068
rect 250312 218028 250904 218056
rect 250312 218016 250318 218028
rect 250898 218016 250904 218028
rect 250956 218016 250962 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 256050 218016 256056 218068
rect 256108 218056 256114 218068
rect 256510 218056 256516 218068
rect 256108 218028 256516 218056
rect 256108 218016 256114 218028
rect 256510 218016 256516 218028
rect 256568 218016 256574 218068
rect 256878 218016 256884 218068
rect 256936 218056 256942 218068
rect 257522 218056 257528 218068
rect 256936 218028 257528 218056
rect 256936 218016 256942 218028
rect 257522 218016 257528 218028
rect 257580 218016 257586 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259362 218056 259368 218068
rect 258592 218028 259368 218056
rect 258592 218016 258598 218028
rect 259362 218016 259368 218028
rect 259420 218016 259426 218068
rect 260190 218016 260196 218068
rect 260248 218056 260254 218068
rect 260742 218056 260748 218068
rect 260248 218028 260748 218056
rect 260248 218016 260254 218028
rect 260742 218016 260748 218028
rect 260800 218016 260806 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 268930 218056 268936 218068
rect 268528 218028 268936 218056
rect 268528 218016 268534 218028
rect 268930 218016 268936 218028
rect 268988 218016 268994 218068
rect 269298 218016 269304 218068
rect 269356 218056 269362 218068
rect 270218 218056 270224 218068
rect 269356 218028 270224 218056
rect 269356 218016 269362 218028
rect 270218 218016 270224 218028
rect 270276 218016 270282 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 272518 218056 272524 218068
rect 271012 218028 272524 218056
rect 271012 218016 271018 218028
rect 272518 218016 272524 218028
rect 272576 218016 272582 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278590 218056 278596 218068
rect 277636 218028 278596 218056
rect 277636 218016 277642 218028
rect 278590 218016 278596 218028
rect 278648 218016 278654 218068
rect 280890 218016 280896 218068
rect 280948 218056 280954 218068
rect 281442 218056 281448 218068
rect 280948 218028 281448 218056
rect 280948 218016 280954 218028
rect 281442 218016 281448 218028
rect 281500 218016 281506 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282730 218056 282736 218068
rect 281776 218028 282736 218056
rect 281776 218016 281782 218028
rect 282730 218016 282736 218028
rect 282788 218016 282794 218068
rect 283374 218016 283380 218068
rect 283432 218056 283438 218068
rect 284294 218056 284300 218068
rect 283432 218028 284300 218056
rect 283432 218016 283438 218028
rect 284294 218016 284300 218028
rect 284352 218016 284358 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288066 218056 288072 218068
rect 287572 218028 288072 218056
rect 287572 218016 287578 218028
rect 288066 218016 288072 218028
rect 288124 218016 288130 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289630 218056 289636 218068
rect 289228 218028 289636 218056
rect 289228 218016 289234 218028
rect 289630 218016 289636 218028
rect 289688 218016 289694 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 291102 218056 291108 218068
rect 290056 218028 291108 218056
rect 290056 218016 290062 218028
rect 291102 218016 291108 218028
rect 291160 218016 291166 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299382 218056 299388 218068
rect 298336 218028 299388 218056
rect 298336 218016 298342 218028
rect 299382 218016 299388 218028
rect 299440 218016 299446 218068
rect 299934 218016 299940 218068
rect 299992 218056 299998 218068
rect 300670 218056 300676 218068
rect 299992 218028 300676 218056
rect 299992 218016 299998 218028
rect 300670 218016 300676 218028
rect 300728 218016 300734 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306190 218056 306196 218068
rect 305788 218028 306196 218056
rect 305788 218016 305794 218028
rect 306190 218016 306196 218028
rect 306248 218016 306254 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 308214 218016 308220 218068
rect 308272 218056 308278 218068
rect 308858 218056 308864 218068
rect 308272 218028 308864 218056
rect 308272 218016 308278 218028
rect 308858 218016 308864 218028
rect 308916 218016 308922 218068
rect 309870 218016 309876 218068
rect 309928 218056 309934 218068
rect 310330 218056 310336 218068
rect 309928 218028 310336 218056
rect 309928 218016 309934 218028
rect 310330 218016 310336 218028
rect 310388 218016 310394 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 312906 218056 312912 218068
rect 312412 218028 312912 218056
rect 312412 218016 312418 218028
rect 312906 218016 312912 218028
rect 312964 218016 312970 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315482 218056 315488 218068
rect 314896 218028 315488 218056
rect 314896 218016 314902 218028
rect 315482 218016 315488 218028
rect 315540 218016 315546 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 317966 218056 317972 218068
rect 317380 218028 317972 218056
rect 317380 218016 317386 218028
rect 317966 218016 317972 218028
rect 318024 218016 318030 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 320082 218056 320088 218068
rect 319036 218028 320088 218056
rect 319036 218016 319042 218028
rect 320082 218016 320088 218028
rect 320140 218016 320146 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 323118 218016 323124 218068
rect 323176 218056 323182 218068
rect 323946 218056 323952 218068
rect 323176 218028 323952 218056
rect 323176 218016 323182 218028
rect 323946 218016 323952 218028
rect 324004 218016 324010 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325510 218056 325516 218068
rect 324832 218028 325516 218056
rect 324832 218016 324838 218028
rect 325510 218016 325516 218028
rect 325568 218016 325574 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 330570 218016 330576 218068
rect 330628 218056 330634 218068
rect 331030 218056 331036 218068
rect 330628 218028 331036 218056
rect 330628 218016 330634 218028
rect 331030 218016 331036 218028
rect 331088 218016 331094 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335170 218056 335176 218068
rect 334768 218028 335176 218056
rect 334768 218016 334774 218028
rect 335170 218016 335176 218028
rect 335228 218016 335234 218068
rect 337194 218016 337200 218068
rect 337252 218056 337258 218068
rect 337746 218056 337752 218068
rect 337252 218028 337752 218056
rect 337252 218016 337258 218028
rect 337746 218016 337752 218028
rect 337804 218016 337810 218068
rect 338850 218016 338856 218068
rect 338908 218056 338914 218068
rect 339402 218056 339408 218068
rect 338908 218028 339408 218056
rect 338908 218016 338914 218028
rect 339402 218016 339408 218028
rect 339460 218016 339466 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 345474 218016 345480 218068
rect 345532 218056 345538 218068
rect 347222 218056 347228 218068
rect 345532 218028 347228 218056
rect 345532 218016 345538 218028
rect 347222 218016 347228 218028
rect 347280 218016 347286 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 349614 218016 349620 218068
rect 349672 218056 349678 218068
rect 350166 218056 350172 218068
rect 349672 218028 350172 218056
rect 349672 218016 349678 218028
rect 350166 218016 350172 218028
rect 350224 218016 350230 218068
rect 352098 218016 352104 218068
rect 352156 218056 352162 218068
rect 353294 218056 353300 218068
rect 352156 218028 353300 218056
rect 352156 218016 352162 218028
rect 353294 218016 353300 218028
rect 353352 218016 353358 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 357250 218056 357256 218068
rect 356296 218028 357256 218056
rect 356296 218016 356302 218028
rect 357250 218016 357256 218028
rect 357308 218016 357314 218068
rect 357894 218016 357900 218068
rect 357952 218056 357958 218068
rect 358538 218056 358544 218068
rect 357952 218028 358544 218056
rect 357952 218016 357958 218028
rect 358538 218016 358544 218028
rect 358596 218016 358602 218068
rect 359550 218016 359556 218068
rect 359608 218056 359614 218068
rect 360102 218056 360108 218068
rect 359608 218028 360108 218056
rect 359608 218016 359614 218028
rect 360102 218016 360108 218028
rect 360160 218016 360166 218068
rect 360378 218016 360384 218068
rect 360436 218056 360442 218068
rect 361022 218056 361028 218068
rect 360436 218028 361028 218056
rect 360436 218016 360442 218028
rect 361022 218016 361028 218028
rect 361080 218016 361086 218068
rect 367830 218016 367836 218068
rect 367888 218056 367894 218068
rect 368382 218056 368388 218068
rect 367888 218028 368388 218056
rect 367888 218016 367894 218028
rect 368382 218016 368388 218028
rect 368440 218016 368446 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373534 218056 373540 218068
rect 372856 218028 373540 218056
rect 372856 218016 372862 218028
rect 373534 218016 373540 218028
rect 373592 218016 373598 218068
rect 374454 218016 374460 218068
rect 374512 218056 374518 218068
rect 375006 218056 375012 218068
rect 374512 218028 375012 218056
rect 374512 218016 374518 218028
rect 375006 218016 375012 218028
rect 375064 218016 375070 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376662 218056 376668 218068
rect 376168 218028 376668 218056
rect 376168 218016 376174 218028
rect 376662 218016 376668 218028
rect 376720 218016 376726 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379238 218056 379244 218068
rect 378652 218028 379244 218056
rect 378652 218016 378658 218028
rect 379238 218016 379244 218028
rect 379296 218016 379302 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 382090 218056 382096 218068
rect 381136 218028 382096 218056
rect 381136 218016 381142 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 385218 218016 385224 218068
rect 385276 218056 385282 218068
rect 386046 218056 386052 218068
rect 385276 218028 386052 218056
rect 385276 218016 385282 218028
rect 386046 218016 386052 218028
rect 386104 218016 386110 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390462 218056 390468 218068
rect 389416 218028 390468 218056
rect 389416 218016 389422 218028
rect 390462 218016 390468 218028
rect 390520 218016 390526 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393130 218056 393136 218068
rect 392728 218028 393136 218056
rect 392728 218016 392734 218028
rect 393130 218016 393136 218028
rect 393188 218016 393194 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394510 218056 394516 218068
rect 393556 218028 394516 218056
rect 393556 218016 393562 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395798 218056 395804 218068
rect 395212 218028 395804 218056
rect 395212 218016 395218 218028
rect 395798 218016 395804 218028
rect 395856 218016 395862 218068
rect 397638 218016 397644 218068
rect 397696 218056 397702 218068
rect 401318 218056 401324 218068
rect 397696 218028 401324 218056
rect 397696 218016 397702 218028
rect 401318 218016 401324 218028
rect 401376 218016 401382 218068
rect 401778 218016 401784 218068
rect 401836 218056 401842 218068
rect 402790 218056 402796 218068
rect 401836 218028 402796 218056
rect 401836 218016 401842 218028
rect 402790 218016 402796 218028
rect 402848 218016 402854 218068
rect 403434 218016 403440 218068
rect 403492 218056 403498 218068
rect 403986 218056 403992 218068
rect 403492 218028 403992 218056
rect 403492 218016 403498 218028
rect 403986 218016 403992 218028
rect 404044 218016 404050 218068
rect 405090 218016 405096 218068
rect 405148 218056 405154 218068
rect 405550 218056 405556 218068
rect 405148 218028 405556 218056
rect 405148 218016 405154 218028
rect 405550 218016 405556 218028
rect 405608 218016 405614 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 428458 218056 428464 218068
rect 427504 218028 428464 218056
rect 427504 218016 427510 218028
rect 428458 218016 428464 218028
rect 428516 218016 428522 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 435726 218016 435732 218068
rect 435784 218056 435790 218068
rect 436278 218056 436284 218068
rect 435784 218028 436284 218056
rect 435784 218016 435790 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436554 218016 436560 218068
rect 436612 218056 436618 218068
rect 437474 218056 437480 218068
rect 436612 218028 437480 218056
rect 436612 218016 436618 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438210 218016 438216 218068
rect 438268 218056 438274 218068
rect 438854 218056 438860 218068
rect 438268 218028 438860 218056
rect 438268 218016 438274 218028
rect 438854 218016 438860 218028
rect 438912 218016 438918 218068
rect 439866 218016 439872 218068
rect 439924 218056 439930 218068
rect 440326 218056 440332 218068
rect 439924 218028 440332 218056
rect 439924 218016 439930 218028
rect 440326 218016 440332 218028
rect 440384 218016 440390 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 455598 218016 455604 218068
rect 455656 218056 455662 218068
rect 457162 218056 457168 218068
rect 455656 218028 457168 218056
rect 455656 218016 455662 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 492030 218016 492036 218068
rect 492088 218056 492094 218068
rect 505646 218056 505652 218068
rect 492088 218028 505652 218056
rect 492088 218016 492094 218028
rect 505646 218016 505652 218028
rect 505704 218016 505710 218068
rect 507670 218016 507676 218068
rect 507728 218056 507734 218068
rect 563348 218056 563376 218096
rect 507728 218028 563376 218056
rect 572272 218056 572300 218096
rect 615678 218056 615684 218068
rect 572272 218028 615684 218056
rect 507728 218016 507734 218028
rect 615678 218016 615684 218028
rect 615736 218016 615742 218068
rect 646590 218016 646596 218068
rect 646648 218056 646654 218068
rect 653398 218056 653404 218068
rect 646648 218028 653404 218056
rect 646648 218016 646654 218028
rect 653398 218016 653404 218028
rect 653456 218016 653462 218068
rect 676214 218016 676220 218068
rect 676272 218056 676278 218068
rect 676858 218056 676864 218068
rect 676272 218028 676864 218056
rect 676272 218016 676278 218028
rect 676858 218016 676864 218028
rect 676916 218016 676922 218068
rect 563514 217948 563520 218000
rect 563572 217988 563578 218000
rect 572070 217988 572076 218000
rect 563572 217960 572076 217988
rect 563572 217948 563578 217960
rect 572070 217948 572076 217960
rect 572128 217948 572134 218000
rect 131022 217812 131028 217864
rect 131080 217852 131086 217864
rect 197722 217852 197728 217864
rect 131080 217824 197728 217852
rect 131080 217812 131086 217824
rect 197722 217812 197728 217824
rect 197780 217812 197786 217864
rect 523034 217812 523040 217864
rect 523092 217852 523098 217864
rect 524230 217852 524236 217864
rect 523092 217824 524236 217852
rect 523092 217812 523098 217824
rect 524230 217812 524236 217824
rect 524288 217812 524294 217864
rect 535454 217812 535460 217864
rect 535512 217852 535518 217864
rect 536650 217852 536656 217864
rect 535512 217824 536656 217852
rect 535512 217812 535518 217824
rect 536650 217812 536656 217824
rect 536708 217812 536714 217864
rect 536834 217812 536840 217864
rect 536892 217852 536898 217864
rect 536892 217824 598428 217852
rect 536892 217812 536898 217824
rect 116946 217676 116952 217728
rect 117004 217716 117010 217728
rect 189258 217716 189264 217728
rect 117004 217688 189264 217716
rect 117004 217676 117010 217688
rect 189258 217676 189264 217688
rect 189316 217676 189322 217728
rect 525978 217676 525984 217728
rect 526036 217716 526042 217728
rect 526530 217716 526536 217728
rect 526036 217688 526536 217716
rect 526036 217676 526042 217688
rect 526530 217676 526536 217688
rect 526588 217676 526594 217728
rect 535914 217676 535920 217728
rect 535972 217716 535978 217728
rect 598198 217716 598204 217728
rect 535972 217688 598204 217716
rect 535972 217676 535978 217688
rect 598198 217676 598204 217688
rect 598256 217676 598262 217728
rect 598400 217716 598428 217824
rect 598566 217812 598572 217864
rect 598624 217852 598630 217864
rect 598624 217824 603258 217852
rect 598624 217812 598630 217824
rect 598400 217688 600728 217716
rect 600700 217648 600728 217688
rect 601510 217676 601516 217728
rect 601568 217716 601574 217728
rect 602338 217716 602344 217728
rect 601568 217688 602344 217716
rect 601568 217676 601574 217688
rect 602338 217676 602344 217688
rect 602396 217676 602402 217728
rect 603230 217716 603258 217824
rect 603350 217812 603356 217864
rect 603408 217852 603414 217864
rect 613378 217852 613384 217864
rect 603408 217824 613384 217852
rect 603408 217812 603414 217824
rect 613378 217812 613384 217824
rect 613436 217812 613442 217864
rect 603994 217716 604000 217728
rect 603230 217688 604000 217716
rect 603994 217676 604000 217688
rect 604052 217676 604058 217728
rect 604454 217676 604460 217728
rect 604512 217716 604518 217728
rect 616874 217716 616880 217728
rect 604512 217688 616880 217716
rect 604512 217676 604518 217688
rect 616874 217676 616880 217688
rect 616932 217676 616938 217728
rect 600700 217620 601096 217648
rect 103698 217540 103704 217592
rect 103756 217580 103762 217592
rect 178402 217580 178408 217592
rect 103756 217552 178408 217580
rect 103756 217540 103762 217552
rect 178402 217540 178408 217552
rect 178460 217540 178466 217592
rect 530578 217540 530584 217592
rect 530636 217580 530642 217592
rect 530946 217580 530952 217592
rect 530636 217552 530952 217580
rect 530636 217540 530642 217552
rect 530946 217540 530952 217552
rect 531004 217580 531010 217592
rect 536834 217580 536840 217592
rect 531004 217552 536840 217580
rect 531004 217540 531010 217552
rect 536834 217540 536840 217552
rect 536892 217540 536898 217592
rect 538214 217540 538220 217592
rect 538272 217580 538278 217592
rect 539134 217580 539140 217592
rect 538272 217552 539140 217580
rect 538272 217540 538278 217552
rect 539134 217540 539140 217552
rect 539192 217540 539198 217592
rect 545758 217540 545764 217592
rect 545816 217580 545822 217592
rect 600130 217580 600136 217592
rect 545816 217552 600136 217580
rect 545816 217540 545822 217552
rect 600130 217540 600136 217552
rect 600188 217540 600194 217592
rect 601068 217580 601096 217620
rect 603442 217580 603448 217592
rect 601068 217552 603448 217580
rect 603442 217540 603448 217552
rect 603500 217540 603506 217592
rect 675846 217540 675852 217592
rect 675904 217580 675910 217592
rect 676674 217580 676680 217592
rect 675904 217552 676680 217580
rect 675904 217540 675910 217552
rect 676674 217540 676680 217552
rect 676732 217540 676738 217592
rect 93762 217404 93768 217456
rect 93820 217444 93826 217456
rect 171226 217444 171232 217456
rect 93820 217416 171232 217444
rect 93820 217404 93826 217416
rect 171226 217404 171232 217416
rect 171284 217404 171290 217456
rect 526530 217404 526536 217456
rect 526588 217444 526594 217456
rect 601510 217444 601516 217456
rect 526588 217416 601516 217444
rect 526588 217404 526594 217416
rect 601510 217404 601516 217416
rect 601568 217404 601574 217456
rect 601878 217404 601884 217456
rect 601936 217444 601942 217456
rect 628282 217444 628288 217456
rect 601936 217416 628288 217444
rect 601936 217404 601942 217416
rect 628282 217404 628288 217416
rect 628340 217404 628346 217456
rect 170306 217308 170312 217320
rect 93826 217280 170312 217308
rect 92060 217200 92066 217252
rect 92118 217240 92124 217252
rect 93826 217240 93854 217280
rect 170306 217268 170312 217280
rect 170364 217268 170370 217320
rect 533430 217268 533436 217320
rect 533488 217308 533494 217320
rect 598566 217308 598572 217320
rect 533488 217280 598572 217308
rect 533488 217268 533494 217280
rect 598566 217268 598572 217280
rect 598624 217268 598630 217320
rect 598750 217268 598756 217320
rect 598808 217308 598814 217320
rect 598808 217280 599348 217308
rect 598808 217268 598814 217280
rect 92118 217212 93854 217240
rect 92118 217200 92124 217212
rect 436094 217200 436100 217252
rect 436152 217240 436158 217252
rect 437336 217240 437342 217252
rect 436152 217212 437342 217240
rect 436152 217200 436158 217212
rect 437336 217200 437342 217212
rect 437394 217200 437400 217252
rect 448514 217200 448520 217252
rect 448572 217240 448578 217252
rect 449756 217240 449762 217252
rect 448572 217212 449762 217240
rect 448572 217200 448578 217212
rect 449756 217200 449762 217212
rect 449814 217200 449820 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 489914 217200 489920 217252
rect 489972 217240 489978 217252
rect 491156 217240 491162 217252
rect 489972 217212 491162 217240
rect 489972 217200 489978 217212
rect 491156 217200 491162 217212
rect 491214 217200 491220 217252
rect 498194 217200 498200 217252
rect 498252 217240 498258 217252
rect 499436 217240 499442 217252
rect 498252 217212 499442 217240
rect 498252 217200 498258 217212
rect 499436 217200 499442 217212
rect 499494 217200 499500 217252
rect 511028 217132 511034 217184
rect 511086 217172 511092 217184
rect 562134 217172 562140 217184
rect 511086 217144 562140 217172
rect 511086 217132 511092 217144
rect 562134 217132 562140 217144
rect 562192 217132 562198 217184
rect 562502 217172 562508 217184
rect 562382 217144 562508 217172
rect 503162 217064 503168 217116
rect 503220 217104 503226 217116
rect 503576 217104 503582 217116
rect 503220 217076 503582 217104
rect 503220 217064 503226 217076
rect 503576 217064 503582 217076
rect 503634 217104 503640 217116
rect 503634 217076 505094 217104
rect 503634 217064 503640 217076
rect 505066 217036 505094 217076
rect 562382 217036 562410 217144
rect 562502 217132 562508 217144
rect 562560 217132 562566 217184
rect 562686 217132 562692 217184
rect 562744 217132 562750 217184
rect 563054 217132 563060 217184
rect 563112 217172 563118 217184
rect 599118 217172 599124 217184
rect 563112 217144 599124 217172
rect 563112 217132 563118 217144
rect 599118 217132 599124 217144
rect 599176 217132 599182 217184
rect 599320 217172 599348 217280
rect 600130 217268 600136 217320
rect 600188 217308 600194 217320
rect 606754 217308 606760 217320
rect 600188 217280 606760 217308
rect 600188 217268 600194 217280
rect 606754 217268 606760 217280
rect 606812 217268 606818 217320
rect 642174 217268 642180 217320
rect 642232 217308 642238 217320
rect 658918 217308 658924 217320
rect 642232 217280 658924 217308
rect 642232 217268 642238 217280
rect 658918 217268 658924 217280
rect 658976 217268 658982 217320
rect 601326 217172 601332 217184
rect 599320 217144 601332 217172
rect 601326 217132 601332 217144
rect 601384 217132 601390 217184
rect 601510 217132 601516 217184
rect 601568 217172 601574 217184
rect 604546 217172 604552 217184
rect 601568 217144 604552 217172
rect 601568 217132 601574 217144
rect 604546 217132 604552 217144
rect 604604 217132 604610 217184
rect 505066 217008 562410 217036
rect 562704 217036 562732 217132
rect 608962 217036 608968 217048
rect 562704 217008 608968 217036
rect 608962 216996 608968 217008
rect 609020 216996 609026 217048
rect 609882 216996 609888 217048
rect 609940 217036 609946 217048
rect 614114 217036 614120 217048
rect 609940 217008 614120 217036
rect 609940 216996 609946 217008
rect 614114 216996 614120 217008
rect 614172 216996 614178 217048
rect 574094 216860 574100 216912
rect 574152 216900 574158 216912
rect 597554 216900 597560 216912
rect 574152 216872 597560 216900
rect 574152 216860 574158 216872
rect 597554 216860 597560 216872
rect 597612 216860 597618 216912
rect 598198 216860 598204 216912
rect 598256 216900 598262 216912
rect 600774 216900 600780 216912
rect 598256 216872 600780 216900
rect 598256 216860 598262 216872
rect 600774 216860 600780 216872
rect 600832 216860 600838 216912
rect 612274 216900 612280 216912
rect 600976 216872 612280 216900
rect 594794 216724 594800 216776
rect 594852 216764 594858 216776
rect 600976 216764 601004 216872
rect 612274 216860 612280 216872
rect 612332 216860 612338 216912
rect 594852 216736 601004 216764
rect 594852 216724 594858 216736
rect 601326 216724 601332 216776
rect 601384 216764 601390 216776
rect 623866 216764 623872 216776
rect 601384 216736 623872 216764
rect 601384 216724 601390 216736
rect 623866 216724 623872 216736
rect 623924 216724 623930 216776
rect 648246 216588 648252 216640
rect 648304 216628 648310 216640
rect 656158 216628 656164 216640
rect 648304 216600 656164 216628
rect 648304 216588 648310 216600
rect 656158 216588 656164 216600
rect 656216 216588 656222 216640
rect 675938 215500 675944 215552
rect 675996 215540 676002 215552
rect 677042 215540 677048 215552
rect 675996 215512 677048 215540
rect 675996 215500 676002 215512
rect 677042 215500 677048 215512
rect 677100 215500 677106 215552
rect 575474 214820 575480 214872
rect 575532 214860 575538 214872
rect 622394 214860 622400 214872
rect 575532 214832 622400 214860
rect 575532 214820 575538 214832
rect 622394 214820 622400 214832
rect 622452 214820 622458 214872
rect 649718 214820 649724 214872
rect 649776 214860 649782 214872
rect 657722 214860 657728 214872
rect 649776 214832 657728 214860
rect 649776 214820 649782 214832
rect 657722 214820 657728 214832
rect 657780 214820 657786 214872
rect 574278 214684 574284 214736
rect 574336 214724 574342 214736
rect 616690 214724 616696 214736
rect 574336 214696 616696 214724
rect 574336 214684 574342 214696
rect 616690 214684 616696 214696
rect 616748 214684 616754 214736
rect 617058 214684 617064 214736
rect 617116 214724 617122 214736
rect 617794 214724 617800 214736
rect 617116 214696 617800 214724
rect 617116 214684 617122 214696
rect 617794 214684 617800 214696
rect 617852 214684 617858 214736
rect 621014 214684 621020 214736
rect 621072 214724 621078 214736
rect 621658 214724 621664 214736
rect 621072 214696 621664 214724
rect 621072 214684 621078 214696
rect 621658 214684 621664 214696
rect 621716 214684 621722 214736
rect 630030 214684 630036 214736
rect 630088 214724 630094 214736
rect 632882 214724 632888 214736
rect 630088 214696 632888 214724
rect 630088 214684 630094 214696
rect 632882 214684 632888 214696
rect 632940 214684 632946 214736
rect 644566 214684 644572 214736
rect 644624 214724 644630 214736
rect 654778 214724 654784 214736
rect 644624 214696 654784 214724
rect 644624 214684 644630 214696
rect 654778 214684 654784 214696
rect 654836 214684 654842 214736
rect 574462 214548 574468 214600
rect 574520 214588 574526 214600
rect 625522 214588 625528 214600
rect 574520 214560 625528 214588
rect 574520 214548 574526 214560
rect 625522 214548 625528 214560
rect 625580 214548 625586 214600
rect 654870 214548 654876 214600
rect 654928 214588 654934 214600
rect 664438 214588 664444 214600
rect 654928 214560 664444 214588
rect 654928 214548 654934 214560
rect 664438 214548 664444 214560
rect 664496 214548 664502 214600
rect 664806 214548 664812 214600
rect 664864 214588 664870 214600
rect 665818 214588 665824 214600
rect 664864 214560 665824 214588
rect 664864 214548 664870 214560
rect 665818 214548 665824 214560
rect 665876 214548 665882 214600
rect 610066 214412 610072 214464
rect 610124 214452 610130 214464
rect 610618 214452 610624 214464
rect 610124 214424 610624 214452
rect 610124 214412 610130 214424
rect 610618 214412 610624 214424
rect 610676 214412 610682 214464
rect 616690 214412 616696 214464
rect 616748 214452 616754 214464
rect 624418 214452 624424 214464
rect 616748 214424 624424 214452
rect 616748 214412 616754 214424
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 626350 214276 626356 214328
rect 626408 214316 626414 214328
rect 628834 214316 628840 214328
rect 626408 214288 628840 214316
rect 626408 214276 626414 214288
rect 628834 214276 628840 214288
rect 628892 214276 628898 214328
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 41690 213976 41696 213988
rect 35860 213948 41696 213976
rect 35860 213936 35866 213948
rect 41690 213936 41696 213948
rect 41748 213936 41754 213988
rect 627454 213936 627460 213988
rect 627512 213976 627518 213988
rect 629386 213976 629392 213988
rect 627512 213948 629392 213976
rect 627512 213936 627518 213948
rect 629386 213936 629392 213948
rect 629444 213936 629450 213988
rect 663150 213868 663156 213920
rect 663208 213908 663214 213920
rect 663702 213908 663708 213920
rect 663208 213880 663708 213908
rect 663208 213868 663214 213880
rect 663702 213868 663708 213880
rect 663760 213868 663766 213920
rect 659562 213596 659568 213648
rect 659620 213636 659626 213648
rect 665542 213636 665548 213648
rect 659620 213608 665548 213636
rect 659620 213596 659626 213608
rect 665542 213596 665548 213608
rect 665600 213596 665606 213648
rect 574094 213460 574100 213512
rect 574152 213500 574158 213512
rect 594794 213500 594800 213512
rect 574152 213472 594800 213500
rect 574152 213460 574158 213472
rect 594794 213460 594800 213472
rect 594852 213460 594858 213512
rect 647142 213460 647148 213512
rect 647200 213500 647206 213512
rect 649902 213500 649908 213512
rect 647200 213472 649908 213500
rect 647200 213460 647206 213472
rect 649902 213460 649908 213472
rect 649960 213460 649966 213512
rect 574646 213324 574652 213376
rect 574704 213364 574710 213376
rect 612826 213364 612832 213376
rect 574704 213336 612832 213364
rect 574704 213324 574710 213336
rect 612826 213324 612832 213336
rect 612884 213324 612890 213376
rect 651098 213324 651104 213376
rect 651156 213364 651162 213376
rect 657538 213364 657544 213376
rect 651156 213336 657544 213364
rect 651156 213324 651162 213336
rect 657538 213324 657544 213336
rect 657596 213324 657602 213376
rect 574830 213188 574836 213240
rect 574888 213228 574894 213240
rect 616138 213228 616144 213240
rect 574888 213200 616144 213228
rect 574888 213188 574894 213200
rect 616138 213188 616144 213200
rect 616196 213188 616202 213240
rect 643830 213188 643836 213240
rect 643888 213228 643894 213240
rect 650638 213228 650644 213240
rect 643888 213200 650644 213228
rect 643888 213188 643894 213200
rect 650638 213188 650644 213200
rect 650696 213188 650702 213240
rect 658182 212848 658188 212900
rect 658240 212888 658246 212900
rect 659102 212888 659108 212900
rect 658240 212860 659108 212888
rect 658240 212848 658246 212860
rect 659102 212848 659108 212860
rect 659160 212848 659166 212900
rect 650454 212712 650460 212764
rect 650512 212752 650518 212764
rect 651282 212752 651288 212764
rect 650512 212724 651288 212752
rect 650512 212712 650518 212724
rect 651282 212712 651288 212724
rect 651340 212712 651346 212764
rect 664254 212712 664260 212764
rect 664312 212752 664318 212764
rect 665082 212752 665088 212764
rect 664312 212724 665088 212752
rect 664312 212712 664318 212724
rect 665082 212712 665088 212724
rect 665140 212712 665146 212764
rect 632698 212508 632704 212560
rect 632756 212548 632762 212560
rect 634354 212548 634360 212560
rect 632756 212520 634360 212548
rect 632756 212508 632762 212520
rect 634354 212508 634360 212520
rect 634412 212508 634418 212560
rect 630674 212372 630680 212424
rect 630732 212412 630738 212424
rect 631594 212412 631600 212424
rect 630732 212384 631600 212412
rect 630732 212372 630738 212384
rect 631594 212372 631600 212384
rect 631652 212372 631658 212424
rect 35802 211556 35808 211608
rect 35860 211596 35866 211608
rect 39574 211596 39580 211608
rect 35860 211568 39580 211596
rect 35860 211556 35866 211568
rect 39574 211556 39580 211568
rect 39632 211556 39638 211608
rect 35618 211284 35624 211336
rect 35676 211324 35682 211336
rect 41690 211324 41696 211336
rect 35676 211296 41696 211324
rect 35676 211284 35682 211296
rect 41690 211284 41696 211296
rect 41748 211284 41754 211336
rect 35434 211148 35440 211200
rect 35492 211188 35498 211200
rect 41322 211188 41328 211200
rect 35492 211160 41328 211188
rect 35492 211148 35498 211160
rect 41322 211148 41328 211160
rect 41380 211148 41386 211200
rect 578510 211148 578516 211200
rect 578568 211188 578574 211200
rect 580902 211188 580908 211200
rect 578568 211160 580908 211188
rect 578568 211148 578574 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 680354 211148 680360 211200
rect 680412 211188 680418 211200
rect 683114 211188 683120 211200
rect 680412 211160 683120 211188
rect 680412 211148 680418 211160
rect 683114 211148 683120 211160
rect 683172 211148 683178 211200
rect 633434 211012 633440 211064
rect 633492 211052 633498 211064
rect 633802 211052 633808 211064
rect 633492 211024 633808 211052
rect 633492 211012 633498 211024
rect 633802 211012 633808 211024
rect 633860 211012 633866 211064
rect 635550 210128 635556 210180
rect 635608 210168 635614 210180
rect 636562 210168 636568 210180
rect 635608 210140 636568 210168
rect 635608 210128 635614 210140
rect 636562 210128 636568 210140
rect 636620 210128 636626 210180
rect 35802 209788 35808 209840
rect 35860 209828 35866 209840
rect 40218 209828 40224 209840
rect 35860 209800 40224 209828
rect 35860 209788 35866 209800
rect 40218 209788 40224 209800
rect 40276 209788 40282 209840
rect 579522 209788 579528 209840
rect 579580 209828 579586 209840
rect 582282 209828 582288 209840
rect 579580 209800 582288 209828
rect 579580 209788 579586 209800
rect 582282 209788 582288 209800
rect 582340 209788 582346 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 581638 208564 581644 208616
rect 581696 208604 581702 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652018 209516 652024 209568
rect 652076 209556 652082 209568
rect 652076 209528 654134 209556
rect 652076 209516 652082 209528
rect 654106 209080 654134 209528
rect 667566 209080 667572 209092
rect 654106 209052 667572 209080
rect 667566 209040 667572 209052
rect 667624 209040 667630 209092
rect 581696 208576 625154 208604
rect 581696 208564 581702 208576
rect 35802 208496 35808 208548
rect 35860 208536 35866 208548
rect 40494 208536 40500 208548
rect 35860 208508 40500 208536
rect 35860 208496 35866 208508
rect 40494 208496 40500 208508
rect 40552 208496 40558 208548
rect 35618 208360 35624 208412
rect 35676 208400 35682 208412
rect 40034 208400 40040 208412
rect 35676 208372 40040 208400
rect 35676 208360 35682 208372
rect 40034 208360 40040 208372
rect 40092 208360 40098 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 35802 207136 35808 207188
rect 35860 207176 35866 207188
rect 40770 207176 40776 207188
rect 35860 207148 40776 207176
rect 35860 207136 35866 207148
rect 40770 207136 40776 207148
rect 40828 207136 40834 207188
rect 580902 206864 580908 206916
rect 580960 206904 580966 206916
rect 589458 206904 589464 206916
rect 580960 206876 589464 206904
rect 580960 206864 580966 206876
rect 589458 206864 589464 206876
rect 589516 206864 589522 206916
rect 35802 205776 35808 205828
rect 35860 205816 35866 205828
rect 40954 205816 40960 205828
rect 35860 205788 40960 205816
rect 35860 205776 35866 205788
rect 40954 205776 40960 205788
rect 41012 205776 41018 205828
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 582282 205504 582288 205556
rect 582340 205544 582346 205556
rect 589458 205544 589464 205556
rect 582340 205516 589464 205544
rect 582340 205504 582346 205516
rect 589458 205504 589464 205516
rect 589516 205504 589522 205556
rect 35802 204552 35808 204604
rect 35860 204592 35866 204604
rect 40402 204592 40408 204604
rect 35860 204564 40408 204592
rect 35860 204552 35866 204564
rect 40402 204552 40408 204564
rect 40460 204552 40466 204604
rect 41690 204388 41696 204400
rect 36004 204360 41696 204388
rect 35618 204280 35624 204332
rect 35676 204320 35682 204332
rect 36004 204320 36032 204360
rect 41690 204348 41696 204360
rect 41748 204348 41754 204400
rect 42058 204348 42064 204400
rect 42116 204388 42122 204400
rect 43346 204388 43352 204400
rect 42116 204360 43352 204388
rect 42116 204348 42122 204360
rect 43346 204348 43352 204360
rect 43404 204348 43410 204400
rect 35676 204292 36032 204320
rect 35676 204280 35682 204292
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 42426 190136 42432 190188
rect 42484 190176 42490 190188
rect 42978 190176 42984 190188
rect 42484 190148 42984 190176
rect 42484 190136 42490 190148
rect 42978 190136 42984 190148
rect 43036 190136 43042 190188
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 42426 187620 42432 187672
rect 42484 187660 42490 187672
rect 43162 187660 43168 187672
rect 42484 187632 43168 187660
rect 42484 187620 42490 187632
rect 43162 187620 43168 187632
rect 43220 187620 43226 187672
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 582374 168376 582380 168428
rect 582432 168416 582438 168428
rect 589458 168416 589464 168428
rect 582432 168388 589464 168416
rect 582432 168376 582438 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579982 167016 579988 167068
rect 580040 167056 580046 167068
rect 589458 167056 589464 167068
rect 580040 167028 589464 167056
rect 580040 167016 580046 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589642 166308 589648 166320
rect 579580 166280 589648 166308
rect 579580 166268 579586 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 579338 165180 579344 165232
rect 579396 165220 579402 165232
rect 582374 165220 582380 165232
rect 579396 165192 582380 165220
rect 579396 165180 579402 165192
rect 582374 165180 582380 165192
rect 582432 165180 582438 165232
rect 668210 165180 668216 165232
rect 668268 165220 668274 165232
rect 669590 165220 669596 165232
rect 668268 165192 669596 165220
rect 668268 165180 668274 165192
rect 669590 165180 669596 165192
rect 669648 165180 669654 165232
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 578234 163616 578240 163668
rect 578292 163656 578298 163668
rect 579982 163656 579988 163668
rect 578292 163628 579988 163656
rect 578292 163616 578298 163628
rect 579982 163616 579988 163628
rect 580040 163616 580046 163668
rect 668210 163276 668216 163328
rect 668268 163316 668274 163328
rect 669774 163316 669780 163328
rect 668268 163288 669780 163316
rect 668268 163276 668274 163288
rect 669774 163276 669780 163288
rect 669832 163276 669838 163328
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 675846 162800 675852 162852
rect 675904 162840 675910 162852
rect 678238 162840 678244 162852
rect 675904 162812 678244 162840
rect 675904 162800 675910 162812
rect 678238 162800 678244 162812
rect 678296 162800 678302 162852
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 668210 160012 668216 160064
rect 668268 160052 668274 160064
rect 670326 160052 670332 160064
rect 668268 160024 670332 160052
rect 668268 160012 668274 160024
rect 670326 160012 670332 160024
rect 670384 160012 670390 160064
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 158720 585784 158772
rect 585836 158760 585842 158772
rect 589458 158760 589464 158772
rect 585836 158732 589464 158760
rect 585836 158720 585842 158732
rect 589458 158720 589464 158732
rect 589516 158720 589522 158772
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 668302 155116 668308 155168
rect 668360 155156 668366 155168
rect 670786 155156 670792 155168
rect 668360 155128 670792 155156
rect 668360 155116 668366 155128
rect 670786 155116 670792 155128
rect 670844 155116 670850 155168
rect 578326 154640 578332 154692
rect 578384 154680 578390 154692
rect 580534 154680 580540 154692
rect 578384 154652 580540 154680
rect 578384 154640 578390 154652
rect 580534 154640 580540 154652
rect 580592 154640 580598 154692
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580258 151784 580264 151836
rect 580316 151824 580322 151836
rect 589458 151824 589464 151836
rect 580316 151796 589464 151824
rect 580316 151784 580322 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 585778 150600 585784 150612
rect 578936 150572 585784 150600
rect 578936 150560 578942 150572
rect 585778 150560 585784 150572
rect 585836 150560 585842 150612
rect 585134 149064 585140 149116
rect 585192 149104 585198 149116
rect 589458 149104 589464 149116
rect 585192 149076 589464 149104
rect 585192 149064 585198 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 668210 148724 668216 148776
rect 668268 148764 668274 148776
rect 670142 148764 670148 148776
rect 668268 148736 670148 148764
rect 668268 148724 668274 148736
rect 670142 148724 670148 148736
rect 670200 148724 670206 148776
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 578878 146276 578884 146328
rect 578936 146316 578942 146328
rect 585134 146316 585140 146328
rect 578936 146288 585140 146316
rect 578936 146276 578942 146288
rect 585134 146276 585140 146288
rect 585192 146276 585198 146328
rect 584766 144916 584772 144968
rect 584824 144956 584830 144968
rect 589458 144956 589464 144968
rect 584824 144928 589464 144956
rect 584824 144916 584830 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 585778 143556 585784 143608
rect 585836 143596 585842 143608
rect 589458 143596 589464 143608
rect 585836 143568 589464 143596
rect 585836 143556 585842 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 580442 140768 580448 140820
rect 580500 140808 580506 140820
rect 589458 140808 589464 140820
rect 580500 140780 589464 140808
rect 580500 140768 580506 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580258 140740 580264 140752
rect 578660 140712 580264 140740
rect 578660 140700 578666 140712
rect 580258 140700 580264 140712
rect 580316 140700 580322 140752
rect 583018 139408 583024 139460
rect 583076 139448 583082 139460
rect 589458 139448 589464 139460
rect 583076 139420 589464 139448
rect 583076 139408 583082 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579522 138660 579528 138712
rect 579580 138700 579586 138712
rect 588538 138700 588544 138712
rect 579580 138672 588544 138700
rect 579580 138660 579586 138672
rect 588538 138660 588544 138672
rect 588596 138660 588602 138712
rect 579062 137300 579068 137352
rect 579120 137340 579126 137352
rect 584766 137340 584772 137352
rect 579120 137312 584772 137340
rect 579120 137300 579126 137312
rect 584766 137300 584772 137312
rect 584824 137300 584830 137352
rect 584582 136620 584588 136672
rect 584640 136660 584646 136672
rect 589458 136660 589464 136672
rect 584640 136632 589464 136660
rect 584640 136620 584646 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 668210 136212 668216 136264
rect 668268 136252 668274 136264
rect 669958 136252 669964 136264
rect 668268 136224 669964 136252
rect 668268 136212 668274 136224
rect 669958 136212 669964 136224
rect 670016 136212 670022 136264
rect 580258 134512 580264 134564
rect 580316 134552 580322 134564
rect 589458 134552 589464 134564
rect 580316 134524 589464 134552
rect 580316 134512 580322 134524
rect 589458 134512 589464 134524
rect 589516 134512 589522 134564
rect 585962 132472 585968 132524
rect 586020 132512 586026 132524
rect 589458 132512 589464 132524
rect 586020 132484 589464 132512
rect 586020 132472 586026 132484
rect 589458 132472 589464 132484
rect 589516 132472 589522 132524
rect 581822 131248 581828 131300
rect 581880 131288 581886 131300
rect 589458 131288 589464 131300
rect 581880 131260 589464 131288
rect 581880 131248 581886 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 578878 131112 578884 131164
rect 578936 131152 578942 131164
rect 585778 131152 585784 131164
rect 578936 131124 585784 131152
rect 578936 131112 578942 131124
rect 585778 131112 585784 131124
rect 585836 131112 585842 131164
rect 668578 129684 668584 129736
rect 668636 129724 668642 129736
rect 670786 129724 670792 129736
rect 668636 129696 670792 129724
rect 668636 129684 668642 129696
rect 670786 129684 670792 129696
rect 670844 129684 670850 129736
rect 583386 129140 583392 129192
rect 583444 129180 583450 129192
rect 590378 129180 590384 129192
rect 583444 129152 590384 129180
rect 583444 129140 583450 129152
rect 590378 129140 590384 129152
rect 590436 129140 590442 129192
rect 579522 129004 579528 129056
rect 579580 129044 579586 129056
rect 587158 129044 587164 129056
rect 579580 129016 587164 129044
rect 579580 129004 579586 129016
rect 587158 129004 587164 129016
rect 587216 129004 587222 129056
rect 587802 126964 587808 127016
rect 587860 127004 587866 127016
rect 589458 127004 589464 127016
rect 587860 126976 589464 127004
rect 587860 126964 587866 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 578326 125604 578332 125656
rect 578384 125644 578390 125656
rect 580442 125644 580448 125656
rect 578384 125616 580448 125644
rect 578384 125604 578390 125616
rect 580442 125604 580448 125616
rect 580500 125604 580506 125656
rect 675938 125264 675944 125316
rect 675996 125304 676002 125316
rect 676582 125304 676588 125316
rect 675996 125276 676588 125304
rect 675996 125264 676002 125276
rect 676582 125264 676588 125276
rect 676640 125264 676646 125316
rect 579062 124856 579068 124908
rect 579120 124896 579126 124908
rect 587802 124896 587808 124908
rect 579120 124868 587808 124896
rect 579120 124856 579126 124868
rect 587802 124856 587808 124868
rect 587860 124856 587866 124908
rect 578694 124108 578700 124160
rect 578752 124148 578758 124160
rect 583018 124148 583024 124160
rect 578752 124120 583024 124148
rect 578752 124108 578758 124120
rect 583018 124108 583024 124120
rect 583076 124108 583082 124160
rect 675846 123360 675852 123412
rect 675904 123400 675910 123412
rect 676398 123400 676404 123412
rect 675904 123372 676404 123400
rect 675904 123360 675910 123372
rect 676398 123360 676404 123372
rect 676456 123360 676462 123412
rect 584398 122816 584404 122868
rect 584456 122856 584462 122868
rect 589458 122856 589464 122868
rect 584456 122828 589464 122856
rect 584456 122816 584462 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 578878 122136 578884 122188
rect 578936 122176 578942 122188
rect 584582 122176 584588 122188
rect 578936 122148 584588 122176
rect 578936 122136 578942 122148
rect 584582 122136 584588 122148
rect 584640 122136 584646 122188
rect 580626 122000 580632 122052
rect 580684 122040 580690 122052
rect 590102 122040 590108 122052
rect 580684 122012 590108 122040
rect 580684 122000 580690 122012
rect 590102 122000 590108 122012
rect 590160 122000 590166 122052
rect 587342 121456 587348 121508
rect 587400 121496 587406 121508
rect 589274 121496 589280 121508
rect 587400 121468 589280 121496
rect 587400 121456 587406 121468
rect 589274 121456 589280 121468
rect 589332 121456 589338 121508
rect 583202 120708 583208 120760
rect 583260 120748 583266 120760
rect 590562 120748 590568 120760
rect 583260 120720 590568 120748
rect 583260 120708 583266 120720
rect 590562 120708 590568 120720
rect 590620 120708 590626 120760
rect 578510 118532 578516 118584
rect 578568 118572 578574 118584
rect 580258 118572 580264 118584
rect 578568 118544 580264 118572
rect 578568 118532 578574 118544
rect 580258 118532 580264 118544
rect 580316 118532 580322 118584
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 583386 116940 583392 116952
rect 579580 116912 583392 116940
rect 579580 116900 579586 116912
rect 583386 116900 583392 116912
rect 583444 116900 583450 116952
rect 675846 116492 675852 116544
rect 675904 116532 675910 116544
rect 676858 116532 676864 116544
rect 675904 116504 676864 116532
rect 675904 116492 675910 116504
rect 676858 116492 676864 116504
rect 676916 116492 676922 116544
rect 585778 115948 585784 116000
rect 585836 115988 585842 116000
rect 589458 115988 589464 116000
rect 585836 115960 589464 115988
rect 585836 115948 585842 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 584582 115200 584588 115252
rect 584640 115240 584646 115252
rect 589642 115240 589648 115252
rect 584640 115212 589648 115240
rect 584640 115200 584646 115212
rect 589642 115200 589648 115212
rect 589700 115200 589706 115252
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 583018 113160 583024 113212
rect 583076 113200 583082 113212
rect 589458 113200 589464 113212
rect 583076 113172 589464 113200
rect 583076 113160 583082 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579522 112820 579528 112872
rect 579580 112860 579586 112872
rect 585962 112860 585968 112872
rect 579580 112832 585968 112860
rect 579580 112820 579586 112832
rect 585962 112820 585968 112832
rect 586020 112820 586026 112872
rect 586146 112412 586152 112464
rect 586204 112452 586210 112464
rect 590102 112452 590108 112464
rect 586204 112424 590108 112452
rect 586204 112412 586210 112424
rect 590102 112412 590108 112424
rect 590160 112412 590166 112464
rect 668210 111460 668216 111512
rect 668268 111500 668274 111512
rect 670694 111500 670700 111512
rect 668268 111472 670700 111500
rect 668268 111460 668274 111472
rect 670694 111460 670700 111472
rect 670752 111460 670758 111512
rect 581638 110440 581644 110492
rect 581696 110480 581702 110492
rect 589458 110480 589464 110492
rect 581696 110452 589464 110480
rect 581696 110440 581702 110452
rect 589458 110440 589464 110452
rect 589516 110440 589522 110492
rect 579338 110236 579344 110288
rect 579396 110276 579402 110288
rect 581822 110276 581828 110288
rect 579396 110248 581828 110276
rect 579396 110236 579402 110248
rect 581822 110236 581828 110248
rect 581880 110236 581886 110288
rect 580442 109080 580448 109132
rect 580500 109120 580506 109132
rect 589458 109120 589464 109132
rect 580500 109092 589464 109120
rect 580500 109080 580506 109092
rect 589458 109080 589464 109092
rect 589516 109080 589522 109132
rect 578326 108944 578332 108996
rect 578384 108984 578390 108996
rect 580626 108984 580632 108996
rect 578384 108956 580632 108984
rect 578384 108944 578390 108956
rect 580626 108944 580632 108956
rect 580684 108944 580690 108996
rect 667934 108808 667940 108860
rect 667992 108848 667998 108860
rect 669958 108848 669964 108860
rect 667992 108820 669964 108848
rect 667992 108808 667998 108820
rect 669958 108808 669964 108820
rect 670016 108808 670022 108860
rect 582282 107652 582288 107704
rect 582340 107692 582346 107704
rect 589458 107692 589464 107704
rect 582340 107664 589464 107692
rect 582340 107652 582346 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 580258 106292 580264 106344
rect 580316 106332 580322 106344
rect 589458 106332 589464 106344
rect 580316 106304 589464 106332
rect 580316 106292 580322 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 579338 105612 579344 105664
rect 579396 105652 579402 105664
rect 582282 105652 582288 105664
rect 579396 105624 582288 105652
rect 579396 105612 579402 105624
rect 582282 105612 582288 105624
rect 582340 105612 582346 105664
rect 587158 104864 587164 104916
rect 587216 104904 587222 104916
rect 589826 104904 589832 104916
rect 587216 104876 589832 104904
rect 587216 104864 587222 104876
rect 589826 104864 589832 104876
rect 589884 104864 589890 104916
rect 578510 103368 578516 103420
rect 578568 103408 578574 103420
rect 588722 103408 588728 103420
rect 578568 103380 588728 103408
rect 578568 103368 578574 103380
rect 588722 103368 588728 103380
rect 588780 103368 588786 103420
rect 579154 102076 579160 102128
rect 579212 102116 579218 102128
rect 584398 102116 584404 102128
rect 579212 102088 584404 102116
rect 579212 102076 579218 102088
rect 584398 102076 584404 102088
rect 584456 102076 584462 102128
rect 584398 100104 584404 100156
rect 584456 100144 584462 100156
rect 589458 100144 589464 100156
rect 584456 100116 589464 100144
rect 584456 100104 584462 100116
rect 589458 100104 589464 100116
rect 589516 100104 589522 100156
rect 578602 99968 578608 100020
rect 578660 100008 578666 100020
rect 587342 100008 587348 100020
rect 578660 99980 587348 100008
rect 578660 99968 578666 99980
rect 587342 99968 587348 99980
rect 587400 99968 587406 100020
rect 592678 99968 592684 100020
rect 592736 100008 592742 100020
rect 667934 100008 667940 100020
rect 592736 99980 667940 100008
rect 592736 99968 592742 99980
rect 667934 99968 667940 99980
rect 667992 99968 667998 100020
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 579522 99220 579528 99272
rect 579580 99260 579586 99272
rect 583202 99260 583208 99272
rect 579580 99232 583208 99260
rect 579580 99220 579586 99232
rect 583202 99220 583208 99232
rect 583260 99220 583266 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 624602 99016 624608 99068
rect 624660 99056 624666 99068
rect 634998 99056 635004 99068
rect 624660 99028 635004 99056
rect 624660 99016 624666 99028
rect 634998 99016 635004 99028
rect 635056 99016 635062 99068
rect 625062 98880 625068 98932
rect 625120 98920 625126 98932
rect 636286 98920 636292 98932
rect 625120 98892 636292 98920
rect 625120 98880 625126 98892
rect 636286 98880 636292 98892
rect 636344 98880 636350 98932
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 647142 98744 647148 98796
rect 647200 98784 647206 98796
rect 661954 98784 661960 98796
rect 647200 98756 661960 98784
rect 647200 98744 647206 98756
rect 661954 98744 661960 98756
rect 662012 98744 662018 98796
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 646590 98648 646596 98660
rect 630548 98620 646596 98648
rect 630548 98608 630554 98620
rect 646590 98608 646596 98620
rect 646648 98608 646654 98660
rect 631410 98268 631416 98320
rect 631468 98308 631474 98320
rect 642174 98308 642180 98320
rect 631468 98280 642180 98308
rect 631468 98268 631474 98280
rect 642174 98268 642180 98280
rect 642232 98268 642238 98320
rect 633618 98132 633624 98184
rect 633676 98172 633682 98184
rect 640702 98172 640708 98184
rect 633676 98144 640708 98172
rect 633676 98132 633682 98144
rect 640702 98132 640708 98144
rect 640760 98132 640766 98184
rect 631980 98076 632192 98104
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625798 97968 625804 97980
rect 618772 97940 625804 97968
rect 618772 97928 618778 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 629754 97928 629760 97980
rect 629812 97968 629818 97980
rect 631980 97968 632008 98076
rect 632164 98036 632192 98076
rect 645302 98036 645308 98048
rect 632164 98008 645308 98036
rect 645302 97996 645308 98008
rect 645360 97996 645366 98048
rect 629812 97940 632008 97968
rect 629812 97928 629818 97940
rect 659194 97928 659200 97980
rect 659252 97968 659258 97980
rect 664162 97968 664168 97980
rect 659252 97940 664168 97968
rect 659252 97928 659258 97940
rect 664162 97928 664168 97940
rect 664220 97928 664226 97980
rect 620186 97792 620192 97844
rect 620244 97832 620250 97844
rect 626350 97832 626356 97844
rect 620244 97804 626356 97832
rect 620244 97792 620250 97804
rect 626350 97792 626356 97804
rect 626408 97792 626414 97844
rect 628282 97792 628288 97844
rect 628340 97832 628346 97844
rect 631410 97832 631416 97844
rect 628340 97804 631416 97832
rect 628340 97792 628346 97804
rect 631410 97792 631416 97804
rect 631468 97792 631474 97844
rect 632698 97792 632704 97844
rect 632756 97832 632762 97844
rect 647694 97832 647700 97844
rect 632756 97804 647700 97832
rect 632756 97792 632762 97804
rect 647694 97792 647700 97804
rect 647752 97792 647758 97844
rect 653950 97792 653956 97844
rect 654008 97832 654014 97844
rect 654318 97832 654324 97844
rect 654008 97804 654324 97832
rect 654008 97792 654014 97804
rect 654318 97792 654324 97804
rect 654376 97792 654382 97844
rect 655422 97792 655428 97844
rect 655480 97832 655486 97844
rect 655480 97804 659792 97832
rect 655480 97792 655486 97804
rect 631226 97656 631232 97708
rect 631284 97696 631290 97708
rect 647326 97696 647332 97708
rect 631284 97668 647332 97696
rect 631284 97656 631290 97668
rect 647326 97656 647332 97668
rect 647384 97656 647390 97708
rect 651834 97656 651840 97708
rect 651892 97696 651898 97708
rect 659562 97696 659568 97708
rect 651892 97668 659568 97696
rect 651892 97656 651898 97668
rect 659562 97656 659568 97668
rect 659620 97656 659626 97708
rect 659764 97696 659792 97804
rect 659930 97792 659936 97844
rect 659988 97832 659994 97844
rect 665358 97832 665364 97844
rect 659988 97804 665364 97832
rect 659988 97792 659994 97804
rect 665358 97792 665364 97804
rect 665416 97792 665422 97844
rect 662506 97696 662512 97708
rect 659764 97668 662512 97696
rect 662506 97656 662512 97668
rect 662564 97656 662570 97708
rect 627546 97520 627552 97572
rect 627604 97560 627610 97572
rect 633618 97560 633624 97572
rect 627604 97532 633624 97560
rect 627604 97520 627610 97532
rect 633618 97520 633624 97532
rect 633676 97520 633682 97572
rect 633802 97520 633808 97572
rect 633860 97560 633866 97572
rect 637758 97560 637764 97572
rect 633860 97532 637764 97560
rect 633860 97520 633866 97532
rect 637758 97520 637764 97532
rect 637816 97520 637822 97572
rect 643002 97520 643008 97572
rect 643060 97560 643066 97572
rect 657998 97560 658004 97572
rect 643060 97532 658004 97560
rect 643060 97520 643066 97532
rect 657998 97520 658004 97532
rect 658056 97520 658062 97572
rect 658182 97520 658188 97572
rect 658240 97560 658246 97572
rect 663058 97560 663064 97572
rect 658240 97532 663064 97560
rect 658240 97520 658246 97532
rect 663058 97520 663064 97532
rect 663116 97520 663122 97572
rect 605466 97384 605472 97436
rect 605524 97424 605530 97436
rect 611906 97424 611912 97436
rect 605524 97396 611912 97424
rect 605524 97384 605530 97396
rect 611906 97384 611912 97396
rect 611964 97384 611970 97436
rect 612642 97384 612648 97436
rect 612700 97424 612706 97436
rect 620278 97424 620284 97436
rect 612700 97396 620284 97424
rect 612700 97384 612706 97396
rect 620278 97384 620284 97396
rect 620336 97384 620342 97436
rect 621658 97384 621664 97436
rect 621716 97424 621722 97436
rect 629294 97424 629300 97436
rect 621716 97396 629300 97424
rect 621716 97384 621722 97396
rect 629294 97384 629300 97396
rect 629352 97384 629358 97436
rect 631962 97384 631968 97436
rect 632020 97424 632026 97436
rect 648614 97424 648620 97436
rect 632020 97396 648620 97424
rect 632020 97384 632026 97396
rect 648614 97384 648620 97396
rect 648672 97384 648678 97436
rect 650362 97384 650368 97436
rect 650420 97424 650426 97436
rect 658274 97424 658280 97436
rect 650420 97396 658280 97424
rect 650420 97384 650426 97396
rect 658274 97384 658280 97396
rect 658332 97384 658338 97436
rect 623130 97248 623136 97300
rect 623188 97288 623194 97300
rect 632054 97288 632060 97300
rect 623188 97260 632060 97288
rect 623188 97248 623194 97260
rect 632054 97248 632060 97260
rect 632112 97248 632118 97300
rect 633250 97248 633256 97300
rect 633308 97288 633314 97300
rect 650546 97288 650552 97300
rect 633308 97260 650552 97288
rect 633308 97248 633314 97260
rect 650546 97248 650552 97260
rect 650604 97248 650610 97300
rect 656802 97180 656808 97232
rect 656860 97220 656866 97232
rect 661402 97220 661408 97232
rect 656860 97192 661408 97220
rect 656860 97180 656866 97192
rect 661402 97180 661408 97192
rect 661460 97180 661466 97232
rect 626074 97112 626080 97164
rect 626132 97152 626138 97164
rect 633802 97152 633808 97164
rect 626132 97124 633808 97152
rect 626132 97112 626138 97124
rect 633802 97112 633808 97124
rect 633860 97112 633866 97164
rect 634170 97112 634176 97164
rect 634228 97152 634234 97164
rect 649074 97152 649080 97164
rect 634228 97124 649080 97152
rect 634228 97112 634234 97124
rect 649074 97112 649080 97124
rect 649132 97112 649138 97164
rect 657998 97044 658004 97096
rect 658056 97084 658062 97096
rect 659838 97084 659844 97096
rect 658056 97056 659844 97084
rect 658056 97044 658062 97056
rect 659838 97044 659844 97056
rect 659896 97044 659902 97096
rect 634722 96976 634728 97028
rect 634780 97016 634786 97028
rect 647142 97016 647148 97028
rect 634780 96988 647148 97016
rect 634780 96976 634786 96988
rect 647142 96976 647148 96988
rect 647200 96976 647206 97028
rect 597646 96908 597652 96960
rect 597704 96948 597710 96960
rect 598198 96948 598204 96960
rect 597704 96920 598204 96948
rect 597704 96908 597710 96920
rect 598198 96908 598204 96920
rect 598256 96908 598262 96960
rect 598934 96908 598940 96960
rect 598992 96948 598998 96960
rect 599670 96948 599676 96960
rect 598992 96920 599676 96948
rect 598992 96908 598998 96920
rect 599670 96908 599676 96920
rect 599728 96908 599734 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 607122 96948 607128 96960
rect 606260 96920 607128 96948
rect 606260 96908 606266 96920
rect 607122 96908 607128 96920
rect 607180 96908 607186 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 654778 96908 654784 96960
rect 654836 96948 654842 96960
rect 655422 96948 655428 96960
rect 654836 96920 655428 96948
rect 654836 96908 654842 96920
rect 655422 96908 655428 96920
rect 655480 96908 655486 96960
rect 656710 96908 656716 96960
rect 656768 96948 656774 96960
rect 660114 96948 660120 96960
rect 656768 96920 660120 96948
rect 656768 96908 656774 96920
rect 660114 96908 660120 96920
rect 660172 96908 660178 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 626810 96840 626816 96892
rect 626868 96880 626874 96892
rect 639230 96880 639236 96892
rect 626868 96852 639236 96880
rect 626868 96840 626874 96852
rect 639230 96840 639236 96852
rect 639288 96840 639294 96892
rect 644290 96772 644296 96824
rect 644348 96812 644354 96824
rect 658826 96812 658832 96824
rect 644348 96784 658832 96812
rect 644348 96772 644354 96784
rect 658826 96772 658832 96784
rect 658884 96772 658890 96824
rect 609146 96704 609152 96756
rect 609204 96744 609210 96756
rect 609698 96744 609704 96756
rect 609204 96716 609704 96744
rect 609204 96704 609210 96716
rect 609698 96704 609704 96716
rect 609756 96704 609762 96756
rect 640058 96568 640064 96620
rect 640116 96608 640122 96620
rect 645118 96608 645124 96620
rect 640116 96580 645124 96608
rect 640116 96568 640122 96580
rect 645118 96568 645124 96580
rect 645176 96568 645182 96620
rect 646406 96568 646412 96620
rect 646464 96608 646470 96620
rect 652202 96608 652208 96620
rect 646464 96580 652208 96608
rect 646464 96568 646470 96580
rect 652202 96568 652208 96580
rect 652260 96568 652266 96620
rect 652570 96568 652576 96620
rect 652628 96608 652634 96620
rect 664346 96608 664352 96620
rect 652628 96580 664352 96608
rect 652628 96568 652634 96580
rect 664346 96568 664352 96580
rect 664404 96568 664410 96620
rect 638586 96432 638592 96484
rect 638644 96472 638650 96484
rect 641346 96472 641352 96484
rect 638644 96444 641352 96472
rect 638644 96432 638650 96444
rect 641346 96432 641352 96444
rect 641404 96432 641410 96484
rect 641530 96432 641536 96484
rect 641588 96472 641594 96484
rect 648430 96472 648436 96484
rect 641588 96444 648436 96472
rect 641588 96432 641594 96444
rect 648430 96432 648436 96444
rect 648488 96432 648494 96484
rect 648890 96432 648896 96484
rect 648948 96472 648954 96484
rect 664530 96472 664536 96484
rect 648948 96444 664536 96472
rect 648948 96432 648954 96444
rect 664530 96432 664536 96444
rect 664588 96432 664594 96484
rect 637574 96296 637580 96348
rect 637632 96336 637638 96348
rect 660666 96336 660672 96348
rect 637632 96308 660672 96336
rect 637632 96296 637638 96308
rect 660666 96296 660672 96308
rect 660724 96296 660730 96348
rect 644934 96160 644940 96212
rect 644992 96200 644998 96212
rect 648062 96200 648068 96212
rect 644992 96172 648068 96200
rect 644992 96160 644998 96172
rect 648062 96160 648068 96172
rect 648120 96160 648126 96212
rect 648430 96160 648436 96212
rect 648488 96200 648494 96212
rect 663794 96200 663800 96212
rect 648488 96172 663800 96200
rect 648488 96160 648494 96172
rect 663794 96160 663800 96172
rect 663852 96160 663858 96212
rect 591298 96024 591304 96076
rect 591356 96064 591362 96076
rect 602614 96064 602620 96076
rect 591356 96036 602620 96064
rect 591356 96024 591362 96036
rect 602614 96024 602620 96036
rect 602672 96024 602678 96076
rect 610618 96024 610624 96076
rect 610676 96064 610682 96076
rect 621658 96064 621664 96076
rect 610676 96036 621664 96064
rect 610676 96024 610682 96036
rect 621658 96024 621664 96036
rect 621716 96024 621722 96076
rect 640518 96024 640524 96076
rect 640576 96064 640582 96076
rect 645578 96064 645584 96076
rect 640576 96036 645584 96064
rect 640576 96024 640582 96036
rect 645578 96024 645584 96036
rect 645636 96024 645642 96076
rect 647510 96024 647516 96076
rect 647568 96064 647574 96076
rect 663978 96064 663984 96076
rect 647568 96036 663984 96064
rect 647568 96024 647574 96036
rect 663978 96024 663984 96036
rect 664036 96024 664042 96076
rect 594058 95888 594064 95940
rect 594116 95928 594122 95940
rect 668026 95928 668032 95940
rect 594116 95900 668032 95928
rect 594116 95888 594122 95900
rect 668026 95888 668032 95900
rect 668084 95888 668090 95940
rect 639046 95752 639052 95804
rect 639104 95792 639110 95804
rect 648614 95792 648620 95804
rect 639104 95764 648620 95792
rect 639104 95752 639110 95764
rect 648614 95752 648620 95764
rect 648672 95752 648678 95804
rect 653306 95752 653312 95804
rect 653364 95792 653370 95804
rect 665174 95792 665180 95804
rect 653364 95764 665180 95792
rect 653364 95752 653370 95764
rect 665174 95752 665180 95764
rect 665232 95752 665238 95804
rect 645118 95616 645124 95668
rect 645176 95656 645182 95668
rect 652018 95656 652024 95668
rect 645176 95628 652024 95656
rect 645176 95616 645182 95628
rect 652018 95616 652024 95628
rect 652076 95616 652082 95668
rect 652386 95616 652392 95668
rect 652444 95656 652450 95668
rect 656342 95656 656348 95668
rect 652444 95628 656348 95656
rect 652444 95616 652450 95628
rect 656342 95616 656348 95628
rect 656400 95616 656406 95668
rect 648062 95480 648068 95532
rect 648120 95520 648126 95532
rect 656158 95520 656164 95532
rect 648120 95492 656164 95520
rect 648120 95480 648126 95492
rect 656158 95480 656164 95492
rect 656216 95480 656222 95532
rect 641346 95412 641352 95464
rect 641404 95412 641410 95464
rect 643462 95412 643468 95464
rect 643520 95452 643526 95464
rect 647878 95452 647884 95464
rect 643520 95424 647884 95452
rect 643520 95412 643526 95424
rect 647878 95412 647884 95424
rect 647936 95412 647942 95464
rect 641364 95316 641392 95412
rect 641364 95288 646958 95316
rect 578326 95140 578332 95192
rect 578384 95180 578390 95192
rect 584582 95180 584588 95192
rect 578384 95152 584588 95180
rect 578384 95140 578390 95152
rect 584582 95140 584588 95152
rect 584640 95140 584646 95192
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 625430 95180 625436 95192
rect 620980 95152 625436 95180
rect 620980 95140 620986 95152
rect 625430 95140 625436 95152
rect 625488 95140 625494 95192
rect 646930 95180 646958 95288
rect 647510 95276 647516 95328
rect 647568 95316 647574 95328
rect 652386 95316 652392 95328
rect 647568 95288 652392 95316
rect 647568 95276 647574 95288
rect 652386 95276 652392 95288
rect 652444 95276 652450 95328
rect 647510 95180 647516 95192
rect 646930 95152 647516 95180
rect 647510 95140 647516 95152
rect 647568 95140 647574 95192
rect 650270 95180 650276 95192
rect 649966 95152 650276 95180
rect 647142 95004 647148 95056
rect 647200 95044 647206 95056
rect 649966 95044 649994 95152
rect 650270 95140 650276 95152
rect 650328 95140 650334 95192
rect 647200 95016 649994 95044
rect 647200 95004 647206 95016
rect 616506 94936 616512 94988
rect 616564 94976 616570 94988
rect 624970 94976 624976 94988
rect 616564 94948 624976 94976
rect 616564 94936 616570 94948
rect 624970 94936 624976 94948
rect 625028 94936 625034 94988
rect 607674 94460 607680 94512
rect 607732 94500 607738 94512
rect 620830 94500 620836 94512
rect 607732 94472 620836 94500
rect 607732 94460 607738 94472
rect 620830 94460 620836 94472
rect 620888 94460 620894 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626166 93820 626172 93832
rect 619600 93792 626172 93820
rect 619600 93780 619606 93792
rect 626166 93780 626172 93792
rect 626224 93780 626230 93832
rect 651282 93576 651288 93628
rect 651340 93616 651346 93628
rect 654686 93616 654692 93628
rect 651340 93588 654692 93616
rect 651340 93576 651346 93588
rect 654686 93576 654692 93588
rect 654744 93576 654750 93628
rect 579246 93372 579252 93424
rect 579304 93412 579310 93424
rect 586146 93412 586152 93424
rect 579304 93384 586152 93412
rect 579304 93372 579310 93384
rect 586146 93372 586152 93384
rect 586204 93372 586210 93424
rect 609698 93100 609704 93152
rect 609756 93140 609762 93152
rect 618622 93140 618628 93152
rect 609756 93112 618628 93140
rect 609756 93100 609762 93112
rect 618622 93100 618628 93112
rect 618680 93100 618686 93152
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 647510 92420 647516 92472
rect 647568 92460 647574 92472
rect 655422 92460 655428 92472
rect 647568 92432 655428 92460
rect 647568 92420 647574 92432
rect 655422 92420 655428 92432
rect 655480 92420 655486 92472
rect 606938 91740 606944 91792
rect 606996 91780 607002 91792
rect 622394 91780 622400 91792
rect 606996 91752 622400 91780
rect 606996 91740 607002 91752
rect 622394 91740 622400 91752
rect 622452 91740 622458 91792
rect 578602 91128 578608 91180
rect 578660 91168 578666 91180
rect 585778 91168 585784 91180
rect 578660 91140 585784 91168
rect 578660 91128 578666 91140
rect 585778 91128 585784 91140
rect 585836 91128 585842 91180
rect 618162 91128 618168 91180
rect 618220 91168 618226 91180
rect 618220 91140 618392 91168
rect 618220 91128 618226 91140
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 618162 91032 618168 91044
rect 611320 91004 618168 91032
rect 611320 90992 611326 91004
rect 618162 90992 618168 91004
rect 618220 90992 618226 91044
rect 618364 91032 618392 91140
rect 626442 91032 626448 91044
rect 618364 91004 626448 91032
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 648614 90788 648620 90840
rect 648672 90828 648678 90840
rect 655422 90828 655428 90840
rect 648672 90800 655428 90828
rect 648672 90788 648678 90800
rect 655422 90788 655428 90800
rect 655480 90788 655486 90840
rect 620830 89632 620836 89684
rect 620888 89672 620894 89684
rect 626442 89672 626448 89684
rect 620888 89644 626448 89672
rect 620888 89632 620894 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 664162 88788 664168 88800
rect 662380 88760 664168 88788
rect 662380 88748 662386 88760
rect 664162 88748 664168 88760
rect 664220 88748 664226 88800
rect 656342 88612 656348 88664
rect 656400 88652 656406 88664
rect 657446 88652 657452 88664
rect 656400 88624 657452 88652
rect 656400 88612 656406 88624
rect 657446 88612 657452 88624
rect 657504 88612 657510 88664
rect 579246 88272 579252 88324
rect 579304 88312 579310 88324
rect 589918 88312 589924 88324
rect 579304 88284 589924 88312
rect 579304 88272 579310 88284
rect 589918 88272 589924 88284
rect 589976 88272 589982 88324
rect 622394 88272 622400 88324
rect 622452 88312 622458 88324
rect 626442 88312 626448 88324
rect 622452 88284 626448 88312
rect 622452 88272 622458 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 618162 88136 618168 88188
rect 618220 88176 618226 88188
rect 626258 88176 626264 88188
rect 618220 88148 626264 88176
rect 618220 88136 618226 88148
rect 626258 88136 626264 88148
rect 626316 88136 626322 88188
rect 648246 86980 648252 87032
rect 648304 87020 648310 87032
rect 662506 87020 662512 87032
rect 648304 86992 662512 87020
rect 648304 86980 648310 86992
rect 662506 86980 662512 86992
rect 662564 86980 662570 87032
rect 578326 86912 578332 86964
rect 578384 86952 578390 86964
rect 580442 86952 580448 86964
rect 578384 86924 580448 86952
rect 578384 86912 578390 86924
rect 580442 86912 580448 86924
rect 580500 86912 580506 86964
rect 656710 86844 656716 86896
rect 656768 86884 656774 86896
rect 659562 86884 659568 86896
rect 656768 86856 659568 86884
rect 656768 86844 656774 86856
rect 659562 86844 659568 86856
rect 659620 86844 659626 86896
rect 656158 86708 656164 86760
rect 656216 86748 656222 86760
rect 660666 86748 660672 86760
rect 656216 86720 660672 86748
rect 656216 86708 656222 86720
rect 660666 86708 660672 86720
rect 660724 86708 660730 86760
rect 652018 86572 652024 86624
rect 652076 86612 652082 86624
rect 660114 86612 660120 86624
rect 652076 86584 660120 86612
rect 652076 86572 652082 86584
rect 660114 86572 660120 86584
rect 660172 86572 660178 86624
rect 652202 86436 652208 86488
rect 652260 86476 652266 86488
rect 657170 86476 657176 86488
rect 652260 86448 657176 86476
rect 652260 86436 652266 86448
rect 657170 86436 657176 86448
rect 657228 86436 657234 86488
rect 621658 86300 621664 86352
rect 621716 86340 621722 86352
rect 626442 86340 626448 86352
rect 621716 86312 626448 86340
rect 621716 86300 621722 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 647878 86300 647884 86352
rect 647936 86340 647942 86352
rect 661402 86340 661408 86352
rect 647936 86312 661408 86340
rect 647936 86300 647942 86312
rect 661402 86300 661408 86312
rect 661460 86300 661466 86352
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 618622 85348 618628 85400
rect 618680 85388 618686 85400
rect 625246 85388 625252 85400
rect 618680 85360 625252 85388
rect 618680 85348 618686 85360
rect 625246 85348 625252 85360
rect 625304 85348 625310 85400
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 626442 84164 626448 84176
rect 608560 84136 626448 84164
rect 608560 84124 608566 84136
rect 626442 84124 626448 84136
rect 626500 84124 626506 84176
rect 579246 83988 579252 84040
rect 579304 84028 579310 84040
rect 581638 84028 581644 84040
rect 579304 84000 581644 84028
rect 579304 83988 579310 84000
rect 581638 83988 581644 84000
rect 581696 83988 581702 84040
rect 578878 82764 578884 82816
rect 578936 82804 578942 82816
rect 583018 82804 583024 82816
rect 578936 82776 583024 82804
rect 578936 82764 578942 82776
rect 583018 82764 583024 82776
rect 583076 82764 583082 82816
rect 579246 82084 579252 82136
rect 579304 82124 579310 82136
rect 587158 82124 587164 82136
rect 579304 82096 587164 82124
rect 579304 82084 579310 82096
rect 587158 82084 587164 82096
rect 587216 82084 587222 82136
rect 628742 81064 628748 81116
rect 628800 81104 628806 81116
rect 642450 81104 642456 81116
rect 628800 81076 642456 81104
rect 628800 81064 628806 81076
rect 642450 81064 642456 81076
rect 642508 81064 642514 81116
rect 615402 80928 615408 80980
rect 615460 80968 615466 80980
rect 646314 80968 646320 80980
rect 615460 80940 646320 80968
rect 615460 80928 615466 80940
rect 646314 80928 646320 80940
rect 646372 80928 646378 80980
rect 613838 80792 613844 80844
rect 613896 80832 613902 80844
rect 647326 80832 647332 80844
rect 613896 80804 647332 80832
rect 613896 80792 613902 80804
rect 647326 80792 647332 80804
rect 647384 80792 647390 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 614022 79432 614028 79484
rect 614080 79472 614086 79484
rect 646038 79472 646044 79484
rect 614080 79444 646044 79472
rect 614080 79432 614086 79444
rect 646038 79432 646044 79444
rect 646096 79432 646102 79484
rect 583018 79296 583024 79348
rect 583076 79336 583082 79348
rect 600498 79336 600504 79348
rect 583076 79308 600504 79336
rect 583076 79296 583082 79308
rect 600498 79296 600504 79308
rect 600556 79296 600562 79348
rect 612642 79296 612648 79348
rect 612700 79336 612706 79348
rect 648614 79336 648620 79348
rect 612700 79308 648620 79336
rect 612700 79296 612706 79308
rect 648614 79296 648620 79308
rect 648672 79296 648678 79348
rect 578234 78072 578240 78124
rect 578292 78112 578298 78124
rect 580258 78112 580264 78124
rect 578292 78084 580264 78112
rect 578292 78072 578298 78084
rect 580258 78072 580264 78084
rect 580316 78072 580322 78124
rect 633434 78072 633440 78124
rect 633492 78112 633498 78124
rect 645302 78112 645308 78124
rect 633492 78084 645308 78112
rect 633492 78072 633498 78084
rect 645302 78072 645308 78084
rect 645360 78072 645366 78124
rect 631042 77936 631048 77988
rect 631100 77976 631106 77988
rect 643094 77976 643100 77988
rect 631100 77948 643100 77976
rect 631100 77936 631106 77948
rect 643094 77936 643100 77948
rect 643152 77936 643158 77988
rect 628466 77664 628472 77716
rect 628524 77704 628530 77716
rect 632790 77704 632796 77716
rect 628524 77676 632796 77704
rect 628524 77664 628530 77676
rect 632790 77664 632796 77676
rect 632848 77664 632854 77716
rect 624418 77392 624424 77444
rect 624476 77432 624482 77444
rect 628466 77432 628472 77444
rect 624476 77404 628472 77432
rect 624476 77392 624482 77404
rect 628466 77392 628472 77404
rect 628524 77392 628530 77444
rect 625798 77256 625804 77308
rect 625856 77296 625862 77308
rect 631042 77296 631048 77308
rect 625856 77268 631048 77296
rect 625856 77256 625862 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 620278 76780 620284 76832
rect 620336 76820 620342 76832
rect 648982 76820 648988 76832
rect 620336 76792 648988 76820
rect 620336 76780 620342 76792
rect 648982 76780 648988 76792
rect 649040 76780 649046 76832
rect 611998 76644 612004 76696
rect 612056 76684 612062 76696
rect 662414 76684 662420 76696
rect 612056 76656 662420 76684
rect 612056 76644 612062 76656
rect 662414 76644 662420 76656
rect 662472 76644 662478 76696
rect 587158 76508 587164 76560
rect 587216 76548 587222 76560
rect 668210 76548 668216 76560
rect 587216 76520 668216 76548
rect 587216 76508 587222 76520
rect 668210 76508 668216 76520
rect 668268 76508 668274 76560
rect 616782 75420 616788 75472
rect 616840 75460 616846 75472
rect 646682 75460 646688 75472
rect 616840 75432 646688 75460
rect 616840 75420 616846 75432
rect 646682 75420 646688 75432
rect 646740 75420 646746 75472
rect 607122 75284 607128 75336
rect 607180 75324 607186 75336
rect 646498 75324 646504 75336
rect 607180 75296 646504 75324
rect 607180 75284 607186 75296
rect 646498 75284 646504 75296
rect 646556 75284 646562 75336
rect 578878 75148 578884 75200
rect 578936 75188 578942 75200
rect 666554 75188 666560 75200
rect 578936 75160 666560 75188
rect 578936 75148 578942 75160
rect 666554 75148 666560 75160
rect 666612 75148 666618 75200
rect 579522 73108 579528 73160
rect 579580 73148 579586 73160
rect 588538 73148 588544 73160
rect 579580 73120 588544 73148
rect 579580 73108 579586 73120
rect 588538 73108 588544 73120
rect 588596 73108 588602 73160
rect 578510 71544 578516 71596
rect 578568 71584 578574 71596
rect 584398 71584 584404 71596
rect 578568 71556 584404 71584
rect 578568 71544 578574 71556
rect 584398 71544 584404 71556
rect 584456 71544 584462 71596
rect 579522 66852 579528 66904
rect 579580 66892 579586 66904
rect 625982 66892 625988 66904
rect 579580 66864 625988 66892
rect 579580 66852 579586 66864
rect 625982 66852 625988 66864
rect 626040 66852 626046 66904
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 592678 64852 592684 64864
rect 579580 64824 592684 64852
rect 579580 64812 579586 64824
rect 592678 64812 592684 64824
rect 592736 64812 592742 64864
rect 579522 62024 579528 62076
rect 579580 62064 579586 62076
rect 587158 62064 587164 62076
rect 579580 62036 587164 62064
rect 579580 62024 579586 62036
rect 587158 62024 587164 62036
rect 587216 62024 587222 62076
rect 578326 59984 578332 60036
rect 578384 60024 578390 60036
rect 624418 60024 624424 60036
rect 578384 59996 624424 60024
rect 578384 59984 578390 59996
rect 624418 59984 624424 59996
rect 624476 59984 624482 60036
rect 577498 58760 577504 58812
rect 577556 58800 577562 58812
rect 604454 58800 604460 58812
rect 577556 58772 604460 58800
rect 577556 58760 577562 58772
rect 604454 58760 604460 58772
rect 604512 58760 604518 58812
rect 576118 58624 576124 58676
rect 576176 58664 576182 58676
rect 603074 58664 603080 58676
rect 576176 58636 603080 58664
rect 576176 58624 576182 58636
rect 603074 58624 603080 58636
rect 603132 58624 603138 58676
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 594058 57916 594064 57928
rect 579580 57888 594064 57916
rect 579580 57876 579586 57888
rect 594058 57876 594064 57888
rect 594116 57876 594122 57928
rect 574922 57196 574928 57248
rect 574980 57236 574986 57248
rect 600314 57236 600320 57248
rect 574980 57208 600320 57236
rect 574980 57196 574986 57208
rect 600314 57196 600320 57208
rect 600372 57196 600378 57248
rect 574738 55972 574744 56024
rect 574796 56012 574802 56024
rect 598934 56012 598940 56024
rect 574796 55984 598940 56012
rect 574796 55972 574802 55984
rect 598934 55972 598940 55984
rect 598992 55972 598998 56024
rect 574462 55836 574468 55888
rect 574520 55876 574526 55888
rect 601878 55876 601884 55888
rect 574520 55848 601884 55876
rect 574520 55836 574526 55848
rect 601878 55836 601884 55848
rect 601936 55836 601942 55888
rect 463344 55440 481634 55468
rect 463344 53644 463372 55440
rect 463804 55304 473354 55332
rect 463804 53768 463832 55304
rect 473326 55264 473354 55304
rect 478846 55304 479288 55332
rect 478846 55264 478874 55304
rect 473326 55236 478874 55264
rect 473326 55100 478874 55128
rect 473326 54924 473354 55100
rect 471164 54896 473354 54924
rect 478846 54924 478874 55100
rect 479260 55060 479288 55304
rect 481606 55196 481634 55440
rect 596450 55196 596456 55208
rect 481606 55168 596456 55196
rect 596450 55156 596456 55168
rect 596508 55156 596514 55208
rect 597830 55060 597836 55072
rect 479260 55032 597836 55060
rect 597830 55020 597836 55032
rect 597888 55020 597894 55072
rect 597646 54924 597652 54936
rect 478846 54896 597652 54924
rect 466426 53808 471008 53836
rect 466426 53768 466454 53808
rect 463804 53740 464108 53768
rect 464080 53644 464108 53740
rect 464218 53740 466454 53768
rect 463326 53592 463332 53644
rect 463384 53592 463390 53644
rect 463510 53592 463516 53644
rect 463568 53632 463574 53644
rect 463878 53632 463884 53644
rect 463568 53604 463884 53632
rect 463568 53592 463574 53604
rect 463878 53592 463884 53604
rect 463936 53592 463942 53644
rect 464062 53592 464068 53644
rect 464120 53592 464126 53644
rect 460382 53456 460388 53508
rect 460440 53496 460446 53508
rect 464218 53496 464246 53740
rect 470980 53644 471008 53808
rect 471164 53644 471192 54896
rect 597646 54884 597652 54896
rect 597704 54884 597710 54936
rect 599118 54788 599124 54800
rect 471900 54760 478920 54788
rect 471900 53904 471928 54760
rect 478892 54720 478920 54760
rect 479260 54760 599124 54788
rect 479260 54720 479288 54760
rect 599118 54748 599124 54760
rect 599176 54748 599182 54800
rect 478892 54692 479288 54720
rect 623038 54652 623044 54664
rect 479352 54624 623044 54652
rect 479352 54584 479380 54624
rect 623038 54612 623044 54624
rect 623096 54612 623102 54664
rect 474016 54556 479380 54584
rect 474016 53904 474044 54556
rect 625798 54516 625804 54528
rect 479444 54488 625804 54516
rect 479444 54448 479472 54488
rect 625798 54476 625804 54488
rect 625856 54476 625862 54528
rect 471716 53876 471928 53904
rect 472084 53876 474044 53904
rect 476776 54420 479472 54448
rect 471716 53644 471744 53876
rect 472084 53768 472112 53876
rect 471992 53740 472112 53768
rect 471992 53644 472020 53740
rect 476776 53644 476804 54420
rect 596266 54380 596272 54392
rect 479536 54352 596272 54380
rect 479536 54312 479564 54352
rect 596266 54340 596272 54352
rect 596324 54340 596330 54392
rect 479444 54284 479564 54312
rect 465902 53592 465908 53644
rect 465960 53632 465966 53644
rect 470318 53632 470324 53644
rect 465960 53604 470324 53632
rect 465960 53592 465966 53604
rect 470318 53592 470324 53604
rect 470376 53592 470382 53644
rect 470962 53592 470968 53644
rect 471020 53592 471026 53644
rect 471146 53592 471152 53644
rect 471204 53592 471210 53644
rect 471698 53592 471704 53644
rect 471756 53592 471762 53644
rect 471974 53592 471980 53644
rect 472032 53592 472038 53644
rect 476758 53592 476764 53644
rect 476816 53592 476822 53644
rect 479444 53632 479472 54284
rect 583018 54244 583024 54256
rect 479628 54216 583024 54244
rect 479628 53644 479656 54216
rect 583018 54204 583024 54216
rect 583076 54204 583082 54256
rect 580442 54108 580448 54120
rect 480088 54080 580448 54108
rect 480088 53768 480116 54080
rect 580442 54068 580448 54080
rect 580500 54068 580506 54120
rect 574738 53972 574744 53984
rect 479996 53740 480116 53768
rect 480180 53944 574744 53972
rect 479996 53644 480024 53740
rect 480180 53644 480208 53944
rect 574738 53932 574744 53944
rect 574796 53932 574802 53984
rect 574922 53836 574928 53848
rect 482986 53808 574928 53836
rect 476960 53604 479472 53632
rect 460440 53468 464246 53496
rect 460440 53456 460446 53468
rect 464982 53456 464988 53508
rect 465040 53496 465046 53508
rect 476960 53496 476988 53604
rect 479610 53592 479616 53644
rect 479668 53592 479674 53644
rect 479978 53592 479984 53644
rect 480036 53592 480042 53644
rect 480162 53592 480168 53644
rect 480220 53592 480226 53644
rect 465040 53468 476988 53496
rect 465040 53456 465046 53468
rect 477972 53400 478184 53428
rect 50522 53320 50528 53372
rect 50580 53360 50586 53372
rect 130378 53360 130384 53372
rect 50580 53332 130384 53360
rect 50580 53320 50586 53332
rect 130378 53320 130384 53332
rect 130436 53320 130442 53372
rect 462222 53320 462228 53372
rect 462280 53360 462286 53372
rect 477972 53360 478000 53400
rect 462280 53332 478000 53360
rect 478156 53360 478184 53400
rect 482986 53360 483014 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 478156 53332 483014 53360
rect 462280 53320 462286 53332
rect 48958 53184 48964 53236
rect 49016 53224 49022 53236
rect 128998 53224 129004 53236
rect 49016 53196 129004 53224
rect 49016 53184 49022 53196
rect 128998 53184 129004 53196
rect 129056 53184 129062 53236
rect 463142 53184 463148 53236
rect 463200 53224 463206 53236
rect 479610 53224 479616 53236
rect 463200 53196 479616 53224
rect 463200 53184 463206 53196
rect 479610 53184 479616 53196
rect 479668 53184 479674 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 47578 53048 47584 53100
rect 47636 53088 47642 53100
rect 129182 53088 129188 53100
rect 47636 53060 129188 53088
rect 47636 53048 47642 53060
rect 129182 53048 129188 53060
rect 129240 53048 129246 53100
rect 461302 53048 461308 53100
rect 461360 53088 461366 53100
rect 480162 53088 480168 53100
rect 461360 53060 480168 53088
rect 461360 53048 461366 53060
rect 480162 53048 480168 53060
rect 480220 53048 480226 53100
rect 463326 52912 463332 52964
rect 463384 52952 463390 52964
rect 463786 52952 463792 52964
rect 463384 52924 463792 52952
rect 463384 52912 463390 52924
rect 463786 52912 463792 52924
rect 463844 52912 463850 52964
rect 459140 52776 459146 52828
rect 459198 52816 459204 52828
rect 459198 52788 463694 52816
rect 459198 52776 459204 52788
rect 463666 52680 463694 52788
rect 465120 52776 465126 52828
rect 465178 52816 465184 52828
rect 479978 52816 479984 52828
rect 465178 52788 479984 52816
rect 465178 52776 465184 52788
rect 479978 52776 479984 52788
rect 480036 52776 480042 52828
rect 471698 52680 471704 52692
rect 463666 52652 471704 52680
rect 471698 52640 471704 52652
rect 471756 52640 471762 52692
rect 50338 51824 50344 51876
rect 50396 51864 50402 51876
rect 129366 51864 129372 51876
rect 50396 51836 129372 51864
rect 50396 51824 50402 51836
rect 129366 51824 129372 51836
rect 129424 51824 129430 51876
rect 46198 51688 46204 51740
rect 46256 51728 46262 51740
rect 130562 51728 130568 51740
rect 46256 51700 130568 51728
rect 46256 51688 46262 51700
rect 130562 51688 130568 51700
rect 130620 51688 130626 51740
rect 145374 51688 145380 51740
rect 145432 51728 145438 51740
rect 306006 51728 306012 51740
rect 145432 51700 306012 51728
rect 145432 51688 145438 51700
rect 306006 51688 306012 51700
rect 306064 51688 306070 51740
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 49142 50328 49148 50380
rect 49200 50368 49206 50380
rect 131022 50368 131028 50380
rect 49200 50340 131028 50368
rect 49200 50328 49206 50340
rect 131022 50328 131028 50340
rect 131080 50328 131086 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 51718 49104 51724 49156
rect 51776 49144 51782 49156
rect 129642 49144 129648 49156
rect 51776 49116 129648 49144
rect 51776 49104 51782 49116
rect 129642 49104 129648 49116
rect 129700 49104 129706 49156
rect 45462 48968 45468 49020
rect 45520 49008 45526 49020
rect 128814 49008 128820 49020
rect 45520 48980 128820 49008
rect 45520 48968 45526 48980
rect 128814 48968 128820 48980
rect 128872 48968 128878 49020
rect 128814 47812 128820 47864
rect 128872 47852 128878 47864
rect 130746 47852 130752 47864
rect 128872 47824 130752 47852
rect 128872 47812 128878 47824
rect 130746 47812 130752 47824
rect 130804 47812 130810 47864
rect 625982 46452 625988 46504
rect 626040 46492 626046 46504
rect 661770 46492 661776 46504
rect 626040 46464 661776 46492
rect 626040 46452 626046 46464
rect 661770 46452 661776 46464
rect 661828 46452 661834 46504
rect 128998 46044 129004 46096
rect 129056 46084 129062 46096
rect 131758 46084 131764 46096
rect 129056 46056 131764 46084
rect 129056 46044 129062 46056
rect 131758 46044 131764 46056
rect 131816 46044 131822 46096
rect 130562 45908 130568 45960
rect 130620 45948 130626 45960
rect 132494 45948 132500 45960
rect 130620 45920 132500 45948
rect 130620 45908 130626 45920
rect 132494 45908 132500 45920
rect 132552 45908 132558 45960
rect 129642 45364 129648 45416
rect 129700 45404 129706 45416
rect 129700 45376 131206 45404
rect 129700 45364 129706 45376
rect 131178 45336 131206 45376
rect 131178 45308 131298 45336
rect 43806 45160 43812 45212
rect 43864 45200 43870 45212
rect 131114 45200 131120 45212
rect 43864 45172 131120 45200
rect 43864 45160 43870 45172
rect 131114 45160 131120 45172
rect 131172 45160 131178 45212
rect 131270 45090 131298 45308
rect 131390 45296 131396 45348
rect 131448 45336 131454 45348
rect 132954 45336 132960 45348
rect 131448 45308 132960 45336
rect 131448 45296 131454 45308
rect 132954 45296 132960 45308
rect 133012 45296 133018 45348
rect 131390 45160 131396 45212
rect 131448 45200 131454 45212
rect 133138 45200 133144 45212
rect 131448 45172 133144 45200
rect 131448 45160 131454 45172
rect 133138 45160 133144 45172
rect 133196 45160 133202 45212
rect 129366 45024 129372 45076
rect 129424 45064 129430 45076
rect 129424 45036 131068 45064
rect 129424 45024 129430 45036
rect 131040 45020 131068 45036
rect 131040 44992 131330 45020
rect 131592 44804 131620 44922
rect 131574 44752 131580 44804
rect 131632 44752 131638 44804
rect 131776 44696 131804 44838
rect 131758 44644 131764 44696
rect 131816 44644 131822 44696
rect 131960 44668 131988 44754
rect 131942 44616 131948 44668
rect 132000 44616 132006 44668
rect 129182 44480 129188 44532
rect 129240 44520 129246 44532
rect 129240 44492 132172 44520
rect 129240 44480 129246 44492
rect 132144 44452 132172 44492
rect 132236 44452 132264 44670
rect 132144 44424 132264 44452
rect 43622 44276 43628 44328
rect 43680 44316 43686 44328
rect 129090 44316 129096 44328
rect 43680 44288 129096 44316
rect 43680 44276 43686 44288
rect 129090 44276 129096 44288
rect 129148 44276 129154 44328
rect 130746 44276 130752 44328
rect 130804 44316 130810 44328
rect 132374 44316 132402 44586
rect 132466 44488 132526 44516
rect 132466 44396 132494 44488
rect 132466 44356 132500 44396
rect 132494 44344 132500 44356
rect 132552 44344 132558 44396
rect 130804 44288 132402 44316
rect 130804 44276 130810 44288
rect 43438 44140 43444 44192
rect 43496 44180 43502 44192
rect 131574 44180 131580 44192
rect 43496 44152 131580 44180
rect 43496 44140 43502 44152
rect 131574 44140 131580 44152
rect 131632 44140 131638 44192
rect 132742 44180 132770 44390
rect 132954 44252 132960 44304
rect 133012 44252 133018 44304
rect 131776 44152 132770 44180
rect 130378 44004 130384 44056
rect 130436 44044 130442 44056
rect 131776 44044 131804 44152
rect 133138 44140 133144 44192
rect 133196 44140 133202 44192
rect 130436 44016 131804 44044
rect 130436 44004 130442 44016
rect 440234 43596 440240 43648
rect 440292 43636 440298 43648
rect 441062 43636 441068 43648
rect 440292 43608 441068 43636
rect 440292 43596 440298 43608
rect 441062 43596 441068 43608
rect 441120 43596 441126 43648
rect 187326 42712 187332 42764
rect 187384 42752 187390 42764
rect 431218 42752 431224 42764
rect 187384 42724 431224 42752
rect 187384 42712 187390 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 441062 42712 441068 42764
rect 441120 42752 441126 42764
rect 449158 42752 449164 42764
rect 441120 42724 449164 42752
rect 441120 42712 441126 42724
rect 449158 42712 449164 42724
rect 449216 42712 449222 42764
rect 459554 42440 459560 42492
rect 459612 42480 459618 42492
rect 460106 42480 460112 42492
rect 459612 42452 460112 42480
rect 459612 42440 459618 42452
rect 460106 42440 460112 42452
rect 460164 42440 460170 42492
rect 454494 42304 454500 42356
rect 454552 42344 454558 42356
rect 463050 42344 463056 42356
rect 454552 42316 463056 42344
rect 454552 42304 454558 42316
rect 463050 42304 463056 42316
rect 463108 42304 463114 42356
rect 661402 42129 661408 42181
rect 661460 42129 661466 42181
rect 431218 41964 431224 42016
rect 431276 42004 431282 42016
rect 441062 42004 441068 42016
rect 431276 41976 441068 42004
rect 431276 41964 431282 41976
rect 441062 41964 441068 41976
rect 441120 41964 441126 42016
rect 449158 41964 449164 42016
rect 449216 42004 449222 42016
rect 459370 42004 459376 42016
rect 449216 41976 459376 42004
rect 449216 41964 449222 41976
rect 459370 41964 459376 41976
rect 459428 41964 459434 42016
rect 404630 41828 404636 41880
rect 404688 41828 404694 41880
rect 404648 41732 404676 41828
rect 420730 41732 420736 41744
rect 404648 41704 420736 41732
rect 420730 41692 420736 41704
rect 420788 41692 420794 41744
rect 427078 41692 427084 41744
rect 427136 41732 427142 41744
rect 459186 41732 459192 41744
rect 427136 41704 459192 41732
rect 427136 41692 427142 41704
rect 459186 41692 459192 41704
rect 459244 41692 459250 41744
rect 311066 41556 311072 41608
rect 311124 41596 311130 41608
rect 454494 41596 454500 41608
rect 311124 41568 454500 41596
rect 311124 41556 311130 41568
rect 454494 41556 454500 41568
rect 454552 41556 454558 41608
rect 420730 41420 420736 41472
rect 420788 41460 420794 41472
rect 427078 41460 427084 41472
rect 420788 41432 424272 41460
rect 420788 41420 420794 41432
rect 424244 41392 424272 41432
rect 424612 41432 427084 41460
rect 424612 41392 424640 41432
rect 427078 41420 427084 41432
rect 427136 41420 427142 41472
rect 424244 41364 424640 41392
<< via1 >>
rect 652024 896996 652076 897048
rect 676036 897064 676088 897116
rect 654784 895772 654836 895824
rect 675852 895772 675904 895824
rect 672724 895636 672776 895688
rect 676036 895636 676088 895688
rect 672540 894412 672592 894464
rect 675852 894412 675904 894464
rect 673368 894276 673420 894328
rect 676036 894276 676088 894328
rect 671988 892984 672040 893036
rect 676036 892984 676088 893036
rect 670884 892848 670936 892900
rect 675852 892848 675904 892900
rect 674932 890332 674984 890384
rect 676036 890332 676088 890384
rect 676220 890128 676272 890180
rect 676864 890128 676916 890180
rect 674472 888904 674524 888956
rect 676036 888904 676088 888956
rect 676220 888700 676272 888752
rect 677048 888700 677100 888752
rect 674288 887272 674340 887324
rect 676036 887272 676088 887324
rect 673184 886864 673236 886916
rect 676036 886864 676088 886916
rect 671804 885640 671856 885692
rect 676036 885640 676088 885692
rect 653404 880472 653456 880524
rect 675576 880472 675628 880524
rect 675944 880404 675996 880456
rect 679624 880404 679676 880456
rect 675392 879316 675444 879368
rect 676864 879316 676916 879368
rect 675760 879180 675812 879232
rect 678244 879180 678296 879232
rect 675208 879044 675260 879096
rect 676404 879044 676456 879096
rect 674794 878636 674846 878688
rect 677048 878636 677100 878688
rect 675944 878432 675996 878484
rect 675484 877752 675536 877804
rect 675208 874284 675260 874336
rect 675208 874148 675260 874200
rect 675024 874012 675076 874064
rect 675392 874012 675444 874064
rect 674840 873672 674892 873724
rect 675392 873672 675444 873724
rect 657544 869388 657596 869440
rect 675024 869388 675076 869440
rect 674840 869252 674892 869304
rect 675300 869252 675352 869304
rect 651472 868844 651524 868896
rect 654784 868844 654836 868896
rect 654140 868028 654192 868080
rect 675024 868028 675076 868080
rect 674840 867552 674892 867604
rect 675208 867552 675260 867604
rect 651472 866600 651524 866652
rect 672724 866600 672776 866652
rect 651380 865172 651432 865224
rect 653404 865172 653456 865224
rect 651472 863812 651524 863864
rect 657544 863812 657596 863864
rect 651472 862452 651524 862504
rect 654140 862452 654192 862504
rect 35624 817096 35676 817148
rect 35808 817096 35860 817148
rect 46204 817096 46256 817148
rect 61384 816960 61436 817012
rect 35624 815736 35676 815788
rect 44824 815736 44876 815788
rect 35808 815600 35860 815652
rect 45008 815600 45060 815652
rect 35624 814376 35676 814428
rect 44272 814376 44324 814428
rect 35808 814240 35860 814292
rect 44548 814240 44600 814292
rect 41328 812812 41380 812864
rect 43260 812812 43312 812864
rect 41144 810704 41196 810756
rect 42524 810704 42576 810756
rect 41144 807440 41196 807492
rect 43076 807440 43128 807492
rect 40960 807304 41012 807356
rect 45192 807304 45244 807356
rect 31760 806624 31812 806676
rect 35624 806624 35676 806676
rect 44824 806556 44876 806608
rect 62764 806556 62816 806608
rect 41328 805944 41380 805996
rect 43812 805944 43864 805996
rect 35624 802544 35676 802596
rect 33048 802408 33100 802460
rect 42156 802408 42208 802460
rect 42340 802408 42392 802460
rect 33784 801184 33836 801236
rect 40132 801184 40184 801236
rect 31024 801048 31076 801100
rect 43628 801048 43680 801100
rect 39304 800844 39356 800896
rect 41972 800844 42024 800896
rect 43444 799008 43496 799060
rect 53104 799008 53156 799060
rect 42524 797648 42576 797700
rect 57244 797648 57296 797700
rect 42892 796492 42944 796544
rect 43628 796492 43680 796544
rect 42432 794996 42484 795048
rect 43076 794996 43128 795048
rect 43076 794860 43128 794912
rect 45192 794860 45244 794912
rect 42432 794044 42484 794096
rect 43076 794044 43128 794096
rect 669228 790916 669280 790968
rect 675208 790916 675260 790968
rect 653404 790780 653456 790832
rect 675392 790780 675444 790832
rect 53104 790712 53156 790764
rect 62212 790712 62264 790764
rect 42248 789692 42300 789744
rect 42248 789488 42300 789540
rect 670608 789352 670660 789404
rect 675116 789352 675168 789404
rect 57244 789148 57296 789200
rect 62120 789148 62172 789200
rect 42616 786632 42668 786684
rect 62120 786632 62172 786684
rect 46204 785136 46256 785188
rect 62120 785136 62172 785188
rect 673000 783844 673052 783896
rect 675116 783844 675168 783896
rect 670424 782484 670476 782536
rect 675300 782484 675352 782536
rect 655520 781056 655572 781108
rect 675024 781056 675076 781108
rect 673552 779968 673604 780020
rect 675116 779968 675168 780020
rect 655152 778472 655204 778524
rect 675024 778472 675076 778524
rect 651472 777588 651524 777640
rect 660304 777588 660356 777640
rect 670240 776976 670292 777028
rect 675024 776976 675076 777028
rect 651472 775684 651524 775736
rect 669964 775684 670016 775736
rect 668400 775548 668452 775600
rect 675024 775548 675076 775600
rect 651380 775276 651432 775328
rect 653404 775276 653456 775328
rect 35808 774188 35860 774240
rect 41696 774188 41748 774240
rect 42064 774188 42116 774240
rect 60004 774188 60056 774240
rect 651472 774120 651524 774172
rect 655520 774120 655572 774172
rect 651472 773780 651524 773832
rect 655152 773780 655204 773832
rect 35808 773372 35860 773424
rect 40500 773372 40552 773424
rect 35532 773100 35584 773152
rect 40500 773100 40552 773152
rect 35348 772964 35400 773016
rect 41696 772964 41748 773016
rect 42064 772964 42116 773016
rect 46204 772964 46256 773016
rect 35164 772828 35216 772880
rect 61384 772828 61436 772880
rect 41696 772692 41748 772744
rect 42064 772692 42116 772744
rect 35808 771808 35860 771860
rect 39580 771808 39632 771860
rect 35624 771536 35676 771588
rect 41328 771604 41380 771656
rect 42064 771468 42116 771520
rect 44548 771468 44600 771520
rect 35808 771400 35860 771452
rect 41696 771400 41748 771452
rect 35808 770448 35860 770500
rect 40040 770448 40092 770500
rect 35624 770176 35676 770228
rect 40316 770176 40368 770228
rect 35808 770040 35860 770092
rect 41696 770040 41748 770092
rect 42064 770040 42116 770092
rect 44272 770040 44324 770092
rect 35808 768952 35860 769004
rect 39764 768952 39816 769004
rect 35532 768816 35584 768868
rect 40684 768816 40736 768868
rect 35348 768680 35400 768732
rect 41696 768680 41748 768732
rect 35808 767456 35860 767508
rect 36544 767456 36596 767508
rect 35624 767320 35676 767372
rect 41696 767252 41748 767304
rect 35808 766028 35860 766080
rect 39304 766028 39356 766080
rect 35808 764804 35860 764856
rect 40408 764804 40460 764856
rect 35808 764532 35860 764584
rect 41696 764532 41748 764584
rect 37096 763648 37148 763700
rect 39304 763648 39356 763700
rect 35808 763240 35860 763292
rect 41696 763240 41748 763292
rect 35808 761880 35860 761932
rect 39948 761880 40000 761932
rect 33048 760996 33100 761048
rect 41512 760996 41564 761048
rect 35164 759568 35216 759620
rect 40500 759500 40552 759552
rect 39304 757732 39356 757784
rect 41604 757732 41656 757784
rect 44732 755488 44784 755540
rect 62764 755488 62816 755540
rect 43444 754876 43496 754928
rect 45100 754876 45152 754928
rect 42340 753924 42392 753976
rect 43628 753924 43680 753976
rect 42248 753516 42300 753568
rect 45284 753516 45336 753568
rect 61384 746988 61436 747040
rect 62396 746988 62448 747040
rect 45100 746512 45152 746564
rect 62120 746512 62172 746564
rect 671068 745220 671120 745272
rect 675116 745220 675168 745272
rect 42524 743996 42576 744048
rect 62120 743860 62172 743912
rect 46204 743724 46256 743776
rect 62120 743724 62172 743776
rect 671344 743724 671396 743776
rect 675484 743724 675536 743776
rect 672356 742432 672408 742484
rect 675392 742432 675444 742484
rect 60004 742364 60056 742416
rect 62120 742364 62172 742416
rect 668768 741072 668820 741124
rect 675300 741072 675352 741124
rect 669780 739916 669832 739968
rect 675392 739916 675444 739968
rect 652024 736176 652076 736228
rect 653404 736176 653456 736228
rect 657544 735564 657596 735616
rect 672172 735700 672224 735752
rect 672172 734544 672224 734596
rect 675300 734544 675352 734596
rect 669596 734408 669648 734460
rect 675116 734408 675168 734460
rect 654784 734136 654836 734188
rect 675116 734272 675168 734324
rect 651472 733388 651524 733440
rect 668584 733388 668636 733440
rect 651472 732776 651524 732828
rect 661684 732776 661736 732828
rect 674472 731824 674524 731876
rect 675300 731824 675352 731876
rect 651472 731416 651524 731468
rect 658924 731416 658976 731468
rect 651472 731280 651524 731332
rect 671344 731280 671396 731332
rect 42064 731144 42116 731196
rect 61384 731144 61436 731196
rect 35808 731076 35860 731128
rect 41696 731076 41748 731128
rect 674840 731076 674892 731128
rect 675208 730872 675260 730924
rect 35808 730532 35860 730584
rect 39948 730532 40000 730584
rect 674840 730464 674892 730516
rect 675300 730464 675352 730516
rect 35624 730260 35676 730312
rect 41696 730260 41748 730312
rect 671252 730056 671304 730108
rect 675300 730056 675352 730108
rect 651472 729988 651524 730040
rect 657544 729988 657596 730040
rect 35440 729376 35492 729428
rect 41696 729376 41748 729428
rect 42064 729308 42116 729360
rect 62764 729308 62816 729360
rect 35808 729036 35860 729088
rect 41696 729036 41748 729088
rect 35624 728764 35676 728816
rect 39580 728764 39632 728816
rect 35256 728628 35308 728680
rect 41696 728628 41748 728680
rect 42064 728628 42116 728680
rect 43076 728628 43128 728680
rect 672724 728628 672776 728680
rect 675300 728628 675352 728680
rect 651472 728492 651524 728544
rect 654784 728492 654836 728544
rect 671804 728288 671856 728340
rect 673184 728084 673236 728136
rect 42064 727880 42116 727932
rect 44272 727880 44324 727932
rect 675852 727880 675904 727932
rect 683304 727880 683356 727932
rect 35808 727812 35860 727864
rect 41512 727812 41564 727864
rect 35624 727540 35676 727592
rect 40408 727540 40460 727592
rect 35808 727404 35860 727456
rect 41696 727404 41748 727456
rect 35808 727268 35860 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 45008 727268 45060 727320
rect 676036 726520 676088 726572
rect 683488 726520 683540 726572
rect 41328 726180 41380 726232
rect 41696 726180 41748 726232
rect 41144 725908 41196 725960
rect 41604 725908 41656 725960
rect 674380 721692 674432 721744
rect 675116 721692 675168 721744
rect 674380 721216 674432 721268
rect 675116 721216 675168 721268
rect 674380 720808 674432 720860
rect 675116 720808 675168 720860
rect 674380 720468 674432 720520
rect 675392 720468 675444 720520
rect 653404 716252 653456 716304
rect 674012 716252 674064 716304
rect 35164 715776 35216 715828
rect 41696 715776 41748 715828
rect 669964 715708 670016 715760
rect 673276 715708 673328 715760
rect 33784 715640 33836 715692
rect 37740 715640 37792 715692
rect 33048 715504 33100 715556
rect 39856 715504 39908 715556
rect 660304 714824 660356 714876
rect 674012 714892 674064 714944
rect 670884 713668 670936 713720
rect 674012 713668 674064 713720
rect 671344 713192 671396 713244
rect 674012 713192 674064 713244
rect 671988 712376 672040 712428
rect 674012 712376 674064 712428
rect 43628 712104 43680 712156
rect 50344 712104 50396 712156
rect 42248 711696 42300 711748
rect 42248 711084 42300 711136
rect 669228 710676 669280 710728
rect 674012 710676 674064 710728
rect 670424 710404 670476 710456
rect 674012 710404 674064 710456
rect 668400 709996 668452 710048
rect 674012 709996 674064 710048
rect 670608 709588 670660 709640
rect 674012 709588 674064 709640
rect 43628 709316 43680 709368
rect 44456 709316 44508 709368
rect 42248 709180 42300 709232
rect 44640 709180 44692 709232
rect 671620 707956 671672 708008
rect 674012 707956 674064 708008
rect 42616 707412 42668 707464
rect 42432 707072 42484 707124
rect 42616 706664 42668 706716
rect 42432 706596 42484 706648
rect 670240 705304 670292 705356
rect 674012 705304 674064 705356
rect 675852 705168 675904 705220
rect 683120 705168 683172 705220
rect 50344 705100 50396 705152
rect 62120 705100 62172 705152
rect 670608 703808 670660 703860
rect 674012 703808 674064 703860
rect 44456 703740 44508 703792
rect 62120 703740 62172 703792
rect 42708 701020 42760 701072
rect 62212 701020 62264 701072
rect 654784 701020 654836 701072
rect 673552 701020 673604 701072
rect 46204 698164 46256 698216
rect 62120 698164 62172 698216
rect 666468 697076 666520 697128
rect 673552 697076 673604 697128
rect 656808 690004 656860 690056
rect 673552 690004 673604 690056
rect 674288 690004 674340 690056
rect 675116 690004 675168 690056
rect 652760 688780 652812 688832
rect 673552 688780 673604 688832
rect 651656 688644 651708 688696
rect 660304 688644 660356 688696
rect 651472 687896 651524 687948
rect 667204 687896 667256 687948
rect 42708 687284 42760 687336
rect 61384 687216 61436 687268
rect 674472 687216 674524 687268
rect 675116 687216 675168 687268
rect 651472 687148 651524 687200
rect 654784 687148 654836 687200
rect 43444 686468 43496 686520
rect 62764 686468 62816 686520
rect 41144 685992 41196 686044
rect 41696 685992 41748 686044
rect 42064 685992 42116 686044
rect 44640 685992 44692 686044
rect 670240 685924 670292 685976
rect 673184 685924 673236 685976
rect 40868 685856 40920 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 45192 685856 45244 685908
rect 651472 685516 651524 685568
rect 656808 685516 656860 685568
rect 41052 684700 41104 684752
rect 41696 684700 41748 684752
rect 40868 684564 40920 684616
rect 41696 684496 41748 684548
rect 42064 684496 42116 684548
rect 45192 684496 45244 684548
rect 41328 683408 41380 683460
rect 41696 683408 41748 683460
rect 675852 682524 675904 682576
rect 683212 682524 683264 682576
rect 683396 682388 683448 682440
rect 675852 682252 675904 682304
rect 40960 679124 41012 679176
rect 41328 679124 41380 679176
rect 41144 678988 41196 679040
rect 41696 678988 41748 679040
rect 42064 678988 42116 679040
rect 45008 678988 45060 679040
rect 40960 677696 41012 677748
rect 41604 677696 41656 677748
rect 35164 672868 35216 672920
rect 38936 672868 38988 672920
rect 33784 672732 33836 672784
rect 38200 672732 38252 672784
rect 668584 671100 668636 671152
rect 674012 671100 674064 671152
rect 661684 670692 661736 670744
rect 673644 670692 673696 670744
rect 671804 670080 671856 670132
rect 674012 670080 674064 670132
rect 658924 669468 658976 669520
rect 673644 669468 673696 669520
rect 45376 669332 45428 669384
rect 53104 669332 53156 669384
rect 670424 669332 670476 669384
rect 674012 669332 674064 669384
rect 670976 669196 671028 669248
rect 671804 669196 671856 669248
rect 671344 668516 671396 668568
rect 674012 668516 674064 668568
rect 671620 668176 671672 668228
rect 673644 668176 673696 668228
rect 45744 667904 45796 667956
rect 57244 667904 57296 667956
rect 671344 667904 671396 667956
rect 674012 667904 674064 667956
rect 42248 667428 42300 667480
rect 45376 667428 45428 667480
rect 671988 666884 672040 666936
rect 674012 666884 674064 666936
rect 670976 666544 671028 666596
rect 673644 666544 673696 666596
rect 669780 665592 669832 665644
rect 674012 665592 674064 665644
rect 671804 665252 671856 665304
rect 673644 665252 673696 665304
rect 672356 665116 672408 665168
rect 673368 665116 673420 665168
rect 42248 664844 42300 664896
rect 43996 664844 44048 664896
rect 42248 664164 42300 664216
rect 42708 664164 42760 664216
rect 42248 663008 42300 663060
rect 43628 663008 43680 663060
rect 668768 662940 668820 662992
rect 674012 662940 674064 662992
rect 669596 662532 669648 662584
rect 674012 662532 674064 662584
rect 669044 661580 669096 661632
rect 674012 661580 674064 661632
rect 667848 661104 667900 661156
rect 674012 661104 674064 661156
rect 53104 660900 53156 660952
rect 62120 660900 62172 660952
rect 671160 660084 671212 660136
rect 674012 660084 674064 660136
rect 675852 659812 675904 659864
rect 683120 659812 683172 659864
rect 57244 659540 57296 659592
rect 62120 659540 62172 659592
rect 42524 657500 42576 657552
rect 62120 657500 62172 657552
rect 42064 657364 42116 657416
rect 42708 657364 42760 657416
rect 653404 655528 653456 655580
rect 674012 655528 674064 655580
rect 44824 655460 44876 655512
rect 62120 655460 62172 655512
rect 668216 654100 668268 654152
rect 674012 654100 674064 654152
rect 667388 647232 667440 647284
rect 674012 647232 674064 647284
rect 655520 645872 655572 645924
rect 671160 645872 671212 645924
rect 674932 645192 674984 645244
rect 675300 645192 675352 645244
rect 652024 645124 652076 645176
rect 668584 645124 668636 645176
rect 35808 644444 35860 644496
rect 41696 644444 41748 644496
rect 42064 644444 42116 644496
rect 60004 644444 60056 644496
rect 674564 643628 674616 643680
rect 35808 643492 35860 643544
rect 39948 643492 40000 643544
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 44640 643288 44692 643340
rect 674564 643288 674616 643340
rect 675116 643220 675168 643272
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 61384 643084 61436 643136
rect 655336 643084 655388 643136
rect 674012 643084 674064 643136
rect 674472 643084 674524 643136
rect 38568 642472 38620 642524
rect 41696 642472 41748 642524
rect 42064 642336 42116 642388
rect 62764 642336 62816 642388
rect 651472 642336 651524 642388
rect 658924 642336 658976 642388
rect 35624 641996 35676 642048
rect 40132 641996 40184 642048
rect 35808 641724 35860 641776
rect 41696 641724 41748 641776
rect 42064 641724 42116 641776
rect 45192 641724 45244 641776
rect 35808 640704 35860 640756
rect 39764 640704 39816 640756
rect 35440 640432 35492 640484
rect 40040 640432 40092 640484
rect 35624 640296 35676 640348
rect 41696 640296 41748 640348
rect 42064 640296 42116 640348
rect 45284 640296 45336 640348
rect 651472 640296 651524 640348
rect 669964 640296 670016 640348
rect 651380 640092 651432 640144
rect 653404 640092 653456 640144
rect 35808 639140 35860 639192
rect 37924 639072 37976 639124
rect 35808 638936 35860 638988
rect 41420 638868 41472 638920
rect 651656 638868 651708 638920
rect 655336 638868 655388 638920
rect 651472 638732 651524 638784
rect 655520 638732 655572 638784
rect 35808 637712 35860 637764
rect 36544 637712 36596 637764
rect 674564 636964 674616 637016
rect 675484 636964 675536 637016
rect 35624 636896 35676 636948
rect 40684 636896 40736 636948
rect 675852 636828 675904 636880
rect 683396 636828 683448 636880
rect 35532 636488 35584 636540
rect 39856 636420 39908 636472
rect 35808 636216 35860 636268
rect 41696 636216 41748 636268
rect 42064 636216 42116 636268
rect 44548 636216 44600 636268
rect 35808 634924 35860 634976
rect 41604 634924 41656 634976
rect 35808 633700 35860 633752
rect 39580 633632 39632 633684
rect 35624 633428 35676 633480
rect 40132 633428 40184 633480
rect 674932 631796 674984 631848
rect 675484 631796 675536 631848
rect 36544 630708 36596 630760
rect 41604 630708 41656 630760
rect 31944 629892 31996 629944
rect 40224 629892 40276 629944
rect 38568 628260 38620 628312
rect 40500 628260 40552 628312
rect 44180 625812 44232 625864
rect 62948 625812 63000 625864
rect 667204 625812 667256 625864
rect 674012 625812 674064 625864
rect 668584 625540 668636 625592
rect 674012 625540 674064 625592
rect 42248 625336 42300 625388
rect 42524 625336 42576 625388
rect 660304 625132 660356 625184
rect 673460 625200 673512 625252
rect 42524 625064 42576 625116
rect 42708 625064 42760 625116
rect 670424 625064 670476 625116
rect 674012 625064 674064 625116
rect 671160 624656 671212 624708
rect 674012 624656 674064 624708
rect 42340 624384 42392 624436
rect 44180 624384 44232 624436
rect 671620 624316 671672 624368
rect 674012 624316 674064 624368
rect 42248 624044 42300 624096
rect 44456 624044 44508 624096
rect 671620 623840 671672 623892
rect 674012 623840 674064 623892
rect 671344 623500 671396 623552
rect 674012 623500 674064 623552
rect 669596 623024 669648 623076
rect 674012 623024 674064 623076
rect 675852 623024 675904 623076
rect 683120 623024 683172 623076
rect 670976 622684 671028 622736
rect 674012 622684 674064 622736
rect 669780 622208 669832 622260
rect 674012 622208 674064 622260
rect 669412 621188 669464 621240
rect 674012 621188 674064 621240
rect 672172 620576 672224 620628
rect 673092 620576 673144 620628
rect 670240 619828 670292 619880
rect 673092 619828 673144 619880
rect 42248 619624 42300 619676
rect 44364 619624 44416 619676
rect 666468 619624 666520 619676
rect 673460 619624 673512 619676
rect 669228 619012 669280 619064
rect 673460 619012 673512 619064
rect 44180 616768 44232 616820
rect 62120 616768 62172 616820
rect 670792 616564 670844 616616
rect 673460 616564 673512 616616
rect 675852 615476 675904 615528
rect 683120 615476 683172 615528
rect 43076 615408 43128 615460
rect 44088 615408 44140 615460
rect 669412 614864 669464 614916
rect 673460 614864 673512 614916
rect 42616 614116 42668 614168
rect 62120 614116 62172 614168
rect 60004 612620 60056 612672
rect 62120 612620 62172 612672
rect 43812 612552 43864 612604
rect 44088 612348 44140 612400
rect 43904 612212 43956 612264
rect 44456 612212 44508 612264
rect 43766 612144 43818 612196
rect 44088 612008 44140 612060
rect 43996 611736 44048 611788
rect 44088 611532 44140 611584
rect 44456 611396 44508 611448
rect 44211 611328 44263 611380
rect 653404 611328 653456 611380
rect 673460 611328 673512 611380
rect 44318 611124 44370 611176
rect 44916 611124 44968 611176
rect 35808 601672 35860 601724
rect 36544 601672 36596 601724
rect 657544 600448 657596 600500
rect 673460 600448 673512 600500
rect 654784 598952 654836 599004
rect 673460 598952 673512 599004
rect 651472 597524 651524 597576
rect 668584 597524 668636 597576
rect 42984 597388 43036 597440
rect 42984 596980 43036 597032
rect 651472 596164 651524 596216
rect 667204 596164 667256 596216
rect 39948 595756 40000 595808
rect 41696 595756 41748 595808
rect 651656 595416 651708 595468
rect 653404 595416 653456 595468
rect 651472 594872 651524 594924
rect 656164 594872 656216 594924
rect 651472 594668 651524 594720
rect 657544 594668 657596 594720
rect 38568 594260 38620 594312
rect 41604 594260 41656 594312
rect 651472 593036 651524 593088
rect 654784 593036 654836 593088
rect 36544 592900 36596 592952
rect 41696 592900 41748 592952
rect 675852 592832 675904 592884
rect 678244 592832 678296 592884
rect 675852 591404 675904 591456
rect 683396 591404 683448 591456
rect 675852 591268 675904 591320
rect 684224 591268 684276 591320
rect 675852 589228 675904 589280
rect 681004 589228 681056 589280
rect 35440 587256 35492 587308
rect 40684 587256 40736 587308
rect 33048 587120 33100 587172
rect 41512 587120 41564 587172
rect 33784 585896 33836 585948
rect 40132 585896 40184 585948
rect 31024 585760 31076 585812
rect 40592 585760 40644 585812
rect 652024 581000 652076 581052
rect 674012 581000 674064 581052
rect 669964 580252 670016 580304
rect 674012 580252 674064 580304
rect 671160 579980 671212 580032
rect 674012 579980 674064 580032
rect 658924 579640 658976 579692
rect 673644 579640 673696 579692
rect 671620 578756 671672 578808
rect 674012 578756 674064 578808
rect 670148 578348 670200 578400
rect 674012 578348 674064 578400
rect 669964 578212 670016 578264
rect 673460 578212 673512 578264
rect 42248 577804 42300 577856
rect 42708 577804 42760 577856
rect 669780 577396 669832 577448
rect 674012 577396 674064 577448
rect 669596 577124 669648 577176
rect 673644 577124 673696 577176
rect 670240 576988 670292 577040
rect 673414 576988 673466 577040
rect 671160 576852 671212 576904
rect 674012 576920 674064 576972
rect 671988 575900 672040 575952
rect 674012 575900 674064 575952
rect 44640 575424 44692 575476
rect 62120 575424 62172 575476
rect 668216 574404 668268 574456
rect 674012 574404 674064 574456
rect 668860 574132 668912 574184
rect 673644 574132 673696 574184
rect 45560 573996 45612 574048
rect 62120 573996 62172 574048
rect 42156 573452 42208 573504
rect 42616 573452 42668 573504
rect 671804 572840 671856 572892
rect 674012 572840 674064 572892
rect 667388 571684 667440 571736
rect 673644 571684 673696 571736
rect 669044 571412 669096 571464
rect 674012 571412 674064 571464
rect 681004 571276 681056 571328
rect 683120 571276 683172 571328
rect 42064 570936 42116 570988
rect 42616 570936 42668 570988
rect 653404 565836 653456 565888
rect 674012 565836 674064 565888
rect 672724 557812 672776 557864
rect 673276 557812 673328 557864
rect 673828 556588 673880 556640
rect 674012 556588 674064 556640
rect 672724 555432 672776 555484
rect 673276 555432 673328 555484
rect 674656 554888 674708 554940
rect 675116 554888 675168 554940
rect 657820 554752 657872 554804
rect 674012 554820 674064 554872
rect 655152 553392 655204 553444
rect 674012 553392 674064 553444
rect 651472 552644 651524 552696
rect 665824 552644 665876 552696
rect 651472 552032 651524 552084
rect 660304 552032 660356 552084
rect 40040 550944 40092 550996
rect 41696 550944 41748 550996
rect 668860 550604 668912 550656
rect 673460 550604 673512 550656
rect 651380 550332 651432 550384
rect 653404 550332 653456 550384
rect 651472 549040 651524 549092
rect 657820 549040 657872 549092
rect 673184 548904 673236 548956
rect 651472 548768 651524 548820
rect 655152 548768 655204 548820
rect 673000 548496 673052 548548
rect 31760 547408 31812 547460
rect 41696 547408 41748 547460
rect 674288 547408 674340 547460
rect 675484 547544 675536 547596
rect 675852 547544 675904 547596
rect 684224 547544 684276 547596
rect 676036 547408 676088 547460
rect 683396 547408 683448 547460
rect 674288 547136 674340 547188
rect 675484 547272 675536 547324
rect 675852 547272 675904 547324
rect 683212 547272 683264 547324
rect 674288 547000 674340 547052
rect 675484 547000 675536 547052
rect 34428 544348 34480 544400
rect 41328 544348 41380 544400
rect 42984 538160 43036 538212
rect 42800 537888 42852 537940
rect 668584 535644 668636 535696
rect 674012 535644 674064 535696
rect 667204 535440 667256 535492
rect 673828 535440 673880 535492
rect 669964 534488 670016 534540
rect 674012 534488 674064 534540
rect 670148 534352 670200 534404
rect 674012 534352 674064 534404
rect 656164 534216 656216 534268
rect 673460 534216 673512 534268
rect 670792 534080 670844 534132
rect 673828 534080 673880 534132
rect 671620 533536 671672 533588
rect 674012 533536 674064 533588
rect 670240 533332 670292 533384
rect 674012 533332 674064 533384
rect 675852 533332 675904 533384
rect 683580 533332 683632 533384
rect 42432 532720 42484 532772
rect 43168 532720 43220 532772
rect 671804 532720 671856 532772
rect 674012 532720 674064 532772
rect 671160 532516 671212 532568
rect 674012 532516 674064 532568
rect 672448 531904 672500 531956
rect 674012 531904 674064 531956
rect 672632 531700 672684 531752
rect 674012 531700 674064 531752
rect 60004 531224 60056 531276
rect 62120 531224 62172 531276
rect 44732 531088 44784 531140
rect 62120 531088 62172 531140
rect 672724 530204 672776 530256
rect 673460 530204 673512 530256
rect 42156 530068 42208 530120
rect 42984 530068 43036 530120
rect 670424 530068 670476 530120
rect 673828 530068 673880 530120
rect 667572 529932 667624 529984
rect 674012 529932 674064 529984
rect 670976 529660 671028 529712
rect 674012 529660 674064 529712
rect 45100 528572 45152 528624
rect 62120 528572 62172 528624
rect 669228 528572 669280 528624
rect 674012 528572 674064 528624
rect 672264 528436 672316 528488
rect 674012 528436 674064 528488
rect 42064 527756 42116 527808
rect 42616 527756 42668 527808
rect 672724 526464 672776 526516
rect 673276 526464 673328 526516
rect 671344 524628 671396 524680
rect 674012 524628 674064 524680
rect 675852 524560 675904 524612
rect 683120 524560 683172 524612
rect 675852 518848 675904 518900
rect 677692 518848 677744 518900
rect 677876 518780 677928 518832
rect 676036 518644 676088 518696
rect 675300 503888 675352 503940
rect 675484 503888 675536 503940
rect 676128 503752 676180 503804
rect 678244 503752 678296 503804
rect 675300 503616 675352 503668
rect 675484 503616 675536 503668
rect 677416 503616 677468 503668
rect 683396 503616 683448 503668
rect 675852 500760 675904 500812
rect 681004 500760 681056 500812
rect 652024 493280 652076 493332
rect 672908 493280 672960 493332
rect 665824 491444 665876 491496
rect 674012 491444 674064 491496
rect 660304 491308 660356 491360
rect 673828 491308 673880 491360
rect 670792 490900 670844 490952
rect 674012 490900 674064 490952
rect 671620 490084 671672 490136
rect 674012 490084 674064 490136
rect 676036 490016 676088 490068
rect 676588 490016 676640 490068
rect 672632 489608 672684 489660
rect 674012 489608 674064 489660
rect 671804 489268 671856 489320
rect 674012 489268 674064 489320
rect 672448 488452 672500 488504
rect 674012 488452 674064 488504
rect 676220 487160 676272 487212
rect 677508 487160 677560 487212
rect 668400 485800 668452 485852
rect 674012 485800 674064 485852
rect 669044 484508 669096 484560
rect 674012 484508 674064 484560
rect 668860 484372 668912 484424
rect 673828 484372 673880 484424
rect 671988 482332 672040 482384
rect 674012 482332 674064 482384
rect 676128 480360 676180 480412
rect 683120 480360 683172 480412
rect 670608 456356 670660 456408
rect 676220 456152 676272 456204
rect 676174 455948 676226 456000
rect 673276 455812 673328 455864
rect 673828 455812 673880 455864
rect 667848 455608 667900 455660
rect 673276 455336 673328 455388
rect 673388 455200 673440 455252
rect 673276 454996 673328 455048
rect 672080 454792 672132 454844
rect 673046 454588 673098 454640
rect 672954 454316 673006 454368
rect 674288 454316 674340 454368
rect 675484 454316 675536 454368
rect 672816 454044 672868 454096
rect 672448 453908 672500 453960
rect 35808 429156 35860 429208
rect 41696 429156 41748 429208
rect 41328 425076 41380 425128
rect 41696 425076 41748 425128
rect 40960 424260 41012 424312
rect 41512 424260 41564 424312
rect 32036 416168 32088 416220
rect 41696 416168 41748 416220
rect 53840 404268 53892 404320
rect 62120 404268 62172 404320
rect 44824 402908 44876 402960
rect 62120 402908 62172 402960
rect 51080 400188 51132 400240
rect 62120 400188 62172 400240
rect 60004 400052 60056 400104
rect 62120 400052 62172 400104
rect 674840 385568 674892 385620
rect 675300 385568 675352 385620
rect 41328 382236 41380 382288
rect 41696 382236 41748 382288
rect 674472 382168 674524 382220
rect 675392 382168 675444 382220
rect 35808 379652 35860 379704
rect 40592 379652 40644 379704
rect 674380 378088 674432 378140
rect 675116 378088 675168 378140
rect 40224 378020 40276 378072
rect 41696 378020 41748 378072
rect 42064 377952 42116 378004
rect 42708 377952 42760 378004
rect 651472 373940 651524 373992
rect 657544 373940 657596 373992
rect 35164 371832 35216 371884
rect 41696 371832 41748 371884
rect 651472 370948 651524 371000
rect 654784 370948 654836 371000
rect 42248 365236 42300 365288
rect 42248 364896 42300 364948
rect 42248 364284 42300 364336
rect 42708 364148 42760 364200
rect 46572 361496 46624 361548
rect 62120 361496 62172 361548
rect 45376 360136 45428 360188
rect 62120 360136 62172 360188
rect 44640 359592 44692 359644
rect 45376 359592 45428 359644
rect 44824 359456 44876 359508
rect 45468 359456 45520 359508
rect 51724 357416 51776 357468
rect 62120 357416 62172 357468
rect 44640 354696 44692 354748
rect 44824 354696 44876 354748
rect 44732 354424 44784 354476
rect 44855 354424 44907 354476
rect 45836 353880 45888 353932
rect 45836 353676 45888 353728
rect 45303 353472 45355 353524
rect 45422 353200 45474 353252
rect 676036 347420 676088 347472
rect 676496 347420 676548 347472
rect 35808 344564 35860 344616
rect 39856 344564 39908 344616
rect 35624 343612 35676 343664
rect 40040 343612 40092 343664
rect 35808 342184 35860 342236
rect 40224 342184 40276 342236
rect 45468 342184 45520 342236
rect 63132 342184 63184 342236
rect 35808 341504 35860 341556
rect 40224 341504 40276 341556
rect 35808 341028 35860 341080
rect 40132 341028 40184 341080
rect 35532 339600 35584 339652
rect 37096 339600 37148 339652
rect 35808 339464 35860 339516
rect 38844 339464 38896 339516
rect 674840 339328 674892 339380
rect 675484 339328 675536 339380
rect 674380 336540 674432 336592
rect 675392 336540 675444 336592
rect 35808 335316 35860 335368
rect 39856 335316 39908 335368
rect 35808 334092 35860 334144
rect 40316 334092 40368 334144
rect 651380 328244 651432 328296
rect 654784 328244 654836 328296
rect 651380 325592 651432 325644
rect 653404 325592 653456 325644
rect 53840 317364 53892 317416
rect 62120 317364 62172 317416
rect 53104 315936 53156 315988
rect 62120 315936 62172 315988
rect 59912 314712 59964 314764
rect 62120 314712 62172 314764
rect 676220 307776 676272 307828
rect 676864 307776 676916 307828
rect 675852 304104 675904 304156
rect 676220 304104 676272 304156
rect 651380 303492 651432 303544
rect 653404 303492 653456 303544
rect 651472 300772 651524 300824
rect 664444 300772 664496 300824
rect 35624 298732 35676 298784
rect 41604 298732 41656 298784
rect 35808 298256 35860 298308
rect 41604 298256 41656 298308
rect 651472 298120 651524 298172
rect 662420 298120 662472 298172
rect 675852 298052 675904 298104
rect 676864 298052 676916 298104
rect 676128 297916 676180 297968
rect 679624 297916 679676 297968
rect 675944 297440 675996 297492
rect 677600 297440 677652 297492
rect 651472 297032 651524 297084
rect 656164 297032 656216 297084
rect 675484 296352 675536 296404
rect 652668 295944 652720 295996
rect 665824 295944 665876 295996
rect 675484 295740 675536 295792
rect 35808 295604 35860 295656
rect 40684 295604 40736 295656
rect 35440 295468 35492 295520
rect 41328 295468 41380 295520
rect 58624 295400 58676 295452
rect 62120 295400 62172 295452
rect 35624 295332 35676 295384
rect 41604 295332 41656 295384
rect 35808 294108 35860 294160
rect 41696 294108 41748 294160
rect 57244 294040 57296 294092
rect 62120 294040 62172 294092
rect 651472 293972 651524 294024
rect 664444 293972 664496 294024
rect 35808 292884 35860 292936
rect 41512 292816 41564 292868
rect 35808 292544 35860 292596
rect 54484 292544 54536 292596
rect 62304 292544 62356 292596
rect 651472 292544 651524 292596
rect 663064 292544 663116 292596
rect 42064 292408 42116 292460
rect 42984 292408 43036 292460
rect 46204 292408 46256 292460
rect 62120 292408 62172 292460
rect 41604 292204 41656 292256
rect 53104 291116 53156 291168
rect 62120 291116 62172 291168
rect 35808 289892 35860 289944
rect 41696 290096 41748 290148
rect 651472 289824 651524 289876
rect 660304 289824 660356 289876
rect 35624 289076 35676 289128
rect 41696 289008 41748 289060
rect 55864 288464 55916 288516
rect 62120 288464 62172 288516
rect 651472 288396 651524 288448
rect 661684 288396 661736 288448
rect 651472 287036 651524 287088
rect 672264 287036 672316 287088
rect 674380 286968 674432 287020
rect 675116 286968 675168 287020
rect 33784 286288 33836 286340
rect 41696 286288 41748 286340
rect 46204 285676 46256 285728
rect 62120 285676 62172 285728
rect 651472 285676 651524 285728
rect 668124 285676 668176 285728
rect 60004 284384 60056 284436
rect 62120 284384 62172 284436
rect 651472 284316 651524 284368
rect 672080 284316 672132 284368
rect 47768 280304 47820 280356
rect 62120 280304 62172 280356
rect 651472 280304 651524 280356
rect 667204 280304 667256 280356
rect 651656 280168 651708 280220
rect 667388 280168 667440 280220
rect 42248 280100 42300 280152
rect 42984 280100 43036 280152
rect 482836 277312 482888 277364
rect 557540 277312 557592 277364
rect 485688 277176 485740 277228
rect 562324 277176 562376 277228
rect 495072 277040 495124 277092
rect 576492 277040 576544 277092
rect 511632 276904 511684 276956
rect 600136 276904 600188 276956
rect 514484 276768 514536 276820
rect 603632 276768 603684 276820
rect 518716 276632 518768 276684
rect 609612 276632 609664 276684
rect 477040 276496 477092 276548
rect 550456 276496 550508 276548
rect 478512 276360 478564 276412
rect 551652 276360 551704 276412
rect 471612 276224 471664 276276
rect 543372 276224 543424 276276
rect 543372 276088 543424 276140
rect 549260 276088 549312 276140
rect 107200 275952 107252 276004
rect 162124 275952 162176 276004
rect 185216 275952 185268 276004
rect 221280 275952 221332 276004
rect 454408 275952 454460 276004
rect 100116 275816 100168 275868
rect 161388 275816 161440 275868
rect 161572 275816 161624 275868
rect 161756 275816 161808 275868
rect 167000 275816 167052 275868
rect 178132 275816 178184 275868
rect 216680 275816 216732 275868
rect 217140 275816 217192 275868
rect 224040 275816 224092 275868
rect 232504 275816 232556 275868
rect 239864 275816 239916 275868
rect 284576 275816 284628 275868
rect 290096 275816 290148 275868
rect 445024 275816 445076 275868
rect 457444 275952 457496 276004
rect 509056 275952 509108 276004
rect 517152 275952 517204 276004
rect 608416 275952 608468 276004
rect 93032 275680 93084 275732
rect 155960 275680 156012 275732
rect 163136 275680 163188 275732
rect 164056 275680 164108 275732
rect 76472 275544 76524 275596
rect 86224 275544 86276 275596
rect 90732 275544 90784 275596
rect 154764 275544 154816 275596
rect 156880 275544 156932 275596
rect 171048 275680 171100 275732
rect 211068 275680 211120 275732
rect 224224 275680 224276 275732
rect 232780 275680 232832 275732
rect 236092 275680 236144 275732
rect 253388 275680 253440 275732
rect 435640 275680 435692 275732
rect 454408 275680 454460 275732
rect 475384 275816 475436 275868
rect 479524 275816 479576 275868
rect 523316 275816 523368 275868
rect 524144 275816 524196 275868
rect 615500 275816 615552 275868
rect 498476 275680 498528 275732
rect 507860 275680 507912 275732
rect 545764 275680 545816 275732
rect 277492 275612 277544 275664
rect 284300 275612 284352 275664
rect 291660 275612 291712 275664
rect 295340 275612 295392 275664
rect 81256 275408 81308 275460
rect 145564 275408 145616 275460
rect 160468 275408 160520 275460
rect 161848 275408 161900 275460
rect 206376 275544 206428 275596
rect 221924 275544 221976 275596
rect 239404 275544 239456 275596
rect 243176 275544 243228 275596
rect 255320 275544 255372 275596
rect 257344 275544 257396 275596
rect 262864 275544 262916 275596
rect 286876 275544 286928 275596
rect 430212 275544 430264 275596
rect 484308 275544 484360 275596
rect 501604 275544 501656 275596
rect 512644 275544 512696 275596
rect 515404 275544 515456 275596
rect 526812 275544 526864 275596
rect 528192 275544 528244 275596
rect 622584 275544 622636 275596
rect 291752 275476 291804 275528
rect 198740 275408 198792 275460
rect 214840 275408 214892 275460
rect 236644 275408 236696 275460
rect 239588 275408 239640 275460
rect 251916 275408 251968 275460
rect 263232 275408 263284 275460
rect 273260 275408 273312 275460
rect 285680 275408 285732 275460
rect 291200 275408 291252 275460
rect 386052 275408 386104 275460
rect 420460 275408 420512 275460
rect 423404 275408 423456 275460
rect 473360 275408 473412 275460
rect 475384 275408 475436 275460
rect 485044 275408 485096 275460
rect 485228 275408 485280 275460
rect 537484 275408 537536 275460
rect 299940 275340 299992 275392
rect 301228 275340 301280 275392
rect 71780 275272 71832 275324
rect 141056 275272 141108 275324
rect 146208 275272 146260 275324
rect 189080 275272 189132 275324
rect 218336 275272 218388 275324
rect 243084 275272 243136 275324
rect 256148 275272 256200 275324
rect 268844 275272 268896 275324
rect 273904 275272 273956 275324
rect 282920 275272 282972 275324
rect 290464 275272 290516 275324
rect 294144 275272 294196 275324
rect 361212 275272 361264 275324
rect 385040 275272 385092 275324
rect 416412 275272 416464 275324
rect 462964 275272 463016 275324
rect 463148 275272 463200 275324
rect 530400 275272 530452 275324
rect 532332 275272 532384 275324
rect 537300 275272 537352 275324
rect 537576 275272 537628 275324
rect 636752 275408 636804 275460
rect 537944 275272 537996 275324
rect 540980 275272 541032 275324
rect 543004 275272 543056 275324
rect 629668 275272 629720 275324
rect 298744 275204 298796 275256
rect 300032 275204 300084 275256
rect 139124 275136 139176 275188
rect 146944 275136 146996 275188
rect 149796 275136 149848 275188
rect 191748 275136 191800 275188
rect 292856 275136 292908 275188
rect 295800 275136 295852 275188
rect 427084 275136 427136 275188
rect 477224 275136 477276 275188
rect 485044 275136 485096 275188
rect 491392 275136 491444 275188
rect 493324 275136 493376 275188
rect 269212 275068 269264 275120
rect 274916 275068 274968 275120
rect 110788 275000 110840 275052
rect 149704 275000 149756 275052
rect 153384 275000 153436 275052
rect 154488 275000 154540 275052
rect 132040 274864 132092 274916
rect 161664 275000 161716 275052
rect 161848 275000 161900 275052
rect 175924 275000 175976 275052
rect 190000 275000 190052 275052
rect 218704 275000 218756 275052
rect 288072 275000 288124 275052
rect 292672 275000 292724 275052
rect 420644 275000 420696 275052
rect 470140 275000 470192 275052
rect 476120 275000 476172 275052
rect 485228 275000 485280 275052
rect 492404 275000 492456 275052
rect 494888 275000 494940 275052
rect 497464 275136 497516 275188
rect 505560 275136 505612 275188
rect 507492 275136 507544 275188
rect 594248 275136 594300 275188
rect 501972 275000 502024 275052
rect 503444 275000 503496 275052
rect 587072 275000 587124 275052
rect 293960 274932 294012 274984
rect 297180 274932 297232 274984
rect 167552 274864 167604 274916
rect 169024 274864 169076 274916
rect 413468 274864 413520 274916
rect 459468 274864 459520 274916
rect 473360 274864 473412 274916
rect 544568 274864 544620 274916
rect 174636 274796 174688 274848
rect 182732 274796 182784 274848
rect 289268 274796 289320 274848
rect 293408 274796 293460 274848
rect 296352 274796 296404 274848
rect 298376 274796 298428 274848
rect 136824 274728 136876 274780
rect 137652 274728 137704 274780
rect 143908 274728 143960 274780
rect 144368 274728 144420 274780
rect 146944 274728 146996 274780
rect 174452 274728 174504 274780
rect 469864 274728 469916 274780
rect 516232 274728 516284 274780
rect 526444 274728 526496 274780
rect 533896 274728 533948 274780
rect 534724 274728 534776 274780
rect 537944 274728 537996 274780
rect 538128 274728 538180 274780
rect 543004 274728 543056 274780
rect 543188 274728 543240 274780
rect 643836 274728 643888 274780
rect 74172 274660 74224 274712
rect 76748 274660 76800 274712
rect 85948 274660 86000 274712
rect 90364 274660 90416 274712
rect 103704 274660 103756 274712
rect 104808 274660 104860 274712
rect 253848 274660 253900 274712
rect 258356 274660 258408 274712
rect 268016 274660 268068 274712
rect 272432 274660 272484 274712
rect 283380 274660 283432 274712
rect 289176 274660 289228 274712
rect 295156 274660 295208 274712
rect 296812 274660 296864 274712
rect 297548 274660 297600 274712
rect 299572 274660 299624 274712
rect 303436 274660 303488 274712
rect 303988 274660 304040 274712
rect 321192 274660 321244 274712
rect 328276 274660 328328 274712
rect 350724 274660 350776 274712
rect 353116 274660 353168 274712
rect 113456 274592 113508 274644
rect 169944 274592 169996 274644
rect 182916 274592 182968 274644
rect 214564 274592 214616 274644
rect 382924 274592 382976 274644
rect 392124 274592 392176 274644
rect 404176 274592 404228 274644
rect 446496 274592 446548 274644
rect 450544 274592 450596 274644
rect 480720 274592 480772 274644
rect 488356 274592 488408 274644
rect 567016 274592 567068 274644
rect 67088 274320 67140 274372
rect 95884 274456 95936 274508
rect 105176 274456 105228 274508
rect 163320 274456 163372 274508
rect 168748 274456 168800 274508
rect 208492 274456 208544 274508
rect 227812 274456 227864 274508
rect 248880 274456 248932 274508
rect 358084 274456 358136 274508
rect 369584 274456 369636 274508
rect 95424 274320 95476 274372
rect 157616 274320 157668 274372
rect 166356 274320 166408 274372
rect 207296 274320 207348 274372
rect 207756 274320 207808 274372
rect 233884 274320 233936 274372
rect 249064 274320 249116 274372
rect 265256 274320 265308 274372
rect 333796 274320 333848 274372
rect 345940 274320 345992 274372
rect 347044 274320 347096 274372
rect 359004 274320 359056 274372
rect 369124 274320 369176 274372
rect 395620 274456 395672 274508
rect 409236 274456 409288 274508
rect 453580 274456 453632 274508
rect 453764 274456 453816 274508
rect 486608 274456 486660 274508
rect 536748 274456 536800 274508
rect 543694 274456 543746 274508
rect 543832 274456 543884 274508
rect 639144 274456 639196 274508
rect 373264 274320 373316 274372
rect 400312 274320 400364 274372
rect 413836 274320 413888 274372
rect 460664 274320 460716 274372
rect 465724 274320 465776 274372
rect 487804 274320 487856 274372
rect 508596 274320 508648 274372
rect 595076 274320 595128 274372
rect 595444 274320 595496 274372
rect 640340 274320 640392 274372
rect 282184 274252 282236 274304
rect 287704 274252 287756 274304
rect 89444 274184 89496 274236
rect 152004 274184 152056 274236
rect 155684 274184 155736 274236
rect 200120 274184 200172 274236
rect 205364 274184 205416 274236
rect 234712 274184 234764 274236
rect 234896 274184 234948 274236
rect 77668 274048 77720 274100
rect 144920 274048 144972 274100
rect 147404 274048 147456 274100
rect 193404 274048 193456 274100
rect 198280 274048 198332 274100
rect 229192 274048 229244 274100
rect 237288 274048 237340 274100
rect 255320 274184 255372 274236
rect 261024 274184 261076 274236
rect 325332 274184 325384 274236
rect 332968 274184 333020 274236
rect 343456 274184 343508 274236
rect 360200 274184 360252 274236
rect 364984 274184 365036 274236
rect 374368 274184 374420 274236
rect 379336 274184 379388 274236
rect 410984 274184 411036 274236
rect 416596 274184 416648 274236
rect 464160 274184 464212 274236
rect 474648 274184 474700 274236
rect 507860 274184 507912 274236
rect 511816 274184 511868 274236
rect 598940 274184 598992 274236
rect 65892 273912 65944 273964
rect 136824 273912 136876 273964
rect 145104 273912 145156 273964
rect 192392 273912 192444 273964
rect 195888 273912 195940 273964
rect 227904 273912 227956 273964
rect 229008 273912 229060 273964
rect 250444 273912 250496 273964
rect 255412 274048 255464 274100
rect 261208 274048 261260 274100
rect 273536 274048 273588 274100
rect 275100 274048 275152 274100
rect 283472 274048 283524 274100
rect 332324 274048 332376 274100
rect 343640 274048 343692 274100
rect 350356 274048 350408 274100
rect 368480 274048 368532 274100
rect 369308 274048 369360 274100
rect 387340 274048 387392 274100
rect 394332 274048 394384 274100
rect 432236 274048 432288 274100
rect 432604 274048 432656 274100
rect 485504 274048 485556 274100
rect 491208 274048 491260 274100
rect 569960 274048 570012 274100
rect 571800 274048 571852 274100
rect 583576 274048 583628 274100
rect 256976 273912 257028 273964
rect 258540 273912 258592 273964
rect 272064 273912 272116 273964
rect 272708 273912 272760 273964
rect 281816 273912 281868 273964
rect 324044 273912 324096 273964
rect 331772 273912 331824 273964
rect 331956 273912 332008 273964
rect 341248 273912 341300 273964
rect 342076 273912 342128 273964
rect 357808 273912 357860 273964
rect 360108 273912 360160 273964
rect 382648 273912 382700 273964
rect 387432 273912 387484 273964
rect 421656 273912 421708 273964
rect 421840 273912 421892 273964
rect 471244 273912 471296 273964
rect 475752 273912 475804 273964
rect 543372 273912 543424 273964
rect 543832 273912 543884 273964
rect 634360 273912 634412 273964
rect 96620 273776 96672 273828
rect 117964 273776 118016 273828
rect 118240 273776 118292 273828
rect 174176 273776 174228 273828
rect 175924 273776 175976 273828
rect 204260 273776 204312 273828
rect 206560 273776 206612 273828
rect 235448 273776 235500 273828
rect 400036 273776 400088 273828
rect 439320 273776 439372 273828
rect 442264 273776 442316 273828
rect 481916 273776 481968 273828
rect 487068 273776 487120 273828
rect 560300 273776 560352 273828
rect 123760 273640 123812 273692
rect 177488 273640 177540 273692
rect 392584 273640 392636 273692
rect 409788 273640 409840 273692
rect 440884 273640 440936 273692
rect 474832 273640 474884 273692
rect 481364 273640 481416 273692
rect 556344 273640 556396 273692
rect 571800 273776 571852 273828
rect 571984 273776 572036 273828
rect 597744 273776 597796 273828
rect 134432 273504 134484 273556
rect 185124 273504 185176 273556
rect 446404 273504 446456 273556
rect 475936 273504 475988 273556
rect 484308 273504 484360 273556
rect 549904 273504 549956 273556
rect 556804 273504 556856 273556
rect 590660 273640 590712 273692
rect 563704 273504 563756 273556
rect 571984 273504 572036 273556
rect 135628 273368 135680 273420
rect 146944 273368 146996 273420
rect 460020 273368 460072 273420
rect 465724 273368 465776 273420
rect 467564 273368 467616 273420
rect 476120 273368 476172 273420
rect 478696 273368 478748 273420
rect 543694 273368 543746 273420
rect 559932 273368 559984 273420
rect 560300 273368 560352 273420
rect 563428 273368 563480 273420
rect 374644 273300 374696 273352
rect 377864 273300 377916 273352
rect 453304 273300 453356 273352
rect 453764 273300 453816 273352
rect 318616 273232 318668 273284
rect 324688 273232 324740 273284
rect 327540 273232 327592 273284
rect 329472 273232 329524 273284
rect 114376 273164 114428 273216
rect 171600 273164 171652 273216
rect 184112 273164 184164 273216
rect 218888 273164 218940 273216
rect 366364 273164 366416 273216
rect 383844 273164 383896 273216
rect 401508 273164 401560 273216
rect 442908 273164 442960 273216
rect 451188 273164 451240 273216
rect 513840 273164 513892 273216
rect 514024 273164 514076 273216
rect 519728 273164 519780 273216
rect 521476 273164 521528 273216
rect 614304 273164 614356 273216
rect 278596 273096 278648 273148
rect 285864 273096 285916 273148
rect 101312 273028 101364 273080
rect 160928 273028 160980 273080
rect 172244 273028 172296 273080
rect 210608 273028 210660 273080
rect 224040 273028 224092 273080
rect 243268 273028 243320 273080
rect 329472 273028 329524 273080
rect 338856 273028 338908 273080
rect 349804 273028 349856 273080
rect 366088 273028 366140 273080
rect 377404 273028 377456 273080
rect 399208 273028 399260 273080
rect 408224 273028 408276 273080
rect 450820 273028 450872 273080
rect 452292 273028 452344 273080
rect 99012 272892 99064 272944
rect 160100 272892 160152 272944
rect 162768 272892 162820 272944
rect 204720 272892 204772 272944
rect 219532 272892 219584 272944
rect 244464 272892 244516 272944
rect 252652 272892 252704 272944
rect 267924 272892 267976 272944
rect 335268 272892 335320 272944
rect 346860 272892 346912 272944
rect 362776 272892 362828 272944
rect 385868 272892 385920 272944
rect 406844 272892 406896 272944
rect 449992 272892 450044 272944
rect 455236 272892 455288 272944
rect 458088 273028 458140 273080
rect 465540 273028 465592 273080
rect 465724 273028 465776 273080
rect 518532 273028 518584 273080
rect 526812 273028 526864 273080
rect 621388 273028 621440 273080
rect 82452 272756 82504 272808
rect 148416 272756 148468 272808
rect 158076 272756 158128 272808
rect 200672 272756 200724 272808
rect 208860 272756 208912 272808
rect 237380 272756 237432 272808
rect 251456 272756 251508 272808
rect 267004 272756 267056 272808
rect 271512 272756 271564 272808
rect 280344 272756 280396 272808
rect 336372 272756 336424 272808
rect 349528 272756 349580 272808
rect 352564 272756 352616 272808
rect 370780 272756 370832 272808
rect 375196 272756 375248 272808
rect 403900 272756 403952 272808
rect 412272 272756 412324 272808
rect 457076 272756 457128 272808
rect 515036 272892 515088 272944
rect 529848 272892 529900 272944
rect 624976 272892 625028 272944
rect 465724 272756 465776 272808
rect 69388 272620 69440 272672
rect 139400 272620 139452 272672
rect 141516 272620 141568 272672
rect 184940 272620 184992 272672
rect 189080 272620 189132 272672
rect 194048 272620 194100 272672
rect 194692 272620 194744 272672
rect 227168 272620 227220 272672
rect 238484 272620 238536 272672
rect 258080 272620 258132 272672
rect 266820 272620 266872 272672
rect 277584 272620 277636 272672
rect 280988 272620 281040 272672
rect 286324 272620 286376 272672
rect 322756 272620 322808 272672
rect 330576 272620 330628 272672
rect 338028 272620 338080 272672
rect 351920 272620 351972 272672
rect 354496 272620 354548 272672
rect 375564 272620 375616 272672
rect 382004 272620 382056 272672
rect 414572 272620 414624 272672
rect 419172 272620 419224 272672
rect 465356 272620 465408 272672
rect 465540 272620 465592 272672
rect 522120 272756 522172 272808
rect 522764 272756 522816 272808
rect 524144 272756 524196 272808
rect 532516 272756 532568 272808
rect 628472 272756 628524 272808
rect 466092 272620 466144 272672
rect 467380 272620 467432 272672
rect 467748 272620 467800 272672
rect 470416 272620 470468 272672
rect 470600 272620 470652 272672
rect 536288 272620 536340 272672
rect 536564 272620 536616 272672
rect 635556 272620 635608 272672
rect 72976 272484 73028 272536
rect 142160 272484 142212 272536
rect 152188 272484 152240 272536
rect 197544 272484 197596 272536
rect 199476 272484 199528 272536
rect 230572 272484 230624 272536
rect 233700 272484 233752 272536
rect 253940 272484 253992 272536
rect 264428 272484 264480 272536
rect 276020 272484 276072 272536
rect 325516 272484 325568 272536
rect 334164 272484 334216 272536
rect 344652 272484 344704 272536
rect 361396 272484 361448 272536
rect 363788 272484 363840 272536
rect 388536 272484 388588 272536
rect 397276 272484 397328 272536
rect 435824 272484 435876 272536
rect 438768 272484 438820 272536
rect 489874 272484 489926 272536
rect 490012 272484 490064 272536
rect 529204 272484 529256 272536
rect 533712 272484 533764 272536
rect 632060 272484 632112 272536
rect 120264 272348 120316 272400
rect 175280 272348 175332 272400
rect 184940 272348 184992 272400
rect 189172 272348 189224 272400
rect 193588 272348 193640 272400
rect 224224 272348 224276 272400
rect 388996 272348 389048 272400
rect 425152 272348 425204 272400
rect 449808 272348 449860 272400
rect 511448 272348 511500 272400
rect 512644 272348 512696 272400
rect 514024 272348 514076 272400
rect 517336 272348 517388 272400
rect 607220 272348 607272 272400
rect 119068 272212 119120 272264
rect 172520 272212 172572 272264
rect 174452 272212 174504 272264
rect 189356 272212 189408 272264
rect 446956 272212 447008 272264
rect 508044 272212 508096 272264
rect 520096 272212 520148 272264
rect 610716 272212 610768 272264
rect 130844 272076 130896 272128
rect 182456 272076 182508 272128
rect 426348 272076 426400 272128
rect 470554 272076 470606 272128
rect 470784 272076 470836 272128
rect 489874 272076 489926 272128
rect 490012 272076 490064 272128
rect 558736 272076 558788 272128
rect 191472 271940 191524 271992
rect 108396 271804 108448 271856
rect 165896 271804 165948 271856
rect 188804 271804 188856 271856
rect 192576 271804 192628 271856
rect 447784 271940 447836 271992
rect 506756 271940 506808 271992
rect 507124 271940 507176 271992
rect 569408 271940 569460 271992
rect 268844 271872 268896 271924
rect 270500 271872 270552 271924
rect 225052 271804 225104 271856
rect 225420 271804 225472 271856
rect 228364 271804 228416 271856
rect 355324 271804 355376 271856
rect 356612 271804 356664 271856
rect 376576 271804 376628 271856
rect 407488 271804 407540 271856
rect 407764 271804 407816 271856
rect 437020 271804 437072 271856
rect 437204 271804 437256 271856
rect 493692 271804 493744 271856
rect 496544 271804 496596 271856
rect 578516 271804 578568 271856
rect 578884 271804 578936 271856
rect 611912 271804 611964 271856
rect 106096 271668 106148 271720
rect 164976 271668 165028 271720
rect 175740 271668 175792 271720
rect 213000 271668 213052 271720
rect 239864 271668 239916 271720
rect 254124 271668 254176 271720
rect 353944 271668 353996 271720
rect 372804 271668 372856 271720
rect 384948 271668 385000 271720
rect 418068 271668 418120 271720
rect 420184 271668 420236 271720
rect 431132 271668 431184 271720
rect 434628 271668 434680 271720
rect 485228 271668 485280 271720
rect 485412 271668 485464 271720
rect 490012 271668 490064 271720
rect 501972 271668 502024 271720
rect 585968 271668 586020 271720
rect 94228 271532 94280 271584
rect 156144 271532 156196 271584
rect 170128 271532 170180 271584
rect 209780 271532 209832 271584
rect 223120 271532 223172 271584
rect 247224 271532 247276 271584
rect 357164 271532 357216 271584
rect 379060 271532 379112 271584
rect 387616 271532 387668 271584
rect 422852 271532 422904 271584
rect 439964 271532 440016 271584
rect 497280 271532 497332 271584
rect 499304 271532 499356 271584
rect 582380 271532 582432 271584
rect 585784 271532 585836 271584
rect 626080 271532 626132 271584
rect 87144 271396 87196 271448
rect 152188 271396 152240 271448
rect 159272 271396 159324 271448
rect 202328 271396 202380 271448
rect 213644 271396 213696 271448
rect 240416 271396 240468 271448
rect 250260 271396 250312 271448
rect 75368 271260 75420 271312
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 142712 271260 142764 271312
rect 144184 271260 144236 271312
rect 154304 271260 154356 271312
rect 198096 271260 198148 271312
rect 212264 271260 212316 271312
rect 239312 271260 239364 271312
rect 244648 271260 244700 271312
rect 262220 271260 262272 271312
rect 265624 271396 265676 271448
rect 276848 271396 276900 271448
rect 339224 271396 339276 271448
rect 354220 271396 354272 271448
rect 358728 271396 358780 271448
rect 381452 271396 381504 271448
rect 393964 271396 394016 271448
rect 429936 271396 429988 271448
rect 442908 271396 442960 271448
rect 500868 271396 500920 271448
rect 505008 271396 505060 271448
rect 589464 271396 589516 271448
rect 266452 271260 266504 271312
rect 276664 271260 276716 271312
rect 284484 271260 284536 271312
rect 329656 271260 329708 271312
rect 340052 271260 340104 271312
rect 340604 271260 340656 271312
rect 355140 271260 355192 271312
rect 365444 271260 365496 271312
rect 390928 271260 390980 271312
rect 391848 271260 391900 271312
rect 428740 271260 428792 271312
rect 445668 271260 445720 271312
rect 504364 271260 504416 271312
rect 507676 271260 507728 271312
rect 593052 271260 593104 271312
rect 612004 271260 612056 271312
rect 618628 271260 618680 271312
rect 618904 271260 618956 271312
rect 633256 271260 633308 271312
rect 142712 271124 142764 271176
rect 148600 271124 148652 271176
rect 194784 271124 194836 271176
rect 197084 271124 197136 271176
rect 229284 271124 229336 271176
rect 230204 271124 230256 271176
rect 251732 271124 251784 271176
rect 254952 271124 255004 271176
rect 269304 271124 269356 271176
rect 270316 271124 270368 271176
rect 280528 271124 280580 271176
rect 331128 271124 331180 271176
rect 342444 271124 342496 271176
rect 347596 271124 347648 271176
rect 364524 271124 364576 271176
rect 366916 271124 366968 271176
rect 393320 271124 393372 271176
rect 402612 271124 402664 271176
rect 444104 271124 444156 271176
rect 459468 271124 459520 271176
rect 523868 271124 523920 271176
rect 524052 271124 524104 271176
rect 617800 271124 617852 271176
rect 625804 271124 625856 271176
rect 645032 271124 645084 271176
rect 116676 270988 116728 271040
rect 172704 270988 172756 271040
rect 192760 270988 192812 271040
rect 225512 270988 225564 271040
rect 326436 270988 326488 271040
rect 335084 270988 335136 271040
rect 381544 270988 381596 271040
rect 411812 270988 411864 271040
rect 414480 270988 414532 271040
rect 438124 270988 438176 271040
rect 438308 270988 438360 271040
rect 124956 270852 125008 270904
rect 178684 270852 178736 270904
rect 417424 270852 417476 270904
rect 427544 270852 427596 270904
rect 430396 270852 430448 270904
rect 483112 270852 483164 270904
rect 485228 270988 485280 271040
rect 490196 270988 490248 271040
rect 495256 270988 495308 271040
rect 575296 270988 575348 271040
rect 492404 270852 492456 270904
rect 492588 270852 492640 270904
rect 571616 270852 571668 270904
rect 571984 270852 572036 270904
rect 604828 270852 604880 270904
rect 127348 270716 127400 270768
rect 179880 270716 179932 270768
rect 321376 270716 321428 270768
rect 327080 270716 327132 270768
rect 427452 270716 427504 270768
rect 479156 270716 479208 270768
rect 486884 270716 486936 270768
rect 564624 270716 564676 270768
rect 137928 270580 137980 270632
rect 187700 270580 187752 270632
rect 422944 270580 422996 270632
rect 445300 270580 445352 270632
rect 489644 270580 489696 270632
rect 568212 270580 568264 270632
rect 129464 270444 129516 270496
rect 181168 270444 181220 270496
rect 191748 270444 191800 270496
rect 196900 270444 196952 270496
rect 201776 270444 201828 270496
rect 232228 270444 232280 270496
rect 395620 270444 395672 270496
rect 433616 270444 433668 270496
rect 453580 270444 453632 270496
rect 516784 270444 516836 270496
rect 517520 270444 517572 270496
rect 579620 270444 579672 270496
rect 581644 270444 581696 270496
rect 620284 270444 620336 270496
rect 88340 270308 88392 270360
rect 121460 270308 121512 270360
rect 122564 270308 122616 270360
rect 176200 270308 176252 270360
rect 180708 270308 180760 270360
rect 215300 270308 215352 270360
rect 232780 270308 232832 270360
rect 247868 270308 247920 270360
rect 262864 270308 262916 270360
rect 97908 270172 97960 270224
rect 158812 270172 158864 270224
rect 179328 270172 179380 270224
rect 214104 270172 214156 270224
rect 226616 270172 226668 270224
rect 249892 270172 249944 270224
rect 259736 270172 259788 270224
rect 367468 270308 367520 270360
rect 393504 270308 393556 270360
rect 400864 270308 400916 270360
rect 441620 270308 441672 270360
rect 456064 270308 456116 270360
rect 520280 270308 520332 270360
rect 85488 270036 85540 270088
rect 149428 270036 149480 270088
rect 173716 270036 173768 270088
rect 212632 270036 212684 270088
rect 216496 270036 216548 270088
rect 242440 270036 242492 270088
rect 248328 270036 248380 270088
rect 264796 270036 264848 270088
rect 70584 269900 70636 269952
rect 79968 269900 80020 269952
rect 80152 269900 80204 269952
rect 146392 269900 146444 269952
rect 165436 269900 165488 269952
rect 206008 269900 206060 269952
rect 210056 269900 210108 269952
rect 238300 269900 238352 269952
rect 241980 269900 242032 269952
rect 260380 269900 260432 269952
rect 271420 270172 271472 270224
rect 345112 270172 345164 270224
rect 361580 270172 361632 270224
rect 364156 270172 364208 270224
rect 389180 270172 389232 270224
rect 390100 270172 390152 270224
rect 405740 270172 405792 270224
rect 409696 270172 409748 270224
rect 454040 270172 454092 270224
rect 458548 270172 458600 270224
rect 524420 270308 524472 270360
rect 525616 270308 525668 270360
rect 523132 270172 523184 270224
rect 533160 270172 533212 270224
rect 533528 270308 533580 270360
rect 626540 270308 626592 270360
rect 619640 270172 619692 270224
rect 327724 270036 327776 270088
rect 336740 270036 336792 270088
rect 345940 270036 345992 270088
rect 362960 270036 363012 270088
rect 369860 270036 369912 270088
rect 396080 270036 396132 270088
rect 399852 270036 399904 270088
rect 412640 270036 412692 270088
rect 414664 270036 414716 270088
rect 460940 270036 460992 270088
rect 461400 270036 461452 270088
rect 527180 270036 527232 270088
rect 528376 270036 528428 270088
rect 623964 270172 624016 270224
rect 620284 270036 620336 270088
rect 630680 270036 630732 270088
rect 273076 269900 273128 269952
rect 326896 269900 326948 269952
rect 335544 269900 335596 269952
rect 336832 269900 336884 269952
rect 350540 269900 350592 269952
rect 351736 269900 351788 269952
rect 371240 269900 371292 269952
rect 372436 269900 372488 269952
rect 400496 269900 400548 269952
rect 401876 269900 401928 269952
rect 416780 269900 416832 269952
rect 417148 269900 417200 269952
rect 465080 269900 465132 269952
rect 468484 269900 468536 269952
rect 76748 269764 76800 269816
rect 143908 269764 143960 269816
rect 144368 269764 144420 269816
rect 190828 269764 190880 269816
rect 202972 269764 203024 269816
rect 233332 269764 233384 269816
rect 241428 269764 241480 269816
rect 259828 269764 259880 269816
rect 261944 269764 261996 269816
rect 274732 269764 274784 269816
rect 280068 269764 280120 269816
rect 287152 269764 287204 269816
rect 335084 269764 335136 269816
rect 347780 269764 347832 269816
rect 355048 269764 355100 269816
rect 376944 269764 376996 269816
rect 377680 269764 377732 269816
rect 408500 269764 408552 269816
rect 412456 269764 412508 269816
rect 458272 269764 458324 269816
rect 463516 269764 463568 269816
rect 531320 269764 531372 269816
rect 531964 269900 532016 269952
rect 533528 269900 533580 269952
rect 533988 269900 534040 269952
rect 537760 269900 537812 269952
rect 537944 269900 537996 269952
rect 538496 269764 538548 269816
rect 538680 269764 538732 269816
rect 542820 269764 542872 269816
rect 543188 269900 543240 269952
rect 640524 269900 640576 269952
rect 637580 269764 637632 269816
rect 126888 269628 126940 269680
rect 178316 269628 178368 269680
rect 200488 269628 200540 269680
rect 226892 269628 226944 269680
rect 384764 269628 384816 269680
rect 418252 269628 418304 269680
rect 422116 269628 422168 269680
rect 471980 269628 472032 269680
rect 472624 269628 472676 269680
rect 473360 269628 473412 269680
rect 78864 269492 78916 269544
rect 130384 269492 130436 269544
rect 133788 269492 133840 269544
rect 183652 269492 183704 269544
rect 186412 269492 186464 269544
rect 204076 269492 204128 269544
rect 392032 269492 392084 269544
rect 401692 269492 401744 269544
rect 404544 269492 404596 269544
rect 423680 269492 423732 269544
rect 432236 269492 432288 269544
rect 466460 269492 466512 269544
rect 530400 269628 530452 269680
rect 530584 269628 530636 269680
rect 531964 269628 532016 269680
rect 533160 269628 533212 269680
rect 616144 269628 616196 269680
rect 140688 269356 140740 269408
rect 188620 269356 188672 269408
rect 429108 269356 429160 269408
rect 455420 269356 455472 269408
rect 466000 269356 466052 269408
rect 509056 269492 509108 269544
rect 596180 269492 596232 269544
rect 474280 269356 474332 269408
rect 538128 269356 538180 269408
rect 538312 269356 538364 269408
rect 581644 269356 581696 269408
rect 121644 269220 121696 269272
rect 167828 269220 167880 269272
rect 272432 269220 272484 269272
rect 278872 269220 278924 269272
rect 423956 269220 424008 269272
rect 448520 269220 448572 269272
rect 470968 269220 471020 269272
rect 540612 269220 540664 269272
rect 540796 269220 540848 269272
rect 543188 269220 543240 269272
rect 543372 269152 543424 269204
rect 546500 269152 546552 269204
rect 274916 269084 274968 269136
rect 279700 269084 279752 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 42156 269016 42208 269068
rect 43168 269016 43220 269068
rect 84108 269016 84160 269068
rect 137468 269016 137520 269068
rect 137652 269016 137704 269068
rect 186136 269016 186188 269068
rect 379704 269016 379756 269068
rect 404360 269016 404412 269068
rect 436192 269016 436244 269068
rect 491760 269016 491812 269068
rect 498292 269016 498344 269068
rect 581000 269016 581052 269068
rect 273260 268948 273312 269000
rect 275560 268948 275612 269000
rect 111984 268880 112036 268932
rect 168748 268880 168800 268932
rect 382372 268880 382424 268932
rect 415400 268880 415452 268932
rect 433708 268880 433760 268932
rect 488540 268880 488592 268932
rect 500776 268880 500828 268932
rect 583760 268880 583812 268932
rect 115848 268744 115900 268796
rect 110236 268608 110288 268660
rect 102508 268472 102560 268524
rect 162952 268472 163004 268524
rect 92388 268336 92440 268388
rect 155500 268336 155552 268388
rect 211344 268744 211396 268796
rect 223488 268744 223540 268796
rect 389824 268744 389876 268796
rect 425336 268744 425388 268796
rect 441160 268744 441212 268796
rect 499580 268744 499632 268796
rect 503260 268744 503312 268796
rect 587900 268744 587952 268796
rect 167000 268608 167052 268660
rect 184480 268608 184532 268660
rect 187332 268608 187384 268660
rect 219440 268608 219492 268660
rect 245568 268608 245620 268660
rect 263140 268608 263192 268660
rect 403256 268608 403308 268660
rect 440240 268608 440292 268660
rect 443644 268608 443696 268660
rect 502340 268608 502392 268660
rect 505744 268608 505796 268660
rect 590844 268608 590896 268660
rect 171232 268472 171284 268524
rect 176936 268472 176988 268524
rect 215116 268472 215168 268524
rect 220452 268472 220504 268524
rect 245752 268472 245804 268524
rect 338488 268472 338540 268524
rect 350724 268472 350776 268524
rect 359832 268472 359884 268524
rect 379520 268472 379572 268524
rect 397092 268472 397144 268524
rect 433340 268472 433392 268524
rect 448612 268472 448664 268524
rect 509240 268472 509292 268524
rect 513196 268472 513248 268524
rect 601700 268472 601752 268524
rect 167644 268336 167696 268388
rect 168012 268336 168064 268388
rect 203524 268336 203576 268388
rect 203892 268336 203944 268388
rect 230756 268336 230808 268388
rect 231676 268336 231728 268388
rect 253204 268336 253256 268388
rect 258356 268336 258408 268388
rect 268936 268336 268988 268388
rect 348424 268336 348476 268388
rect 367100 268336 367152 268388
rect 372160 268336 372212 268388
rect 397460 268336 397512 268388
rect 408040 268336 408092 268388
rect 451372 268336 451424 268388
rect 464344 268336 464396 268388
rect 532700 268336 532752 268388
rect 541348 268336 541400 268388
rect 641720 268336 641772 268388
rect 128544 268200 128596 268252
rect 150440 268200 150492 268252
rect 151728 268200 151780 268252
rect 196072 268200 196124 268252
rect 419632 268200 419684 268252
rect 467932 268200 467984 268252
rect 493600 268200 493652 268252
rect 574100 268200 574152 268252
rect 163136 268064 163188 268116
rect 168012 268064 168064 268116
rect 412640 268064 412692 268116
rect 447140 268064 447192 268116
rect 495808 268064 495860 268116
rect 576860 268064 576912 268116
rect 198740 267792 198792 267844
rect 201868 267792 201920 267844
rect 117964 267656 118016 267708
rect 159640 267656 159692 267708
rect 167828 267656 167880 267708
rect 177028 267656 177080 267708
rect 181996 267656 182048 267708
rect 95884 267520 95936 267572
rect 138112 267520 138164 267572
rect 150440 267520 150492 267572
rect 181996 267520 182048 267572
rect 182732 267656 182784 267708
rect 214288 267656 214340 267708
rect 378232 267656 378284 267708
rect 392584 267656 392636 267708
rect 398104 267656 398156 267708
rect 414480 267656 414532 267708
rect 423772 267656 423824 267708
rect 440884 267656 440936 267708
rect 442724 267656 442776 267708
rect 493324 267656 493376 267708
rect 497832 267656 497884 267708
rect 517520 267656 517572 267708
rect 529664 267656 529716 267708
rect 585784 267656 585836 267708
rect 219256 267520 219308 267572
rect 340972 267520 341024 267572
rect 355324 267520 355376 267572
rect 370780 267520 370832 267572
rect 377404 267520 377456 267572
rect 380716 267520 380768 267572
rect 399852 267520 399904 267572
rect 410524 267520 410576 267572
rect 429108 267520 429160 267572
rect 445300 267520 445352 267572
rect 497464 267520 497516 267572
rect 514852 267520 514904 267572
rect 571984 267520 572036 267572
rect 86224 267384 86276 267436
rect 144736 267384 144788 267436
rect 146944 267384 146996 267436
rect 186964 267384 187016 267436
rect 236644 267384 236696 267436
rect 241612 267384 241664 267436
rect 315304 267384 315356 267436
rect 318984 267384 319036 267436
rect 350080 267384 350132 267436
rect 358084 267384 358136 267436
rect 362500 267384 362552 267436
rect 369308 267384 369360 267436
rect 371608 267384 371660 267436
rect 373264 267384 373316 267436
rect 383200 267384 383252 267436
rect 401876 267384 401928 267436
rect 405556 267384 405608 267436
rect 423956 267384 424008 267436
rect 432052 267384 432104 267436
rect 453304 267384 453356 267436
rect 460204 267384 460256 267436
rect 515404 267384 515456 267436
rect 519820 267384 519872 267436
rect 578884 267384 578936 267436
rect 104808 267248 104860 267300
rect 164608 267248 164660 267300
rect 169024 267248 169076 267300
rect 209320 267248 209372 267300
rect 218704 267248 218756 267300
rect 223028 267248 223080 267300
rect 223488 267248 223540 267300
rect 239128 267248 239180 267300
rect 314476 267248 314528 267300
rect 318800 267248 318852 267300
rect 353392 267248 353444 267300
rect 364984 267248 365036 267300
rect 373264 267248 373316 267300
rect 392032 267248 392084 267300
rect 403072 267248 403124 267300
rect 422944 267248 422996 267300
rect 424600 267248 424652 267300
rect 446404 267248 446456 267300
rect 448152 267248 448204 267300
rect 457444 267248 457496 267300
rect 470140 267248 470192 267300
rect 534724 267248 534776 267300
rect 543004 267248 543056 267300
rect 625804 267248 625856 267300
rect 79968 267112 80020 267164
rect 140596 267112 140648 267164
rect 144184 267112 144236 267164
rect 191932 267112 191984 267164
rect 192576 267112 192628 267164
rect 223948 267112 224000 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 312820 267112 312872 267164
rect 316040 267112 316092 267164
rect 365812 267112 365864 267164
rect 382924 267112 382976 267164
rect 390652 267112 390704 267164
rect 417424 267112 417476 267164
rect 417976 267112 418028 267164
rect 432236 267112 432288 267164
rect 432880 267112 432932 267164
rect 460020 267112 460072 267164
rect 465172 267112 465224 267164
rect 526444 267112 526496 267164
rect 534724 267112 534776 267164
rect 618904 267112 618956 267164
rect 90364 266976 90416 267028
rect 151360 266976 151412 267028
rect 154488 266976 154540 267028
rect 199384 266976 199436 267028
rect 218888 266976 218940 267028
rect 220084 266976 220136 267028
rect 228364 266976 228416 267028
rect 121460 266840 121512 266892
rect 144920 266840 144972 266892
rect 145380 266840 145432 266892
rect 150532 266840 150584 266892
rect 204076 266840 204128 266892
rect 220912 266840 220964 266892
rect 316960 266976 317012 267028
rect 321928 266976 321980 267028
rect 375748 266976 375800 267028
rect 390100 266976 390152 267028
rect 393136 266976 393188 267028
rect 420184 266976 420236 267028
rect 431224 266976 431276 267028
rect 432604 266976 432656 267028
rect 249064 266840 249116 266892
rect 286324 266840 286376 266892
rect 287980 266840 288032 266892
rect 321928 266840 321980 266892
rect 327540 266840 327592 266892
rect 332692 266840 332744 266892
rect 343824 266840 343876 266892
rect 392308 266840 392360 266892
rect 393964 266840 394016 266892
rect 427912 266840 427964 266892
rect 450544 266976 450596 267028
rect 455052 266976 455104 267028
rect 512644 266976 512696 267028
rect 524788 266976 524840 267028
rect 612004 266976 612056 267028
rect 450268 266840 450320 266892
rect 355876 266772 355928 266824
rect 374644 266772 374696 266824
rect 130384 266704 130436 266756
rect 147220 266704 147272 266756
rect 149704 266704 149756 266756
rect 169576 266704 169628 266756
rect 230756 266704 230808 266756
rect 234160 266704 234212 266756
rect 252008 266704 252060 266756
rect 259000 266704 259052 266756
rect 313648 266704 313700 266756
rect 317420 266704 317472 266756
rect 388168 266704 388220 266756
rect 214564 266636 214616 266688
rect 218428 266636 218480 266688
rect 308680 266636 308732 266688
rect 310520 266636 310572 266688
rect 317788 266636 317840 266688
rect 322940 266636 322992 266688
rect 342628 266636 342680 266688
rect 347044 266636 347096 266688
rect 137468 266568 137520 266620
rect 145380 266568 145432 266620
rect 145564 266568 145616 266620
rect 148048 266568 148100 266620
rect 226892 266568 226944 266620
rect 231676 266568 231728 266620
rect 394792 266704 394844 266756
rect 397092 266704 397144 266756
rect 397460 266704 397512 266756
rect 407764 266704 407816 266756
rect 428740 266704 428792 266756
rect 404544 266568 404596 266620
rect 404728 266568 404780 266620
rect 412640 266568 412692 266620
rect 440332 266704 440384 266756
rect 445024 266704 445076 266756
rect 457720 266704 457772 266756
rect 479524 266704 479576 266756
rect 442264 266568 442316 266620
rect 452752 266568 452804 266620
rect 469864 266568 469916 266620
rect 504824 266840 504876 266892
rect 513932 266840 513984 266892
rect 490012 266704 490064 266756
rect 507124 266704 507176 266756
rect 509884 266704 509936 266756
rect 516508 266704 516560 266756
rect 517336 266704 517388 266756
rect 518992 266840 519044 266892
rect 520096 266840 520148 266892
rect 527272 266840 527324 266892
rect 528192 266840 528244 266892
rect 528928 266840 528980 266892
rect 529848 266840 529900 266892
rect 531412 266840 531464 266892
rect 532516 266840 532568 266892
rect 533068 266840 533120 266892
rect 533988 266840 534040 266892
rect 535552 266840 535604 266892
rect 536748 266840 536800 266892
rect 539692 266840 539744 266892
rect 595444 266840 595496 266892
rect 563704 266704 563756 266756
rect 501604 266568 501656 266620
rect 214104 266500 214156 266552
rect 215944 266500 215996 266552
rect 248880 266500 248932 266552
rect 250720 266500 250772 266552
rect 310336 266500 310388 266552
rect 311900 266500 311952 266552
rect 312268 266500 312320 266552
rect 314660 266500 314712 266552
rect 316132 266500 316184 266552
rect 320180 266500 320232 266552
rect 347412 266500 347464 266552
rect 349804 266500 349856 266552
rect 350908 266500 350960 266552
rect 352564 266500 352616 266552
rect 357532 266500 357584 266552
rect 359832 266500 359884 266552
rect 144920 266432 144972 266484
rect 153844 266432 153896 266484
rect 162124 266364 162176 266416
rect 167092 266364 167144 266416
rect 178684 266364 178736 266416
rect 179512 266364 179564 266416
rect 215300 266364 215352 266416
rect 217600 266364 217652 266416
rect 219440 266364 219492 266416
rect 222568 266364 222620 266416
rect 224224 266364 224276 266416
rect 226708 266364 226760 266416
rect 233884 266364 233936 266416
rect 236644 266364 236696 266416
rect 239588 266364 239640 266416
rect 246580 266364 246632 266416
rect 250444 266364 250496 266416
rect 251548 266364 251600 266416
rect 253388 266364 253440 266416
rect 256516 266364 256568 266416
rect 287704 266364 287756 266416
rect 288808 266364 288860 266416
rect 301044 266364 301096 266416
rect 302056 266364 302108 266416
rect 303712 266364 303764 266416
rect 304540 266364 304592 266416
rect 307852 266364 307904 266416
rect 309140 266364 309192 266416
rect 309508 266364 309560 266416
rect 310980 266364 311032 266416
rect 311164 266364 311216 266416
rect 313280 266364 313332 266416
rect 320272 266364 320324 266416
rect 321376 266364 321428 266416
rect 324412 266364 324464 266416
rect 325332 266364 325384 266416
rect 328552 266364 328604 266416
rect 329472 266364 329524 266416
rect 330208 266364 330260 266416
rect 331956 266364 332008 266416
rect 334348 266364 334400 266416
rect 335268 266364 335320 266416
rect 346768 266364 346820 266416
rect 347596 266364 347648 266416
rect 349252 266364 349304 266416
rect 350356 266364 350408 266416
rect 352564 266364 352616 266416
rect 353944 266364 353996 266416
rect 359188 266364 359240 266416
rect 360108 266364 360160 266416
rect 360016 266228 360068 266280
rect 366364 266500 366416 266552
rect 374920 266500 374972 266552
rect 379704 266500 379756 266552
rect 482560 266500 482612 266552
rect 485044 266500 485096 266552
rect 491668 266432 491720 266484
rect 492588 266432 492640 266484
rect 494152 266432 494204 266484
rect 495256 266432 495308 266484
rect 499948 266432 500000 266484
rect 502432 266432 502484 266484
rect 503444 266432 503496 266484
rect 504088 266432 504140 266484
rect 505008 266432 505060 266484
rect 506572 266432 506624 266484
rect 507676 266432 507728 266484
rect 510712 266568 510764 266620
rect 511816 266568 511868 266620
rect 513932 266568 513984 266620
rect 556804 266568 556856 266620
rect 549904 266432 549956 266484
rect 361672 266364 361724 266416
rect 362776 266364 362828 266416
rect 368296 266364 368348 266416
rect 369124 266364 369176 266416
rect 369400 266364 369452 266416
rect 369860 266364 369912 266416
rect 370320 266364 370372 266416
rect 372160 266364 372212 266416
rect 374092 266364 374144 266416
rect 375196 266364 375248 266416
rect 379888 266364 379940 266416
rect 381544 266364 381596 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387432 266364 387484 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400036 266364 400088 266416
rect 400036 266228 400088 266280
rect 403256 266364 403308 266416
rect 407212 266364 407264 266416
rect 408224 266364 408276 266416
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 425428 266364 425480 266416
rect 427084 266364 427136 266416
rect 429568 266364 429620 266416
rect 430396 266364 430448 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 446128 266364 446180 266416
rect 447784 266364 447836 266416
rect 454408 266364 454460 266416
rect 455236 266364 455288 266416
rect 456892 266364 456944 266416
rect 458088 266364 458140 266416
rect 466828 266364 466880 266416
rect 467748 266364 467800 266416
rect 473452 266364 473504 266416
rect 474648 266364 474700 266416
rect 477592 266364 477644 266416
rect 478512 266364 478564 266416
rect 481732 266364 481784 266416
rect 482836 266364 482888 266416
rect 483388 266364 483440 266416
rect 484308 266364 484360 266416
rect 485872 266364 485924 266416
rect 487068 266364 487120 266416
rect 484216 266228 484268 266280
rect 560484 266296 560536 266348
rect 487528 266160 487580 266212
rect 565820 266160 565872 266212
rect 492496 266024 492548 266076
rect 572720 266024 572772 266076
rect 512368 265888 512420 265940
rect 600320 265888 600372 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 152004 265616 152056 265668
rect 152740 265616 152792 265668
rect 155960 265616 156012 265668
rect 156788 265616 156840 265668
rect 172520 265616 172572 265668
rect 173348 265616 173400 265668
rect 189172 265616 189224 265668
rect 189908 265616 189960 265668
rect 229100 265616 229152 265668
rect 229652 265616 229704 265668
rect 243084 265616 243136 265668
rect 243820 265616 243872 265668
rect 253940 265616 253992 265668
rect 254492 265616 254544 265668
rect 280344 265616 280396 265668
rect 280988 265616 281040 265668
rect 284300 265616 284352 265668
rect 285220 265616 285272 265668
rect 296812 265616 296864 265668
rect 297548 265616 297600 265668
rect 520648 265616 520700 265668
rect 612740 265616 612792 265668
rect 480076 265480 480128 265532
rect 554780 265480 554832 265532
rect 479248 265344 479300 265396
rect 553400 265344 553452 265396
rect 475108 265208 475160 265260
rect 547972 265208 548024 265260
rect 469312 265072 469364 265124
rect 539968 265072 540020 265124
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 676036 259564 676088 259616
rect 676220 259564 676272 259616
rect 554320 259428 554372 259480
rect 560944 259428 560996 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 563704 256708 563756 256760
rect 553492 255552 553544 255604
rect 555424 255552 555476 255604
rect 35808 255416 35860 255468
rect 39764 255416 39816 255468
rect 675852 254600 675904 254652
rect 683028 254600 683080 254652
rect 675024 254260 675076 254312
rect 675484 254260 675536 254312
rect 35808 254056 35860 254108
rect 39580 254056 39632 254108
rect 35808 252696 35860 252748
rect 41696 252696 41748 252748
rect 35624 252560 35676 252612
rect 40960 252560 41012 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 35808 251336 35860 251388
rect 40500 251336 40552 251388
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 35808 249908 35860 249960
rect 39396 249908 39448 249960
rect 35808 248480 35860 248532
rect 39212 248480 39264 248532
rect 35808 247188 35860 247240
rect 41696 247188 41748 247240
rect 35624 247052 35676 247104
rect 41512 247052 41564 247104
rect 558184 246304 558236 246356
rect 647240 246304 647292 246356
rect 553860 245624 553912 245676
rect 596824 245624 596876 245676
rect 554504 244264 554556 244316
rect 573364 244264 573416 244316
rect 674748 242700 674800 242752
rect 675300 242700 675352 242752
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553676 241476 553728 241528
rect 629944 241476 629996 241528
rect 554504 240116 554556 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 668768 236988 668820 237040
rect 671528 236988 671580 237040
rect 672080 236784 672132 236836
rect 671528 236580 671580 236632
rect 672954 236648 673006 236700
rect 671712 236444 671764 236496
rect 673184 236240 673236 236292
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 670976 235900 671028 235952
rect 673276 235900 673328 235952
rect 670148 235764 670200 235816
rect 672080 235764 672132 235816
rect 672632 235696 672684 235748
rect 673092 235492 673144 235544
rect 669596 235288 669648 235340
rect 668216 235084 668268 235136
rect 668400 234812 668452 234864
rect 674088 234676 674140 234728
rect 661684 234608 661736 234660
rect 670424 234608 670476 234660
rect 42432 234540 42484 234592
rect 42984 234540 43036 234592
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 669412 234472 669464 234524
rect 675116 234472 675168 234524
rect 671896 234336 671948 234388
rect 671160 234200 671212 234252
rect 674104 234200 674156 234252
rect 675852 233928 675904 233980
rect 683396 233928 683448 233980
rect 652392 233860 652444 233912
rect 674104 233792 674156 233844
rect 676036 233792 676088 233844
rect 678244 233792 678296 233844
rect 670332 233180 670384 233232
rect 672632 233180 672684 233232
rect 639604 232500 639656 232552
rect 654784 232500 654836 232552
rect 660304 232500 660356 232552
rect 675852 232500 675904 232552
rect 683212 232500 683264 232552
rect 671896 232432 671948 232484
rect 665456 231616 665508 231668
rect 674932 231616 674984 231668
rect 146208 231548 146260 231600
rect 150532 231548 150584 231600
rect 663064 231480 663116 231532
rect 671896 231480 671948 231532
rect 675852 231480 675904 231532
rect 683580 231480 683632 231532
rect 146760 231412 146812 231464
rect 147220 231412 147272 231464
rect 662328 231344 662380 231396
rect 675116 231344 675168 231396
rect 137928 231276 137980 231328
rect 152464 231276 152516 231328
rect 156512 231276 156564 231328
rect 163688 231276 163740 231328
rect 91744 231140 91796 231192
rect 168840 231140 168892 231192
rect 664996 231140 665048 231192
rect 596824 231072 596876 231124
rect 633624 231072 633676 231124
rect 636844 231072 636896 231124
rect 650644 231072 650696 231124
rect 128268 231004 128320 231056
rect 195888 231004 195940 231056
rect 675116 231004 675168 231056
rect 118608 230868 118660 230920
rect 188160 230868 188212 230920
rect 674956 230800 675008 230852
rect 110328 230732 110380 230784
rect 184296 230732 184348 230784
rect 97908 230596 97960 230648
rect 173992 230596 174044 230648
rect 195060 230596 195112 230648
rect 196900 230596 196952 230648
rect 672080 230596 672132 230648
rect 439320 230528 439372 230580
rect 152464 230460 152516 230512
rect 203616 230460 203668 230512
rect 42432 230392 42484 230444
rect 43076 230392 43128 230444
rect 130384 230392 130436 230444
rect 142436 230392 142488 230444
rect 142620 230392 142672 230444
rect 146208 230392 146260 230444
rect 147634 230392 147686 230444
rect 149520 230392 149572 230444
rect 206284 230392 206336 230444
rect 256424 230392 256476 230444
rect 276296 230392 276348 230444
rect 292488 230392 292540 230444
rect 308404 230392 308456 230444
rect 334992 230392 335044 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 526904 230392 526956 230444
rect 536104 230392 536156 230444
rect 674676 230392 674728 230444
rect 387432 230324 387484 230376
rect 388444 230324 388496 230376
rect 398104 230324 398156 230376
rect 399392 230324 399444 230376
rect 436100 230324 436152 230376
rect 436744 230324 436796 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 443828 230324 443880 230376
rect 444840 230324 444892 230376
rect 446404 230324 446456 230376
rect 448704 230324 448756 230376
rect 449624 230324 449676 230376
rect 450544 230324 450596 230376
rect 452844 230324 452896 230376
rect 454316 230324 454368 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 470876 230324 470928 230376
rect 471888 230324 471940 230376
rect 472164 230324 472216 230376
rect 473176 230324 473228 230376
rect 487620 230324 487672 230376
rect 488448 230324 488500 230376
rect 493416 230324 493468 230376
rect 496360 230324 496412 230376
rect 497280 230324 497332 230376
rect 498108 230324 498160 230376
rect 511448 230324 511500 230376
rect 517520 230324 517572 230376
rect 133788 230256 133840 230308
rect 202328 230256 202380 230308
rect 210424 230256 210476 230308
rect 261576 230256 261628 230308
rect 275652 230256 275704 230308
rect 313096 230256 313148 230308
rect 528836 230256 528888 230308
rect 539600 230256 539652 230308
rect 388444 230188 388496 230240
rect 391664 230188 391716 230240
rect 444472 230188 444524 230240
rect 447692 230188 447744 230240
rect 451556 230188 451608 230240
rect 453304 230188 453356 230240
rect 453488 230188 453540 230240
rect 455788 230188 455840 230240
rect 468300 230188 468352 230240
rect 469128 230188 469180 230240
rect 490196 230188 490248 230240
rect 493692 230188 493744 230240
rect 674564 230188 674616 230240
rect 95240 230120 95292 230172
rect 157294 230120 157346 230172
rect 157432 230120 157484 230172
rect 161112 230120 161164 230172
rect 176752 230120 176804 230172
rect 235816 230120 235868 230172
rect 264244 230120 264296 230172
rect 302792 230120 302844 230172
rect 302976 230120 303028 230172
rect 329840 230120 329892 230172
rect 334256 230120 334308 230172
rect 355600 230120 355652 230172
rect 521108 230120 521160 230172
rect 529204 230120 529256 230172
rect 532700 230120 532752 230172
rect 547144 230120 547196 230172
rect 454132 230052 454184 230104
rect 455328 230052 455380 230104
rect 491484 230052 491536 230104
rect 492496 230052 492548 230104
rect 126888 229984 126940 230036
rect 195060 229984 195112 230036
rect 195428 229984 195480 230036
rect 214748 229984 214800 230036
rect 219992 229984 220044 230036
rect 230664 229984 230716 230036
rect 242532 229984 242584 230036
rect 287336 229984 287388 230036
rect 287520 229984 287572 230036
rect 307944 229984 307996 230036
rect 312636 229984 312688 230036
rect 340144 229984 340196 230036
rect 354956 229984 355008 230036
rect 371056 229984 371108 230036
rect 476672 229984 476724 230036
rect 481640 229984 481692 230036
rect 515312 229984 515364 230036
rect 524604 229984 524656 230036
rect 534632 229984 534684 230036
rect 549260 229984 549312 230036
rect 674452 229916 674504 229968
rect 86224 229848 86276 229900
rect 156696 229848 156748 229900
rect 68284 229712 68336 229764
rect 142620 229712 142672 229764
rect 147772 229712 147824 229764
rect 158536 229848 158588 229900
rect 163964 229848 164016 229900
rect 225512 229848 225564 229900
rect 230480 229848 230532 229900
rect 277032 229848 277084 229900
rect 282552 229848 282604 229900
rect 318248 229848 318300 229900
rect 324228 229848 324280 229900
rect 350448 229848 350500 229900
rect 366732 229848 366784 229900
rect 383936 229848 383988 229900
rect 457352 229848 457404 229900
rect 464068 229848 464120 229900
rect 469588 229848 469640 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 82084 229576 82136 229628
rect 147128 229508 147180 229560
rect 157294 229712 157346 229764
rect 166264 229712 166316 229764
rect 171048 229712 171100 229764
rect 219992 229712 220044 229764
rect 148140 229576 148192 229628
rect 155960 229576 156012 229628
rect 157340 229576 157392 229628
rect 102140 229440 102192 229492
rect 144000 229440 144052 229492
rect 144184 229440 144236 229492
rect 146944 229440 146996 229492
rect 111064 229304 111116 229356
rect 147588 229304 147640 229356
rect 147772 229304 147824 229356
rect 210056 229440 210108 229492
rect 214748 229576 214800 229628
rect 246120 229712 246172 229764
rect 256516 229712 256568 229764
rect 297640 229712 297692 229764
rect 318064 229712 318116 229764
rect 220360 229440 220412 229492
rect 220728 229440 220780 229492
rect 266728 229576 266780 229628
rect 296996 229576 297048 229628
rect 323400 229576 323452 229628
rect 345020 229712 345072 229764
rect 360752 229712 360804 229764
rect 361212 229712 361264 229764
rect 378784 229712 378836 229764
rect 391204 229712 391256 229764
rect 398748 229712 398800 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 410892 229712 410944 229764
rect 417424 229712 417476 229764
rect 467012 229712 467064 229764
rect 474004 229712 474056 229764
rect 481824 229848 481876 229900
rect 489920 229848 489972 229900
rect 495992 229848 496044 229900
rect 506572 229848 506624 229900
rect 510804 229848 510856 229900
rect 511908 229848 511960 229900
rect 517244 229848 517296 229900
rect 525984 229848 526036 229900
rect 536564 229848 536616 229900
rect 559564 229848 559616 229900
rect 476028 229780 476080 229832
rect 478604 229780 478656 229832
rect 673460 229780 673512 229832
rect 479248 229712 479300 229764
rect 488080 229712 488132 229764
rect 492128 229712 492180 229764
rect 505192 229712 505244 229764
rect 507584 229712 507636 229764
rect 516784 229712 516836 229764
rect 523040 229712 523092 229764
rect 534816 229712 534868 229764
rect 538496 229712 538548 229764
rect 566464 229712 566516 229764
rect 476764 229644 476816 229696
rect 345296 229576 345348 229628
rect 463792 229576 463844 229628
rect 465724 229576 465776 229628
rect 509516 229576 509568 229628
rect 515404 229576 515456 229628
rect 530124 229576 530176 229628
rect 531136 229576 531188 229628
rect 384304 229508 384356 229560
rect 389088 229508 389140 229560
rect 448980 229508 449032 229560
rect 451924 229508 451976 229560
rect 231124 229440 231176 229492
rect 271880 229440 271932 229492
rect 465448 229440 465500 229492
rect 467472 229440 467524 229492
rect 488264 229440 488316 229492
rect 490380 229440 490432 229492
rect 530768 229440 530820 229492
rect 538312 229576 538364 229628
rect 673920 229576 673972 229628
rect 450912 229372 450964 229424
rect 453028 229372 453080 229424
rect 151176 229304 151228 229356
rect 123484 229168 123536 229220
rect 153384 229168 153436 229220
rect 153844 229304 153896 229356
rect 156512 229304 156564 229356
rect 157064 229304 157116 229356
rect 215208 229304 215260 229356
rect 246488 229304 246540 229356
rect 282184 229304 282236 229356
rect 413836 229304 413888 229356
rect 420000 229304 420052 229356
rect 674104 229304 674156 229356
rect 450268 229236 450320 229288
rect 451740 229236 451792 229288
rect 495348 229236 495400 229288
rect 500224 229236 500276 229288
rect 505652 229236 505704 229288
rect 510620 229236 510672 229288
rect 513380 229236 513432 229288
rect 519360 229236 519412 229288
rect 161756 229168 161808 229220
rect 184664 229168 184716 229220
rect 240968 229168 241020 229220
rect 100668 229032 100720 229084
rect 106188 229032 106240 229084
rect 142988 229032 143040 229084
rect 143448 229032 143500 229084
rect 146208 229032 146260 229084
rect 146392 229032 146444 229084
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 503720 229100 503772 229152
rect 509884 229100 509936 229152
rect 519176 229100 519228 229152
rect 205548 229032 205600 229084
rect 206008 229032 206060 229084
rect 214380 229032 214432 229084
rect 214748 229032 214800 229084
rect 257068 229032 257120 229084
rect 257528 229032 257580 229084
rect 296352 229032 296404 229084
rect 302148 229032 302200 229084
rect 331128 229032 331180 229084
rect 524972 229100 525024 229152
rect 529940 229100 529992 229152
rect 660948 229100 661000 229152
rect 665456 229100 665508 229152
rect 169300 228896 169352 228948
rect 172336 228896 172388 228948
rect 179696 228896 179748 228948
rect 180064 228896 180116 228948
rect 93768 228760 93820 228812
rect 166816 228760 166868 228812
rect 172152 228760 172204 228812
rect 174636 228760 174688 228812
rect 174820 228760 174872 228812
rect 219808 228760 219860 228812
rect 220360 228896 220412 228948
rect 246764 228896 246816 228948
rect 257712 228896 257764 228948
rect 299572 228896 299624 228948
rect 300676 228896 300728 228948
rect 330484 228896 330536 228948
rect 502432 228896 502484 228948
rect 521016 228896 521068 228948
rect 542820 228896 542872 228948
rect 673460 228896 673512 228948
rect 226156 228760 226208 228812
rect 238576 228760 238628 228812
rect 282828 228760 282880 228812
rect 296628 228760 296680 228812
rect 329196 228760 329248 228812
rect 336464 228760 336516 228812
rect 358820 228760 358872 228812
rect 359924 228760 359976 228812
rect 376852 228760 376904 228812
rect 478880 228760 478932 228812
rect 490196 228760 490248 228812
rect 518532 228760 518584 228812
rect 541624 228760 541676 228812
rect 67548 228624 67600 228676
rect 61660 228488 61712 228540
rect 142620 228488 142672 228540
rect 57244 228352 57296 228404
rect 141148 228352 141200 228404
rect 142988 228624 143040 228676
rect 152464 228624 152516 228676
rect 153108 228624 153160 228676
rect 142988 228488 143040 228540
rect 145932 228488 145984 228540
rect 146116 228488 146168 228540
rect 202420 228488 202472 228540
rect 214380 228624 214432 228676
rect 220360 228624 220412 228676
rect 220544 228624 220596 228676
rect 264796 228624 264848 228676
rect 285496 228624 285548 228676
rect 318892 228624 318944 228676
rect 325516 228624 325568 228676
rect 349160 228624 349212 228676
rect 350172 228624 350224 228676
rect 369124 228624 369176 228676
rect 377772 228624 377824 228676
rect 390376 228624 390428 228676
rect 498568 228624 498620 228676
rect 515772 228624 515824 228676
rect 517888 228624 517940 228676
rect 539416 228624 539468 228676
rect 539600 228624 539652 228676
rect 555976 228624 556028 228676
rect 215852 228488 215904 228540
rect 216220 228488 216272 228540
rect 219624 228488 219676 228540
rect 219992 228488 220044 228540
rect 260288 228488 260340 228540
rect 268936 228488 268988 228540
rect 306012 228488 306064 228540
rect 313924 228488 313976 228540
rect 320824 228488 320876 228540
rect 326896 228488 326948 228540
rect 351092 228488 351144 228540
rect 354588 228488 354640 228540
rect 372344 228488 372396 228540
rect 373448 228488 373500 228540
rect 387156 228488 387208 228540
rect 390468 228488 390520 228540
rect 400036 228488 400088 228540
rect 148876 228352 148928 228404
rect 152464 228352 152516 228404
rect 166816 228352 166868 228404
rect 166954 228352 167006 228404
rect 214564 228352 214616 228404
rect 217508 228352 217560 228404
rect 221464 228352 221516 228404
rect 224592 228352 224644 228404
rect 273812 228352 273864 228404
rect 274272 228352 274324 228404
rect 312452 228352 312504 228404
rect 320088 228352 320140 228404
rect 346860 228352 346912 228404
rect 347044 228352 347096 228404
rect 365904 228352 365956 228404
rect 371148 228352 371200 228404
rect 385224 228352 385276 228404
rect 386236 228352 386288 228404
rect 397460 228352 397512 228404
rect 112812 228216 112864 228268
rect 184940 228216 184992 228268
rect 189724 228216 189776 228268
rect 239036 228216 239088 228268
rect 254952 228216 255004 228268
rect 295708 228216 295760 228268
rect 407764 228488 407816 228540
rect 409788 228488 409840 228540
rect 415492 228488 415544 228540
rect 485688 228488 485740 228540
rect 498292 228488 498344 228540
rect 499856 228488 499908 228540
rect 517704 228488 517756 228540
rect 527548 228488 527600 228540
rect 553308 228488 553360 228540
rect 555424 228488 555476 228540
rect 571340 228488 571392 228540
rect 402796 228352 402848 228404
rect 411628 228352 411680 228404
rect 474464 228352 474516 228404
rect 484584 228352 484636 228404
rect 485044 228352 485096 228404
rect 498568 228352 498620 228404
rect 506572 228352 506624 228404
rect 512092 228352 512144 228404
rect 533528 228352 533580 228404
rect 537208 228352 537260 228404
rect 565636 228352 565688 228404
rect 663524 228352 663576 228404
rect 672080 228352 672132 228404
rect 512736 228216 512788 228268
rect 539416 228216 539468 228268
rect 540888 228216 540940 228268
rect 119988 228080 120040 228132
rect 190092 228080 190144 228132
rect 192944 228080 192996 228132
rect 126704 227944 126756 227996
rect 195244 227944 195296 227996
rect 202420 228080 202472 228132
rect 210700 228080 210752 228132
rect 213920 228080 213972 228132
rect 214380 228080 214432 228132
rect 214564 228080 214616 228132
rect 206008 227944 206060 227996
rect 88248 227808 88300 227860
rect 95240 227808 95292 227860
rect 133512 227808 133564 227860
rect 200396 227808 200448 227860
rect 203524 227808 203576 227860
rect 42432 227672 42484 227724
rect 43260 227672 43312 227724
rect 64788 227672 64840 227724
rect 111064 227672 111116 227724
rect 117228 227672 117280 227724
rect 187516 227672 187568 227724
rect 187700 227672 187752 227724
rect 110144 227536 110196 227588
rect 182364 227536 182416 227588
rect 185400 227536 185452 227588
rect 192668 227536 192720 227588
rect 200028 227672 200080 227724
rect 204904 227672 204956 227724
rect 205456 227808 205508 227860
rect 214748 227944 214800 227996
rect 219808 228080 219860 228132
rect 231308 228080 231360 228132
rect 233884 228080 233936 228132
rect 272524 228080 272576 228132
rect 400128 228080 400180 228132
rect 415032 228012 415084 228064
rect 421932 228012 421984 228064
rect 221004 227944 221056 227996
rect 221464 227944 221516 227996
rect 251272 227944 251324 227996
rect 416688 227876 416740 227928
rect 420644 227876 420696 227928
rect 447048 227876 447100 227928
rect 450544 227876 450596 227928
rect 210976 227808 211028 227860
rect 219992 227808 220044 227860
rect 226156 227808 226208 227860
rect 233884 227808 233936 227860
rect 239312 227808 239364 227860
rect 243544 227808 243596 227860
rect 246304 227808 246356 227860
rect 248696 227808 248748 227860
rect 249064 227808 249116 227860
rect 253848 227808 253900 227860
rect 331036 227740 331088 227792
rect 334256 227740 334308 227792
rect 351092 227740 351144 227792
rect 353024 227740 353076 227792
rect 371792 227740 371844 227792
rect 373632 227740 373684 227792
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 420644 227740 420696 227792
rect 423864 227740 423916 227792
rect 471520 227740 471572 227792
rect 479524 227740 479576 227792
rect 489920 227740 489972 227792
rect 494520 227740 494572 227792
rect 660488 227740 660540 227792
rect 665180 227740 665232 227792
rect 668952 227740 669004 227792
rect 672724 227740 672776 227792
rect 217784 227672 217836 227724
rect 219808 227672 219860 227724
rect 228732 227672 228784 227724
rect 228916 227672 228968 227724
rect 268016 227672 268068 227724
rect 291016 227672 291068 227724
rect 322112 227672 322164 227724
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 214748 227536 214800 227588
rect 214932 227536 214984 227588
rect 262220 227536 262272 227588
rect 281356 227536 281408 227588
rect 317604 227536 317656 227588
rect 322112 227536 322164 227588
rect 332416 227536 332468 227588
rect 337752 227536 337804 227588
rect 345020 227536 345072 227588
rect 524604 227536 524656 227588
rect 537484 227536 537536 227588
rect 60648 227400 60700 227452
rect 102140 227400 102192 227452
rect 103428 227400 103480 227452
rect 171232 227400 171284 227452
rect 172152 227400 172204 227452
rect 177212 227400 177264 227452
rect 181352 227400 181404 227452
rect 96436 227264 96488 227316
rect 89628 227128 89680 227180
rect 156696 227128 156748 227180
rect 169484 227264 169536 227316
rect 159640 227128 159692 227180
rect 185584 227264 185636 227316
rect 186136 227400 186188 227452
rect 187700 227400 187752 227452
rect 189908 227400 189960 227452
rect 204720 227400 204772 227452
rect 204904 227400 204956 227452
rect 251916 227400 251968 227452
rect 264796 227400 264848 227452
rect 304724 227400 304776 227452
rect 315488 227400 315540 227452
rect 341432 227400 341484 227452
rect 352564 227400 352616 227452
rect 363328 227400 363380 227452
rect 494704 227400 494756 227452
rect 511080 227400 511132 227452
rect 514024 227400 514076 227452
rect 535736 227400 535788 227452
rect 536104 227400 536156 227452
rect 552664 227400 552716 227452
rect 219532 227264 219584 227316
rect 219992 227264 220044 227316
rect 241612 227264 241664 227316
rect 249248 227264 249300 227316
rect 290556 227264 290608 227316
rect 293776 227264 293828 227316
rect 325332 227264 325384 227316
rect 333888 227264 333940 227316
rect 356244 227264 356296 227316
rect 357256 227264 357308 227316
rect 374276 227264 374328 227316
rect 382096 227264 382148 227316
rect 392952 227264 393004 227316
rect 171600 227128 171652 227180
rect 219808 227128 219860 227180
rect 56508 226992 56560 227044
rect 142160 226992 142212 227044
rect 143264 226992 143316 227044
rect 204076 226992 204128 227044
rect 122748 226856 122800 226908
rect 185400 226856 185452 226908
rect 185584 226856 185636 226908
rect 214104 226992 214156 227044
rect 233700 227128 233752 227180
rect 241152 227128 241204 227180
rect 286692 227128 286744 227180
rect 306196 227128 306248 227180
rect 336924 227128 336976 227180
rect 340696 227128 340748 227180
rect 361396 227128 361448 227180
rect 363512 227128 363564 227180
rect 368480 227128 368532 227180
rect 376668 227128 376720 227180
rect 389732 227128 389784 227180
rect 393136 227128 393188 227180
rect 402612 227264 402664 227316
rect 510620 227264 510672 227316
rect 524420 227264 524472 227316
rect 526260 227264 526312 227316
rect 551560 227264 551612 227316
rect 402244 227128 402296 227180
rect 408408 227128 408460 227180
rect 478604 227128 478656 227180
rect 486792 227128 486844 227180
rect 490380 227128 490432 227180
rect 502984 227128 503036 227180
rect 505008 227128 505060 227180
rect 523040 227128 523092 227180
rect 523684 227128 523736 227180
rect 548340 227128 548392 227180
rect 556804 227128 556856 227180
rect 570604 227128 570656 227180
rect 668584 227128 668636 227180
rect 673276 227128 673328 227180
rect 221832 226992 221884 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 308588 226992 308640 227044
rect 310336 226992 310388 227044
rect 338212 226992 338264 227044
rect 338672 226992 338724 227044
rect 360108 226992 360160 227044
rect 362776 226992 362828 227044
rect 379060 226992 379112 227044
rect 391756 226992 391808 227044
rect 403532 226992 403584 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 486976 226992 487028 227044
rect 500960 226992 501012 227044
rect 506296 226992 506348 227044
rect 526536 226992 526588 227044
rect 533344 226992 533396 227044
rect 560760 226992 560812 227044
rect 652208 226992 652260 227044
rect 129556 226720 129608 226772
rect 197452 226720 197504 226772
rect 204720 226720 204772 226772
rect 214748 226856 214800 226908
rect 219992 226856 220044 226908
rect 214104 226720 214156 226772
rect 218428 226720 218480 226772
rect 219348 226720 219400 226772
rect 267372 226856 267424 226908
rect 378784 226788 378836 226840
rect 385868 226788 385920 226840
rect 673460 226788 673512 226840
rect 235816 226720 235868 226772
rect 280252 226720 280304 226772
rect 136548 226584 136600 226636
rect 203156 226584 203208 226636
rect 204076 226584 204128 226636
rect 208124 226584 208176 226636
rect 212172 226584 212224 226636
rect 214932 226584 214984 226636
rect 219532 226584 219584 226636
rect 223580 226584 223632 226636
rect 225604 226584 225656 226636
rect 238392 226584 238444 226636
rect 259368 226584 259420 226636
rect 298284 226584 298336 226636
rect 673276 226516 673328 226568
rect 106924 226448 106976 226500
rect 146576 226448 146628 226500
rect 150072 226448 150124 226500
rect 213276 226448 213328 226500
rect 216404 226448 216456 226500
rect 220544 226448 220596 226500
rect 220728 226448 220780 226500
rect 228916 226448 228968 226500
rect 369124 226448 369176 226500
rect 376208 226448 376260 226500
rect 403992 226448 404044 226500
rect 412272 226448 412324 226500
rect 474740 226448 474792 226500
rect 482744 226448 482796 226500
rect 386052 226380 386104 226432
rect 391204 226380 391256 226432
rect 672724 226380 672776 226432
rect 407764 226312 407816 226364
rect 408684 226312 408736 226364
rect 481640 226312 481692 226364
rect 487804 226312 487856 226364
rect 488080 226312 488132 226364
rect 490012 226312 490064 226364
rect 122564 226244 122616 226296
rect 193956 226244 194008 226296
rect 194140 226244 194192 226296
rect 204904 226244 204956 226296
rect 205088 226244 205140 226296
rect 254492 226244 254544 226296
rect 260656 226244 260708 226296
rect 298928 226244 298980 226296
rect 308864 226244 308916 226296
rect 336280 226244 336332 226296
rect 388628 226244 388680 226296
rect 394240 226244 394292 226296
rect 72424 226108 72476 226160
rect 141148 226108 141200 226160
rect 141516 226108 141568 226160
rect 145012 226108 145064 226160
rect 145196 226108 145248 226160
rect 146760 226108 146812 226160
rect 148968 226108 149020 226160
rect 213460 226108 213512 226160
rect 213644 226108 213696 226160
rect 219992 226108 220044 226160
rect 222016 226108 222068 226160
rect 269948 226108 270000 226160
rect 270224 226108 270276 226160
rect 287520 226108 287572 226160
rect 288072 226108 288124 226160
rect 322756 226108 322808 226160
rect 525984 226108 526036 226160
rect 539968 226244 540020 226296
rect 563704 226244 563756 226296
rect 568120 226244 568172 226296
rect 83464 225972 83516 226024
rect 163044 225972 163096 226024
rect 196624 225972 196676 226024
rect 236460 225972 236512 226024
rect 252468 225972 252520 226024
rect 293132 225972 293184 226024
rect 299388 225972 299440 226024
rect 328552 225972 328604 226024
rect 335176 225972 335228 226024
rect 356888 225972 356940 226024
rect 361212 225972 361264 226024
rect 377496 225972 377548 226024
rect 498108 225972 498160 226024
rect 514300 225972 514352 226024
rect 516600 225972 516652 226024
rect 538496 226108 538548 226160
rect 672604 226108 672656 226160
rect 672080 226040 672132 226092
rect 538312 225972 538364 226024
rect 557264 225972 557316 226024
rect 76564 225836 76616 225888
rect 158260 225836 158312 225888
rect 169668 225836 169720 225888
rect 171600 225836 171652 225888
rect 171784 225836 171836 225888
rect 204536 225836 204588 225888
rect 204904 225836 204956 225888
rect 213644 225836 213696 225888
rect 219992 225836 220044 225888
rect 244188 225836 244240 225888
rect 261852 225836 261904 225888
rect 300860 225836 300912 225888
rect 312912 225836 312964 225888
rect 341708 225836 341760 225888
rect 341984 225836 342036 225888
rect 365260 225836 365312 225888
rect 375012 225836 375064 225888
rect 387800 225836 387852 225888
rect 394332 225836 394384 225888
rect 403256 225836 403308 225888
rect 501144 225836 501196 225888
rect 519176 225836 519228 225888
rect 521752 225836 521804 225888
rect 545764 225836 545816 225888
rect 672264 225836 672316 225888
rect 458640 225768 458692 225820
rect 462964 225768 463016 225820
rect 66168 225700 66220 225752
rect 149796 225700 149848 225752
rect 151268 225700 151320 225752
rect 58992 225564 59044 225616
rect 141516 225564 141568 225616
rect 141792 225564 141844 225616
rect 203156 225564 203208 225616
rect 204904 225700 204956 225752
rect 248880 225700 248932 225752
rect 251088 225700 251140 225752
rect 294420 225700 294472 225752
rect 296444 225700 296496 225752
rect 327908 225700 327960 225752
rect 329748 225700 329800 225752
rect 353668 225700 353720 225752
rect 365352 225700 365404 225752
rect 383292 225700 383344 225752
rect 387708 225700 387760 225752
rect 397828 225700 397880 225752
rect 481180 225700 481232 225752
rect 492680 225700 492732 225752
rect 493692 225700 493744 225752
rect 505376 225700 505428 225752
rect 508872 225700 508924 225752
rect 529204 225700 529256 225752
rect 535920 225700 535972 225752
rect 563060 225700 563112 225752
rect 672264 225632 672316 225684
rect 217140 225564 217192 225616
rect 217876 225564 217928 225616
rect 266084 225564 266136 225616
rect 267004 225564 267056 225616
rect 274456 225564 274508 225616
rect 278412 225564 278464 225616
rect 313280 225564 313332 225616
rect 327724 225564 327776 225616
rect 352380 225564 352432 225616
rect 352932 225564 352984 225616
rect 371608 225564 371660 225616
rect 382924 225564 382976 225616
rect 396172 225564 396224 225616
rect 410984 225564 411036 225616
rect 416136 225564 416188 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 488724 225564 488776 225616
rect 489368 225564 489420 225616
rect 503168 225564 503220 225616
rect 510160 225564 510212 225616
rect 530584 225564 530636 225616
rect 531412 225564 531464 225616
rect 558184 225564 558236 225616
rect 125232 225428 125284 225480
rect 196164 225428 196216 225480
rect 198004 225428 198056 225480
rect 204904 225428 204956 225480
rect 209596 225428 209648 225480
rect 259644 225428 259696 225480
rect 297364 225428 297416 225480
rect 310520 225428 310572 225480
rect 671896 225428 671948 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 129372 225292 129424 225344
rect 199108 225292 199160 225344
rect 203156 225292 203208 225344
rect 209412 225292 209464 225344
rect 62028 225156 62080 225208
rect 130384 225156 130436 225208
rect 135076 225156 135128 225208
rect 204260 225156 204312 225208
rect 204536 225156 204588 225208
rect 222936 225292 222988 225344
rect 242900 225292 242952 225344
rect 285036 225292 285088 225344
rect 215208 225156 215260 225208
rect 217876 225156 217928 225208
rect 426440 225156 426492 225208
rect 426992 225156 427044 225208
rect 666468 225156 666520 225208
rect 132408 225020 132460 225072
rect 201684 225020 201736 225072
rect 203892 225020 203944 225072
rect 255136 225020 255188 225072
rect 672034 225088 672086 225140
rect 355232 224952 355284 225004
rect 358176 224952 358228 225004
rect 404176 224952 404228 225004
rect 410616 224952 410668 225004
rect 416504 224952 416556 225004
rect 422208 224952 422260 225004
rect 96252 224884 96304 224936
rect 172980 224884 173032 224936
rect 89444 224748 89496 224800
rect 168196 224748 168248 224800
rect 171968 224748 172020 224800
rect 177488 224884 177540 224936
rect 199752 224884 199804 224936
rect 199936 224884 199988 224936
rect 248052 224884 248104 224936
rect 272524 224884 272576 224936
rect 309876 224884 309928 224936
rect 319812 224884 319864 224936
rect 345940 224884 345992 224936
rect 519360 224884 519412 224936
rect 535000 224884 535052 224936
rect 621020 224884 621072 224936
rect 232596 224748 232648 224800
rect 245476 224748 245528 224800
rect 287704 224748 287756 224800
rect 311532 224748 311584 224800
rect 338856 224748 338908 224800
rect 462504 224748 462556 224800
rect 469312 224748 469364 224800
rect 506940 224748 506992 224800
rect 526352 224748 526404 224800
rect 529940 224748 529992 224800
rect 350356 224680 350408 224732
rect 354956 224680 355008 224732
rect 79968 224612 80020 224664
rect 160468 224612 160520 224664
rect 165160 224612 165212 224664
rect 227444 224612 227496 224664
rect 228732 224612 228784 224664
rect 274916 224612 274968 224664
rect 275100 224612 275152 224664
rect 311164 224612 311216 224664
rect 322848 224612 322900 224664
rect 349804 224612 349856 224664
rect 359464 224612 359516 224664
rect 378140 224612 378192 224664
rect 494060 224612 494112 224664
rect 510160 224612 510212 224664
rect 520464 224612 520516 224664
rect 544384 224612 544436 224664
rect 549260 224748 549312 224800
rect 557080 224748 557132 224800
rect 557264 224748 557316 224800
rect 626540 224748 626592 224800
rect 671820 224680 671872 224732
rect 549996 224612 550048 224664
rect 625252 224612 625304 224664
rect 668032 224612 668084 224664
rect 85488 224476 85540 224528
rect 165620 224476 165672 224528
rect 165988 224476 166040 224528
rect 185400 224476 185452 224528
rect 185584 224476 185636 224528
rect 237748 224476 237800 224528
rect 248328 224476 248380 224528
rect 291844 224476 291896 224528
rect 294880 224476 294932 224528
rect 325976 224476 326028 224528
rect 331864 224476 331916 224528
rect 337568 224476 337620 224528
rect 346308 224476 346360 224528
rect 366548 224476 366600 224528
rect 379244 224476 379296 224528
rect 393596 224476 393648 224528
rect 447508 224476 447560 224528
rect 448060 224476 448112 224528
rect 456064 224476 456116 224528
rect 459744 224476 459796 224528
rect 491300 224476 491352 224528
rect 506020 224476 506072 224528
rect 515956 224476 516008 224528
rect 538956 224476 539008 224528
rect 542452 224476 542504 224528
rect 542820 224476 542872 224528
rect 623228 224476 623280 224528
rect 671252 224408 671304 224460
rect 73712 224340 73764 224392
rect 155316 224340 155368 224392
rect 155868 224340 155920 224392
rect 159640 224340 159692 224392
rect 161664 224340 161716 224392
rect 224868 224340 224920 224392
rect 233148 224340 233200 224392
rect 277676 224340 277728 224392
rect 289636 224340 289688 224392
rect 296996 224340 297048 224392
rect 299112 224340 299164 224392
rect 331404 224340 331456 224392
rect 342168 224340 342220 224392
rect 362040 224340 362092 224392
rect 366732 224340 366784 224392
rect 381636 224340 381688 224392
rect 394516 224340 394568 224392
rect 404544 224340 404596 224392
rect 480536 224340 480588 224392
rect 492864 224340 492916 224392
rect 499212 224340 499264 224392
rect 516784 224340 516836 224392
rect 525616 224340 525668 224392
rect 550640 224340 550692 224392
rect 554964 224272 555016 224324
rect 555884 224272 555936 224324
rect 625988 224340 626040 224392
rect 68928 224204 68980 224256
rect 152740 224204 152792 224256
rect 168012 224204 168064 224256
rect 230020 224204 230072 224256
rect 231676 224204 231728 224256
rect 278964 224204 279016 224256
rect 286324 224204 286376 224256
rect 289912 224204 289964 224256
rect 290832 224204 290884 224256
rect 324044 224204 324096 224256
rect 339408 224204 339460 224256
rect 362316 224204 362368 224256
rect 372528 224204 372580 224256
rect 387432 224204 387484 224256
rect 390192 224204 390244 224256
rect 401968 224204 402020 224256
rect 405556 224204 405608 224256
rect 414204 224204 414256 224256
rect 470232 224204 470284 224256
rect 480352 224204 480404 224256
rect 483756 224204 483808 224256
rect 497464 224204 497516 224256
rect 102048 224068 102100 224120
rect 178500 224068 178552 224120
rect 179328 224068 179380 224120
rect 185584 224068 185636 224120
rect 194784 224068 194836 224120
rect 250628 224068 250680 224120
rect 266268 224068 266320 224120
rect 303436 224068 303488 224120
rect 304264 224068 304316 224120
rect 315304 224068 315356 224120
rect 504364 224068 504416 224120
rect 523500 224204 523552 224256
rect 535276 224204 535328 224256
rect 562324 224204 562376 224256
rect 571432 224204 571484 224256
rect 651288 224204 651340 224256
rect 666468 224204 666520 224256
rect 667848 224204 667900 224256
rect 562140 224136 562192 224188
rect 539968 224000 540020 224052
rect 622584 224000 622636 224052
rect 669044 224000 669096 224052
rect 106004 223932 106056 223984
rect 181076 223932 181128 223984
rect 185400 223932 185452 223984
rect 194600 223932 194652 223984
rect 194968 223932 195020 223984
rect 199844 223932 199896 223984
rect 201408 223932 201460 223984
rect 255780 223932 255832 223984
rect 279424 223864 279476 223916
rect 284760 223864 284812 223916
rect 524420 223864 524472 223916
rect 525064 223864 525116 223916
rect 619640 223864 619692 223916
rect 108672 223796 108724 223848
rect 183652 223796 183704 223848
rect 184388 223796 184440 223848
rect 207480 223796 207532 223848
rect 227536 223796 227588 223848
rect 273168 223796 273220 223848
rect 671252 223796 671304 223848
rect 505192 223728 505244 223780
rect 507676 223728 507728 223780
rect 517704 223728 517756 223780
rect 617064 223728 617116 223780
rect 115296 223660 115348 223712
rect 188804 223660 188856 223712
rect 191564 223660 191616 223712
rect 194968 223660 195020 223712
rect 207664 223660 207716 223712
rect 228088 223660 228140 223712
rect 460572 223660 460624 223712
rect 463148 223660 463200 223712
rect 505376 223592 505428 223644
rect 614948 223592 615000 223644
rect 87972 223524 88024 223576
rect 164976 223524 165028 223576
rect 171784 223524 171836 223576
rect 181720 223524 181772 223576
rect 183192 223524 183244 223576
rect 184664 223524 184716 223576
rect 187332 223524 187384 223576
rect 242256 223524 242308 223576
rect 249432 223524 249484 223576
rect 276296 223524 276348 223576
rect 278596 223524 278648 223576
rect 315028 223524 315080 223576
rect 406752 223524 406804 223576
rect 414848 223524 414900 223576
rect 454868 223524 454920 223576
rect 460480 223524 460532 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 671160 223524 671212 223576
rect 562140 223456 562192 223508
rect 563336 223456 563388 223508
rect 88892 223388 88944 223440
rect 107660 223388 107712 223440
rect 108304 223388 108356 223440
rect 175924 223388 175976 223440
rect 184848 223388 184900 223440
rect 239680 223388 239732 223440
rect 244096 223388 244148 223440
rect 286048 223388 286100 223440
rect 81348 223252 81400 223304
rect 151912 223252 151964 223304
rect 68744 223116 68796 223168
rect 146484 223116 146536 223168
rect 146668 223116 146720 223168
rect 156420 223252 156472 223304
rect 156604 223252 156656 223304
rect 161940 223252 161992 223304
rect 162308 223252 162360 223304
rect 186872 223252 186924 223304
rect 188160 223252 188212 223304
rect 245108 223252 245160 223304
rect 250904 223252 250956 223304
rect 291200 223388 291252 223440
rect 316684 223388 316736 223440
rect 327264 223388 327316 223440
rect 517520 223388 517572 223440
rect 532516 223388 532568 223440
rect 534816 223388 534868 223440
rect 547420 223388 547472 223440
rect 671022 223388 671074 223440
rect 297548 223320 297600 223372
rect 305368 223320 305420 223372
rect 288992 223252 289044 223304
rect 295064 223252 295116 223304
rect 307668 223252 307720 223304
rect 335636 223252 335688 223304
rect 337936 223252 337988 223304
rect 359188 223252 359240 223304
rect 493048 223252 493100 223304
rect 508504 223252 508556 223304
rect 514668 223252 514720 223304
rect 535460 223252 535512 223304
rect 75828 222980 75880 223032
rect 154948 223116 155000 223168
rect 156420 223116 156472 223168
rect 176108 223116 176160 223168
rect 181996 223116 182048 223168
rect 240324 223116 240376 223168
rect 241336 223116 241388 223168
rect 283472 223116 283524 223168
rect 288256 223116 288308 223168
rect 321468 223116 321520 223168
rect 323952 223116 324004 223168
rect 348516 223116 348568 223168
rect 358544 223116 358596 223168
rect 374644 223116 374696 223168
rect 483112 223116 483164 223168
rect 496084 223116 496136 223168
rect 503352 223116 503404 223168
rect 521752 223116 521804 223168
rect 529480 223116 529532 223168
rect 555700 223116 555752 223168
rect 669044 223116 669096 223168
rect 152372 222980 152424 223032
rect 71412 222844 71464 222896
rect 151636 222844 151688 222896
rect 151774 222844 151826 222896
rect 156420 222844 156472 222896
rect 157524 222980 157576 223032
rect 219072 222980 219124 223032
rect 245292 222980 245344 223032
rect 289268 222980 289320 223032
rect 291660 222980 291712 223032
rect 300216 222980 300268 223032
rect 315672 222980 315724 223032
rect 344652 222980 344704 223032
rect 171784 222844 171836 222896
rect 172888 222844 172940 222896
rect 212632 222844 212684 222896
rect 213184 222844 213236 222896
rect 233332 222844 233384 222896
rect 234528 222844 234580 222896
rect 281540 222844 281592 222896
rect 282736 222844 282788 222896
rect 316316 222844 316368 222896
rect 321468 222844 321520 222896
rect 346584 222980 346636 223032
rect 349068 222980 349120 223032
rect 367192 222980 367244 223032
rect 368388 222980 368440 223032
rect 382648 222980 382700 223032
rect 383568 222980 383620 223032
rect 394884 222980 394936 223032
rect 486608 222980 486660 223032
rect 500408 222980 500460 223032
rect 508228 222980 508280 223032
rect 527180 222980 527232 223032
rect 532056 222980 532108 223032
rect 559012 222980 559064 223032
rect 345296 222844 345348 222896
rect 347872 222844 347924 222896
rect 85304 222708 85356 222760
rect 156604 222708 156656 222760
rect 156788 222708 156840 222760
rect 159824 222708 159876 222760
rect 165620 222708 165672 222760
rect 192024 222708 192076 222760
rect 193956 222708 194008 222760
rect 247408 222708 247460 222760
rect 284208 222708 284260 222760
rect 316960 222708 317012 222760
rect 347228 222708 347280 222760
rect 367836 222844 367888 222896
rect 375196 222844 375248 222896
rect 391020 222844 391072 222896
rect 395804 222844 395856 222896
rect 406476 222844 406528 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 479892 222844 479944 222896
rect 492036 222844 492088 222896
rect 500776 222844 500828 222896
rect 517520 222844 517572 222896
rect 519820 222844 519872 222896
rect 543280 222844 543332 222896
rect 554044 222844 554096 222896
rect 632704 222844 632756 222896
rect 558184 222708 558236 222760
rect 78588 222572 78640 222624
rect 88892 222572 88944 222624
rect 99288 222572 99340 222624
rect 107660 222572 107712 222624
rect 126520 222572 126572 222624
rect 108304 222436 108356 222488
rect 118424 222436 118476 222488
rect 191380 222572 191432 222624
rect 197176 222572 197228 222624
rect 249984 222572 250036 222624
rect 482744 222572 482796 222624
rect 593972 222572 594024 222624
rect 620284 222708 620336 222760
rect 126520 222300 126572 222352
rect 146668 222436 146720 222488
rect 139124 222300 139176 222352
rect 206836 222436 206888 222488
rect 207848 222436 207900 222488
rect 258356 222436 258408 222488
rect 502432 222436 502484 222488
rect 558184 222436 558236 222488
rect 558552 222436 558604 222488
rect 559840 222436 559892 222488
rect 627092 222572 627144 222624
rect 620284 222436 620336 222488
rect 630680 222436 630732 222488
rect 490012 222368 490064 222420
rect 147128 222300 147180 222352
rect 211988 222300 212040 222352
rect 237012 222300 237064 222352
rect 280896 222300 280948 222352
rect 484584 222300 484636 222352
rect 629852 222300 629904 222352
rect 502432 222164 502484 222216
rect 532516 222164 532568 222216
rect 621204 222164 621256 222216
rect 111984 222096 112036 222148
rect 185860 222096 185912 222148
rect 200396 222096 200448 222148
rect 252928 222096 252980 222148
rect 258080 222096 258132 222148
rect 263876 222096 263928 222148
rect 270040 222096 270092 222148
rect 306380 222096 306432 222148
rect 310704 222096 310756 222148
rect 312636 222096 312688 222148
rect 331404 222096 331456 222148
rect 353944 222096 353996 222148
rect 452568 222096 452620 222148
rect 455604 222096 455656 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 527180 222028 527232 222080
rect 528192 222028 528244 222080
rect 91284 221960 91336 222012
rect 167184 221960 167236 222012
rect 167460 221960 167512 222012
rect 172704 221960 172756 222012
rect 94596 221824 94648 221876
rect 169852 221824 169904 221876
rect 97724 221688 97776 221740
rect 167460 221688 167512 221740
rect 167644 221688 167696 221740
rect 73896 221552 73948 221604
rect 82084 221552 82136 221604
rect 86316 221552 86368 221604
rect 161940 221552 161992 221604
rect 162124 221552 162176 221604
rect 167828 221552 167880 221604
rect 168196 221688 168248 221740
rect 226524 221960 226576 222012
rect 232136 221960 232188 222012
rect 234712 221960 234764 222012
rect 261024 221960 261076 222012
rect 301688 221960 301740 222012
rect 313188 221960 313240 222012
rect 340420 221960 340472 222012
rect 553952 222028 554004 222080
rect 596916 222028 596968 222080
rect 552940 221960 552992 222012
rect 424968 221892 425020 221944
rect 429200 221892 429252 221944
rect 174084 221824 174136 221876
rect 231952 221824 232004 221876
rect 233700 221824 233752 221876
rect 277952 221824 278004 221876
rect 280068 221824 280120 221876
rect 313740 221824 313792 221876
rect 318248 221824 318300 221876
rect 343824 221824 343876 221876
rect 353300 221824 353352 221876
rect 372712 221824 372764 221876
rect 174912 221688 174964 221740
rect 185768 221688 185820 221740
rect 243084 221688 243136 221740
rect 182640 221552 182692 221604
rect 232136 221552 232188 221604
rect 263140 221688 263192 221740
rect 263508 221688 263560 221740
rect 301044 221688 301096 221740
rect 303252 221688 303304 221740
rect 332600 221688 332652 221740
rect 344652 221688 344704 221740
rect 364524 221688 364576 221740
rect 370964 221688 371016 221740
rect 380348 221824 380400 221876
rect 492496 221824 492548 221876
rect 506848 221824 506900 221876
rect 522672 221824 522724 221876
rect 544016 221892 544068 221944
rect 544200 221824 544252 221876
rect 597100 221960 597152 222012
rect 605012 221960 605064 222012
rect 597284 221824 597336 221876
rect 597468 221824 597520 221876
rect 603172 221824 603224 221876
rect 380072 221688 380124 221740
rect 386512 221688 386564 221740
rect 484768 221688 484820 221740
rect 497832 221688 497884 221740
rect 501328 221688 501380 221740
rect 520188 221756 520240 221808
rect 524236 221688 524288 221740
rect 543694 221688 543746 221740
rect 543832 221688 543884 221740
rect 558092 221688 558144 221740
rect 59360 221416 59412 221468
rect 141332 221416 141384 221468
rect 147588 221416 147640 221468
rect 204904 221416 204956 221468
rect 205088 221416 205140 221468
rect 220176 221416 220228 221468
rect 221004 221416 221056 221468
rect 243728 221552 243780 221604
rect 283748 221552 283800 221604
rect 302424 221552 302476 221604
rect 334072 221552 334124 221604
rect 348792 221552 348844 221604
rect 370044 221552 370096 221604
rect 373724 221552 373776 221604
rect 384304 221552 384356 221604
rect 391020 221552 391072 221604
rect 400404 221552 400456 221604
rect 401324 221552 401376 221604
rect 405832 221552 405884 221604
rect 475844 221552 475896 221604
rect 486148 221552 486200 221604
rect 496268 221552 496320 221604
rect 513380 221552 513432 221604
rect 516968 221552 517020 221604
rect 527548 221552 527600 221604
rect 533988 221552 534040 221604
rect 560760 221756 560812 221808
rect 560944 221756 560996 221808
rect 562692 221756 562744 221808
rect 562876 221688 562928 221740
rect 563014 221688 563066 221740
rect 563152 221688 563204 221740
rect 609428 221688 609480 221740
rect 558644 221552 558696 221604
rect 605932 221552 605984 221604
rect 234068 221416 234120 221468
rect 276112 221416 276164 221468
rect 284024 221416 284076 221468
rect 320364 221416 320416 221468
rect 332600 221416 332652 221468
rect 357532 221416 357584 221468
rect 369492 221416 369544 221468
rect 384120 221416 384172 221468
rect 384396 221416 384448 221468
rect 395160 221416 395212 221468
rect 396816 221416 396868 221468
rect 407304 221416 407356 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 468944 221416 468996 221468
rect 476212 221416 476264 221468
rect 483756 221416 483808 221468
rect 538772 221416 538824 221468
rect 538956 221416 539008 221468
rect 543096 221416 543148 221468
rect 544016 221416 544068 221468
rect 597100 221416 597152 221468
rect 543280 221348 543332 221400
rect 543832 221348 543884 221400
rect 597284 221348 597336 221400
rect 606116 221348 606168 221400
rect 104532 221280 104584 221332
rect 176476 221280 176528 221332
rect 111156 221144 111208 221196
rect 167644 221144 167696 221196
rect 167828 221144 167880 221196
rect 185860 221280 185912 221332
rect 234252 221280 234304 221332
rect 237840 221280 237892 221332
rect 243728 221280 243780 221332
rect 266820 221280 266872 221332
rect 303804 221280 303856 221332
rect 177304 221144 177356 221196
rect 185308 221144 185360 221196
rect 523500 221212 523552 221264
rect 601700 221212 601752 221264
rect 124404 221008 124456 221060
rect 193312 221008 193364 221060
rect 204904 221144 204956 221196
rect 211344 221144 211396 221196
rect 211528 221144 211580 221196
rect 260840 221144 260892 221196
rect 517520 221076 517572 221128
rect 518440 221076 518492 221128
rect 600596 221076 600648 221128
rect 205088 221008 205140 221060
rect 218152 221008 218204 221060
rect 221004 221008 221056 221060
rect 223488 221008 223540 221060
rect 268200 221008 268252 221060
rect 83004 220940 83056 220992
rect 521016 220940 521068 220992
rect 601332 220940 601384 220992
rect 151084 220872 151136 220924
rect 155040 220872 155092 220924
rect 162124 220872 162176 220924
rect 163780 220872 163832 220924
rect 80520 220804 80572 220856
rect 86132 220804 86184 220856
rect 167092 220872 167144 220924
rect 222292 220872 222344 220924
rect 227904 220872 227956 220924
rect 234068 220872 234120 220924
rect 253848 220872 253900 220924
rect 258632 220872 258684 220924
rect 101220 220736 101272 220788
rect 166448 220736 166500 220788
rect 418344 220804 418396 220856
rect 424048 220804 424100 220856
rect 456708 220804 456760 220856
rect 462136 220804 462188 220856
rect 466092 220804 466144 220856
rect 471336 220804 471388 220856
rect 515772 220804 515824 220856
rect 600320 220804 600372 220856
rect 76380 220600 76432 220652
rect 156144 220600 156196 220652
rect 156604 220600 156656 220652
rect 166448 220600 166500 220652
rect 167184 220736 167236 220788
rect 176476 220736 176528 220788
rect 176614 220736 176666 220788
rect 180524 220736 180576 220788
rect 180708 220736 180760 220788
rect 236736 220736 236788 220788
rect 254400 220736 254452 220788
rect 296812 220736 296864 220788
rect 340052 220736 340104 220788
rect 342352 220736 342404 220788
rect 414204 220736 414256 220788
rect 418160 220736 418212 220788
rect 431960 220736 432012 220788
rect 434812 220736 434864 220788
rect 474004 220736 474056 220788
rect 475384 220736 475436 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 500224 220736 500276 220788
rect 511816 220736 511868 220788
rect 455328 220668 455380 220720
rect 458824 220668 458876 220720
rect 465724 220668 465776 220720
rect 469588 220668 469640 220720
rect 543832 220668 543884 220720
rect 549076 220668 549128 220720
rect 550640 220668 550692 220720
rect 550824 220668 550876 220720
rect 221280 220600 221332 220652
rect 79692 220464 79744 220516
rect 151728 220464 151780 220516
rect 151912 220464 151964 220516
rect 153568 220464 153620 220516
rect 154212 220464 154264 220516
rect 156788 220464 156840 220516
rect 156972 220464 157024 220516
rect 158904 220464 158956 220516
rect 160836 220464 160888 220516
rect 163780 220464 163832 220516
rect 164148 220464 164200 220516
rect 166908 220464 166960 220516
rect 167092 220464 167144 220516
rect 223764 220600 223816 220652
rect 236184 220600 236236 220652
rect 246488 220600 246540 220652
rect 246948 220600 247000 220652
rect 288624 220600 288676 220652
rect 304908 220600 304960 220652
rect 333244 220600 333296 220652
rect 509884 220600 509936 220652
rect 522580 220600 522632 220652
rect 529020 220600 529072 220652
rect 601516 220736 601568 220788
rect 545028 220532 545080 220584
rect 223764 220464 223816 220516
rect 270592 220464 270644 220516
rect 276756 220464 276808 220516
rect 311348 220464 311400 220516
rect 328092 220464 328144 220516
rect 351276 220464 351328 220516
rect 364524 220464 364576 220516
rect 379704 220464 379756 220516
rect 469128 220464 469180 220516
rect 474556 220464 474608 220516
rect 488448 220464 488500 220516
rect 501880 220464 501932 220516
rect 511632 220464 511684 220516
rect 531688 220464 531740 220516
rect 548340 220464 548392 220516
rect 552848 220464 552900 220516
rect 560576 220464 560628 220516
rect 562876 220464 562928 220516
rect 607312 220600 607364 220652
rect 64604 220328 64656 220380
rect 141976 220328 142028 220380
rect 151774 220328 151826 220380
rect 202420 220328 202472 220380
rect 202788 220328 202840 220380
rect 214564 220328 214616 220380
rect 73068 220192 73120 220244
rect 151084 220260 151136 220312
rect 142344 220124 142396 220176
rect 156604 220192 156656 220244
rect 156788 220192 156840 220244
rect 212908 220192 212960 220244
rect 213828 220192 213880 220244
rect 262404 220328 262456 220380
rect 262680 220328 262732 220380
rect 264244 220328 264296 220380
rect 264612 220328 264664 220380
rect 269304 220328 269356 220380
rect 273444 220328 273496 220380
rect 309232 220328 309284 220380
rect 316500 220328 316552 220380
rect 342904 220328 342956 220380
rect 351276 220328 351328 220380
rect 369308 220328 369360 220380
rect 376944 220328 376996 220380
rect 388444 220328 388496 220380
rect 473176 220328 473228 220380
rect 481180 220328 481232 220380
rect 496452 220328 496504 220380
rect 509332 220328 509384 220380
rect 515404 220328 515456 220380
rect 530032 220328 530084 220380
rect 531136 220328 531188 220380
rect 553400 220328 553452 220380
rect 553952 220328 554004 220380
rect 601148 220464 601200 220516
rect 611452 220464 611504 220516
rect 217140 220192 217192 220244
rect 265164 220192 265216 220244
rect 267648 220192 267700 220244
rect 306840 220192 306892 220244
rect 309048 220192 309100 220244
rect 339684 220192 339736 220244
rect 342996 220192 343048 220244
rect 363328 220192 363380 220244
rect 363696 220192 363748 220244
rect 381084 220192 381136 220244
rect 388444 220192 388496 220244
rect 400956 220192 401008 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 472992 220192 473044 220244
rect 482008 220192 482060 220244
rect 482928 220192 482980 220244
rect 495348 220192 495400 220244
rect 497648 220192 497700 220244
rect 515220 220192 515272 220244
rect 528376 220192 528428 220244
rect 553584 220192 553636 220244
rect 566464 220328 566516 220380
rect 566648 220328 566700 220380
rect 567292 220328 567344 220380
rect 568396 220328 568448 220380
rect 568580 220328 568632 220380
rect 569776 220328 569828 220380
rect 569960 220328 570012 220380
rect 572444 220328 572496 220380
rect 572996 220328 573048 220380
rect 610072 220328 610124 220380
rect 563520 220192 563572 220244
rect 572628 220192 572680 220244
rect 572812 220192 572864 220244
rect 610256 220192 610308 220244
rect 69756 220056 69808 220108
rect 142160 220056 142212 220108
rect 151452 220056 151504 220108
rect 214288 220056 214340 220108
rect 214564 220056 214616 220108
rect 229284 220056 229336 220108
rect 230204 220056 230256 220108
rect 275284 220056 275336 220108
rect 292488 220056 292540 220108
rect 326160 220056 326212 220108
rect 328920 220056 328972 220108
rect 354772 220056 354824 220108
rect 355416 220056 355468 220108
rect 375564 220056 375616 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404728 220056 404780 220108
rect 421656 220056 421708 220108
rect 426716 220056 426768 220108
rect 478328 220056 478380 220108
rect 489460 220056 489512 220108
rect 489644 220056 489696 220108
rect 504364 220056 504416 220108
rect 513104 220056 513156 220108
rect 534172 220056 534224 220108
rect 538128 220056 538180 220108
rect 586520 220056 586572 220108
rect 633440 220056 633492 220108
rect 107844 219920 107896 219972
rect 127624 219920 127676 219972
rect 127808 219920 127860 219972
rect 185768 219920 185820 219972
rect 114468 219784 114520 219836
rect 185124 219784 185176 219836
rect 190092 219784 190144 219836
rect 190644 219920 190696 219972
rect 244464 219920 244516 219972
rect 253572 219920 253624 219972
rect 293316 219920 293368 219972
rect 586336 219988 586388 220040
rect 530032 219852 530084 219904
rect 560208 219852 560260 219904
rect 608692 219852 608744 219904
rect 202788 219784 202840 219836
rect 121092 219648 121144 219700
rect 127624 219648 127676 219700
rect 140780 219648 140832 219700
rect 140964 219648 141016 219700
rect 127808 219512 127860 219564
rect 134340 219512 134392 219564
rect 200764 219512 200816 219564
rect 201132 219648 201184 219700
rect 252744 219784 252796 219836
rect 270776 219784 270828 219836
rect 279148 219784 279200 219836
rect 286692 219784 286744 219836
rect 319076 219784 319128 219836
rect 506020 219716 506072 219768
rect 589280 219716 589332 219768
rect 589648 219716 589700 219768
rect 600780 219716 600832 219768
rect 600964 219716 601016 219768
rect 620468 219852 620520 219904
rect 203156 219648 203208 219700
rect 205824 219512 205876 219564
rect 207204 219648 207256 219700
rect 257252 219648 257304 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 527548 219580 527600 219632
rect 619916 219580 619968 219632
rect 208584 219512 208636 219564
rect 212908 219512 212960 219564
rect 215944 219512 215996 219564
rect 289820 219512 289872 219564
rect 105820 219444 105872 219496
rect 63960 219376 64012 219428
rect 64880 219376 64932 219428
rect 221648 219444 221700 219496
rect 147128 219376 147180 219428
rect 159180 219376 159232 219428
rect 160008 219376 160060 219428
rect 163320 219376 163372 219428
rect 163964 219376 164016 219428
rect 63132 219104 63184 219156
rect 106924 219240 106976 219292
rect 113640 219240 113692 219292
rect 156328 219240 156380 219292
rect 160008 219240 160060 219292
rect 204536 219376 204588 219428
rect 209688 219376 209740 219428
rect 210424 219376 210476 219428
rect 217968 219376 218020 219428
rect 167460 219240 167512 219292
rect 168196 219240 168248 219292
rect 169116 219240 169168 219292
rect 169668 219240 169720 219292
rect 169944 219240 169996 219292
rect 171048 219240 171100 219292
rect 172428 219240 172480 219292
rect 173164 219240 173216 219292
rect 182364 219240 182416 219292
rect 189724 219240 189776 219292
rect 192300 219240 192352 219292
rect 192944 219240 192996 219292
rect 193128 219240 193180 219292
rect 198188 219240 198240 219292
rect 198924 219240 198976 219292
rect 200028 219240 200080 219292
rect 201868 219240 201920 219292
rect 207664 219240 207716 219292
rect 211344 219240 211396 219292
rect 218152 219240 218204 219292
rect 258080 219376 258132 219428
rect 272892 219376 272944 219428
rect 366732 219512 366784 219564
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 223488 219240 223540 219292
rect 239496 219240 239548 219292
rect 272708 219240 272760 219292
rect 70584 219104 70636 219156
rect 117964 219104 118016 219156
rect 132592 219104 132644 219156
rect 177488 219104 177540 219156
rect 179052 219104 179104 219156
rect 196624 219104 196676 219156
rect 199752 219104 199804 219156
rect 243544 219104 243596 219156
rect 272340 219104 272392 219156
rect 289820 219240 289872 219292
rect 297548 219376 297600 219428
rect 304080 219376 304132 219428
rect 308404 219376 308456 219428
rect 320640 219376 320692 219428
rect 279056 219104 279108 219156
rect 286324 219104 286376 219156
rect 292028 219240 292080 219292
rect 313924 219240 313976 219292
rect 341340 219376 341392 219428
rect 342260 219376 342312 219428
rect 343824 219376 343876 219428
rect 347044 219376 347096 219428
rect 366180 219376 366232 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 428280 219376 428332 219428
rect 432144 219512 432196 219564
rect 501144 219512 501196 219564
rect 561680 219308 561732 219360
rect 562324 219308 562376 219360
rect 566924 219308 566976 219360
rect 567108 219308 567160 219360
rect 571892 219308 571944 219360
rect 572260 219308 572312 219360
rect 589464 219444 589516 219496
rect 600964 219444 601016 219496
rect 601516 219444 601568 219496
rect 607496 219444 607548 219496
rect 345296 219240 345348 219292
rect 419172 219240 419224 219292
rect 422668 219240 422720 219292
rect 557816 219240 557868 219292
rect 62304 218968 62356 219020
rect 72424 218968 72476 219020
rect 77208 218968 77260 219020
rect 140044 218968 140096 219020
rect 50712 218832 50764 218884
rect 62764 218832 62816 218884
rect 83832 218832 83884 218884
rect 153844 218968 153896 219020
rect 59820 218696 59872 218748
rect 143724 218832 143776 218884
rect 146760 218832 146812 218884
rect 142620 218696 142672 218748
rect 143264 218696 143316 218748
rect 144276 218696 144328 218748
rect 144828 218696 144880 218748
rect 145104 218696 145156 218748
rect 145932 218696 145984 218748
rect 148416 218696 148468 218748
rect 148968 218696 149020 218748
rect 149244 218696 149296 218748
rect 150072 218696 150124 218748
rect 153384 218832 153436 218884
rect 203524 218968 203576 219020
rect 206376 218968 206428 219020
rect 253848 218968 253900 219020
rect 259184 218968 259236 219020
rect 291660 218968 291712 219020
rect 295800 219104 295852 219156
rect 296720 219104 296772 219156
rect 300492 219104 300544 219156
rect 322112 219104 322164 219156
rect 325332 219104 325384 219156
rect 327724 219104 327776 219156
rect 340512 219104 340564 219156
rect 352564 219104 352616 219156
rect 362040 219104 362092 219156
rect 370964 219104 371016 219156
rect 552664 219104 552716 219156
rect 297364 218968 297416 219020
rect 307392 218968 307444 219020
rect 331864 218968 331916 219020
rect 333704 218968 333756 219020
rect 355232 218968 355284 219020
rect 357072 218968 357124 219020
rect 369124 218968 369176 219020
rect 370320 218968 370372 219020
rect 380072 218968 380124 219020
rect 380256 218968 380308 219020
rect 388628 218968 388680 219020
rect 547420 218968 547472 219020
rect 557632 218968 557684 219020
rect 567108 218968 567160 219020
rect 156328 218832 156380 218884
rect 162308 218832 162360 218884
rect 162492 218832 162544 218884
rect 171600 218832 171652 218884
rect 100392 218560 100444 218612
rect 105820 218560 105872 218612
rect 120264 218560 120316 218612
rect 165804 218696 165856 218748
rect 180064 218832 180116 218884
rect 175740 218696 175792 218748
rect 181168 218696 181220 218748
rect 184388 218696 184440 218748
rect 188988 218832 189040 218884
rect 194140 218832 194192 218884
rect 194324 218832 194376 218884
rect 239312 218832 239364 218884
rect 246120 218832 246172 218884
rect 279056 218832 279108 218884
rect 279240 218832 279292 218884
rect 189632 218696 189684 218748
rect 189816 218696 189868 218748
rect 195428 218696 195480 218748
rect 195612 218696 195664 218748
rect 198004 218696 198056 218748
rect 198188 218696 198240 218748
rect 246304 218696 246356 218748
rect 252744 218696 252796 218748
rect 107016 218424 107068 218476
rect 152372 218424 152424 218476
rect 152556 218424 152608 218476
rect 153108 218424 153160 218476
rect 156696 218424 156748 218476
rect 157248 218424 157300 218476
rect 171048 218560 171100 218612
rect 171600 218560 171652 218612
rect 181352 218560 181404 218612
rect 186504 218560 186556 218612
rect 194324 218560 194376 218612
rect 198096 218560 198148 218612
rect 200396 218560 200448 218612
rect 203064 218560 203116 218612
rect 206192 218560 206244 218612
rect 208032 218560 208084 218612
rect 211528 218560 211580 218612
rect 165620 218424 165672 218476
rect 166632 218424 166684 218476
rect 201868 218424 201920 218476
rect 217324 218560 217376 218612
rect 219624 218560 219676 218612
rect 264612 218560 264664 218612
rect 265992 218560 266044 218612
rect 272340 218560 272392 218612
rect 272708 218560 272760 218612
rect 279424 218560 279476 218612
rect 117964 218288 118016 218340
rect 123484 218288 123536 218340
rect 131856 218288 131908 218340
rect 132408 218288 132460 218340
rect 136824 218288 136876 218340
rect 139492 218288 139544 218340
rect 140136 218288 140188 218340
rect 181168 218288 181220 218340
rect 181536 218288 181588 218340
rect 181996 218288 182048 218340
rect 184020 218288 184072 218340
rect 184940 218288 184992 218340
rect 185676 218288 185728 218340
rect 186136 218288 186188 218340
rect 196440 218288 196492 218340
rect 213000 218424 213052 218476
rect 221648 218424 221700 218476
rect 225972 218424 226024 218476
rect 267004 218424 267056 218476
rect 285864 218832 285916 218884
rect 292028 218832 292080 218884
rect 314016 218832 314068 218884
rect 340052 218832 340104 218884
rect 347044 218832 347096 218884
rect 363512 218832 363564 218884
rect 368664 218832 368716 218884
rect 378784 218832 378836 218884
rect 382740 218832 382792 218884
rect 383568 218832 383620 218884
rect 386880 218832 386932 218884
rect 398104 218832 398156 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412548 218832 412600 218884
rect 291660 218696 291712 218748
rect 324596 218696 324648 218748
rect 327264 218696 327316 218748
rect 351092 218696 351144 218748
rect 353760 218696 353812 218748
rect 371792 218696 371844 218748
rect 383568 218696 383620 218748
rect 396264 218696 396316 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 471336 218696 471388 218748
rect 472900 218696 472952 218748
rect 482744 218696 482796 218748
rect 485320 218696 485372 218748
rect 542820 218696 542872 218748
rect 304264 218560 304316 218612
rect 398472 218560 398524 218612
rect 407764 218560 407816 218612
rect 429936 218560 429988 218612
rect 432144 218560 432196 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 537484 218560 537536 218612
rect 558000 218832 558052 218884
rect 548524 218696 548576 218748
rect 566740 218832 566792 218884
rect 567476 219104 567528 219156
rect 574284 219104 574336 219156
rect 567660 218968 567712 219020
rect 575480 218968 575532 219020
rect 288992 218424 289044 218476
rect 294144 218424 294196 218476
rect 316684 218424 316736 218476
rect 512736 218424 512788 218476
rect 542820 218424 542872 218476
rect 545028 218560 545080 218612
rect 557816 218560 557868 218612
rect 558000 218560 558052 218612
rect 560208 218560 560260 218612
rect 567476 218560 567528 218612
rect 567660 218424 567712 218476
rect 568304 218832 568356 218884
rect 572076 218832 572128 218884
rect 572536 218832 572588 218884
rect 572720 218832 572772 218884
rect 574468 218832 574520 218884
rect 596824 219308 596876 219360
rect 589280 219172 589332 219224
rect 597928 219172 597980 219224
rect 626356 218832 626408 218884
rect 568488 218696 568540 218748
rect 572260 218696 572312 218748
rect 601884 218696 601936 218748
rect 598756 218560 598808 218612
rect 604460 218424 604512 218476
rect 458180 218356 458232 218408
rect 202236 218288 202288 218340
rect 202788 218288 202840 218340
rect 204720 218288 204772 218340
rect 207848 218288 207900 218340
rect 208860 218288 208912 218340
rect 209504 218288 209556 218340
rect 210332 218288 210384 218340
rect 213184 218288 213236 218340
rect 222936 218288 222988 218340
rect 231032 218288 231084 218340
rect 232872 218288 232924 218340
rect 270776 218288 270828 218340
rect 426624 218288 426676 218340
rect 429384 218288 429436 218340
rect 434904 218288 434956 218340
rect 436652 218288 436704 218340
rect 450728 218288 450780 218340
rect 453856 218288 453908 218340
rect 461308 218288 461360 218340
rect 500408 218288 500460 218340
rect 609888 218288 609940 218340
rect 55680 218152 55732 218204
rect 56508 218152 56560 218204
rect 57428 218152 57480 218204
rect 61660 218152 61712 218204
rect 67272 218152 67324 218204
rect 68284 218152 68336 218204
rect 75552 218152 75604 218204
rect 76564 218152 76616 218204
rect 123576 218152 123628 218204
rect 165988 218152 166040 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58164 218016 58216 218068
rect 59360 218016 59412 218068
rect 61476 218016 61528 218068
rect 62028 218016 62080 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 66444 218016 66496 218068
rect 67548 218016 67600 218068
rect 68100 218016 68152 218068
rect 68744 218016 68796 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 83464 218016 83516 218068
rect 84660 218016 84712 218068
rect 85304 218016 85356 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 90456 218016 90508 218068
rect 91744 218016 91796 218068
rect 92940 218016 92992 218068
rect 93768 218016 93820 218068
rect 95424 218016 95476 218068
rect 96252 218016 96304 218068
rect 97080 218016 97132 218068
rect 98000 218016 98052 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 102876 218016 102928 218068
rect 103428 218016 103480 218068
rect 105360 218016 105412 218068
rect 106004 218016 106056 218068
rect 109500 218016 109552 218068
rect 110144 218016 110196 218068
rect 116124 218016 116176 218068
rect 117228 218016 117280 218068
rect 117780 218016 117832 218068
rect 118700 218016 118752 218068
rect 119436 218016 119488 218068
rect 119988 218016 120040 218068
rect 121920 218016 121972 218068
rect 122564 218016 122616 218068
rect 126060 218016 126112 218068
rect 126704 218016 126756 218068
rect 127716 218016 127768 218068
rect 128268 218016 128320 218068
rect 128544 218016 128596 218068
rect 129372 218016 129424 218068
rect 130200 218016 130252 218068
rect 132500 218016 132552 218068
rect 132684 218016 132736 218068
rect 133512 218016 133564 218068
rect 135996 218016 136048 218068
rect 136548 218016 136600 218068
rect 138480 218016 138532 218068
rect 139124 218016 139176 218068
rect 139492 218016 139544 218068
rect 171416 218152 171468 218204
rect 173256 218152 173308 218204
rect 170772 218016 170824 218068
rect 176476 218016 176528 218068
rect 178224 218016 178276 218068
rect 179328 218016 179380 218068
rect 179880 218152 179932 218204
rect 225604 218152 225656 218204
rect 241980 218152 242032 218204
rect 242900 218152 242952 218204
rect 243544 218152 243596 218204
rect 249064 218152 249116 218204
rect 297456 218152 297508 218204
rect 302884 218152 302936 218204
rect 335544 218152 335596 218204
rect 338672 218152 338724 218204
rect 358728 218152 358780 218204
rect 359464 218152 359516 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 400956 218152 401008 218204
rect 402244 218152 402296 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 427912 218152 427964 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 502984 218152 503036 218204
rect 548524 218152 548576 218204
rect 553400 218152 553452 218204
rect 556528 218152 556580 218204
rect 557632 218152 557684 218204
rect 560208 218152 560260 218204
rect 562140 218152 562192 218204
rect 563060 218152 563112 218204
rect 572444 218152 572496 218204
rect 614488 218152 614540 218204
rect 210332 218016 210384 218068
rect 210516 218016 210568 218068
rect 210976 218016 211028 218068
rect 214656 218016 214708 218068
rect 215208 218016 215260 218068
rect 215484 218016 215536 218068
rect 216128 218016 216180 218068
rect 218796 218016 218848 218068
rect 219348 218016 219400 218068
rect 221280 218016 221332 218068
rect 221832 218016 221884 218068
rect 225420 218016 225472 218068
rect 226156 218016 226208 218068
rect 227076 218016 227128 218068
rect 227536 218016 227588 218068
rect 229560 218016 229612 218068
rect 230480 218016 230532 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 235356 218016 235408 218068
rect 235816 218016 235868 218068
rect 240324 218016 240376 218068
rect 241336 218016 241388 218068
rect 243636 218016 243688 218068
rect 244096 218016 244148 218068
rect 244464 218016 244516 218068
rect 245292 218016 245344 218068
rect 247776 218016 247828 218068
rect 248328 218016 248380 218068
rect 248604 218016 248656 218068
rect 249248 218016 249300 218068
rect 250260 218016 250312 218068
rect 250904 218016 250956 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 256056 218016 256108 218068
rect 256516 218016 256568 218068
rect 256884 218016 256936 218068
rect 257528 218016 257580 218068
rect 258540 218016 258592 218068
rect 259368 218016 259420 218068
rect 260196 218016 260248 218068
rect 260748 218016 260800 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 268476 218016 268528 218068
rect 268936 218016 268988 218068
rect 269304 218016 269356 218068
rect 270224 218016 270276 218068
rect 270960 218016 271012 218068
rect 272524 218016 272576 218068
rect 277584 218016 277636 218068
rect 278596 218016 278648 218068
rect 280896 218016 280948 218068
rect 281448 218016 281500 218068
rect 281724 218016 281776 218068
rect 282736 218016 282788 218068
rect 283380 218016 283432 218068
rect 284300 218016 284352 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288072 218016 288124 218068
rect 289176 218016 289228 218068
rect 289636 218016 289688 218068
rect 290004 218016 290056 218068
rect 291108 218016 291160 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 298284 218016 298336 218068
rect 299388 218016 299440 218068
rect 299940 218016 299992 218068
rect 300676 218016 300728 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 305736 218016 305788 218068
rect 306196 218016 306248 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 308220 218016 308272 218068
rect 308864 218016 308916 218068
rect 309876 218016 309928 218068
rect 310336 218016 310388 218068
rect 312360 218016 312412 218068
rect 312912 218016 312964 218068
rect 314844 218016 314896 218068
rect 315488 218016 315540 218068
rect 317328 218016 317380 218068
rect 317972 218016 318024 218068
rect 318984 218016 319036 218068
rect 320088 218016 320140 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 323124 218016 323176 218068
rect 323952 218016 324004 218068
rect 324780 218016 324832 218068
rect 325516 218016 325568 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 330576 218016 330628 218068
rect 331036 218016 331088 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335176 218016 335228 218068
rect 337200 218016 337252 218068
rect 337752 218016 337804 218068
rect 338856 218016 338908 218068
rect 339408 218016 339460 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 345480 218016 345532 218068
rect 347228 218016 347280 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 349620 218016 349672 218068
rect 350172 218016 350224 218068
rect 352104 218016 352156 218068
rect 353300 218016 353352 218068
rect 356244 218016 356296 218068
rect 357256 218016 357308 218068
rect 357900 218016 357952 218068
rect 358544 218016 358596 218068
rect 359556 218016 359608 218068
rect 360108 218016 360160 218068
rect 360384 218016 360436 218068
rect 361028 218016 361080 218068
rect 367836 218016 367888 218068
rect 368388 218016 368440 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373540 218016 373592 218068
rect 374460 218016 374512 218068
rect 375012 218016 375064 218068
rect 376116 218016 376168 218068
rect 376668 218016 376720 218068
rect 378600 218016 378652 218068
rect 379244 218016 379296 218068
rect 381084 218016 381136 218068
rect 382096 218016 382148 218068
rect 385224 218016 385276 218068
rect 386052 218016 386104 218068
rect 389364 218016 389416 218068
rect 390468 218016 390520 218068
rect 392676 218016 392728 218068
rect 393136 218016 393188 218068
rect 393504 218016 393556 218068
rect 394516 218016 394568 218068
rect 395160 218016 395212 218068
rect 395804 218016 395856 218068
rect 397644 218016 397696 218068
rect 401324 218016 401376 218068
rect 401784 218016 401836 218068
rect 402796 218016 402848 218068
rect 403440 218016 403492 218068
rect 403992 218016 404044 218068
rect 405096 218016 405148 218068
rect 405556 218016 405608 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 428464 218016 428516 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 435732 218016 435784 218068
rect 436284 218016 436336 218068
rect 436560 218016 436612 218068
rect 437480 218016 437532 218068
rect 438216 218016 438268 218068
rect 438860 218016 438912 218068
rect 439872 218016 439924 218068
rect 440332 218016 440384 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 455604 218016 455656 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 492036 218016 492088 218068
rect 505652 218016 505704 218068
rect 507676 218016 507728 218068
rect 615684 218016 615736 218068
rect 646596 218016 646648 218068
rect 653404 218016 653456 218068
rect 676220 218016 676272 218068
rect 676864 218016 676916 218068
rect 563520 217948 563572 218000
rect 572076 217948 572128 218000
rect 131028 217812 131080 217864
rect 197728 217812 197780 217864
rect 523040 217812 523092 217864
rect 524236 217812 524288 217864
rect 535460 217812 535512 217864
rect 536656 217812 536708 217864
rect 536840 217812 536892 217864
rect 116952 217676 117004 217728
rect 189264 217676 189316 217728
rect 525984 217676 526036 217728
rect 526536 217676 526588 217728
rect 535920 217676 535972 217728
rect 598204 217676 598256 217728
rect 598572 217812 598624 217864
rect 601516 217676 601568 217728
rect 602344 217676 602396 217728
rect 603356 217812 603408 217864
rect 613384 217812 613436 217864
rect 604000 217676 604052 217728
rect 604460 217676 604512 217728
rect 616880 217676 616932 217728
rect 103704 217540 103756 217592
rect 178408 217540 178460 217592
rect 530584 217540 530636 217592
rect 530952 217540 531004 217592
rect 536840 217540 536892 217592
rect 538220 217540 538272 217592
rect 539140 217540 539192 217592
rect 545764 217540 545816 217592
rect 600136 217540 600188 217592
rect 603448 217540 603500 217592
rect 675852 217540 675904 217592
rect 676680 217540 676732 217592
rect 93768 217404 93820 217456
rect 171232 217404 171284 217456
rect 526536 217404 526588 217456
rect 601516 217404 601568 217456
rect 601884 217404 601936 217456
rect 628288 217404 628340 217456
rect 92066 217200 92118 217252
rect 170312 217268 170364 217320
rect 533436 217268 533488 217320
rect 598572 217268 598624 217320
rect 598756 217268 598808 217320
rect 436100 217200 436152 217252
rect 437342 217200 437394 217252
rect 448520 217200 448572 217252
rect 449762 217200 449814 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 489920 217200 489972 217252
rect 491162 217200 491214 217252
rect 498200 217200 498252 217252
rect 499442 217200 499494 217252
rect 511034 217132 511086 217184
rect 562140 217132 562192 217184
rect 503168 217064 503220 217116
rect 503582 217064 503634 217116
rect 562508 217132 562560 217184
rect 562692 217132 562744 217184
rect 563060 217132 563112 217184
rect 599124 217132 599176 217184
rect 600136 217268 600188 217320
rect 606760 217268 606812 217320
rect 642180 217268 642232 217320
rect 658924 217268 658976 217320
rect 601332 217132 601384 217184
rect 601516 217132 601568 217184
rect 604552 217132 604604 217184
rect 608968 216996 609020 217048
rect 609888 216996 609940 217048
rect 614120 216996 614172 217048
rect 574100 216860 574152 216912
rect 597560 216860 597612 216912
rect 598204 216860 598256 216912
rect 600780 216860 600832 216912
rect 594800 216724 594852 216776
rect 612280 216860 612332 216912
rect 601332 216724 601384 216776
rect 623872 216724 623924 216776
rect 648252 216588 648304 216640
rect 656164 216588 656216 216640
rect 675944 215500 675996 215552
rect 677048 215500 677100 215552
rect 575480 214820 575532 214872
rect 622400 214820 622452 214872
rect 649724 214820 649776 214872
rect 657728 214820 657780 214872
rect 574284 214684 574336 214736
rect 616696 214684 616748 214736
rect 617064 214684 617116 214736
rect 617800 214684 617852 214736
rect 621020 214684 621072 214736
rect 621664 214684 621716 214736
rect 630036 214684 630088 214736
rect 632888 214684 632940 214736
rect 644572 214684 644624 214736
rect 654784 214684 654836 214736
rect 574468 214548 574520 214600
rect 625528 214548 625580 214600
rect 654876 214548 654928 214600
rect 664444 214548 664496 214600
rect 664812 214548 664864 214600
rect 665824 214548 665876 214600
rect 610072 214412 610124 214464
rect 610624 214412 610676 214464
rect 616696 214412 616748 214464
rect 624424 214412 624476 214464
rect 626356 214276 626408 214328
rect 628840 214276 628892 214328
rect 35808 213936 35860 213988
rect 41696 213936 41748 213988
rect 627460 213936 627512 213988
rect 629392 213936 629444 213988
rect 663156 213868 663208 213920
rect 663708 213868 663760 213920
rect 659568 213596 659620 213648
rect 665548 213596 665600 213648
rect 574100 213460 574152 213512
rect 594800 213460 594852 213512
rect 647148 213460 647200 213512
rect 649908 213460 649960 213512
rect 574652 213324 574704 213376
rect 612832 213324 612884 213376
rect 651104 213324 651156 213376
rect 657544 213324 657596 213376
rect 574836 213188 574888 213240
rect 616144 213188 616196 213240
rect 643836 213188 643888 213240
rect 650644 213188 650696 213240
rect 658188 212848 658240 212900
rect 659108 212848 659160 212900
rect 650460 212712 650512 212764
rect 651288 212712 651340 212764
rect 664260 212712 664312 212764
rect 665088 212712 665140 212764
rect 632704 212508 632756 212560
rect 634360 212508 634412 212560
rect 630680 212372 630732 212424
rect 631600 212372 631652 212424
rect 35808 211556 35860 211608
rect 39580 211556 39632 211608
rect 35624 211284 35676 211336
rect 41696 211284 41748 211336
rect 35440 211148 35492 211200
rect 41328 211148 41380 211200
rect 578516 211148 578568 211200
rect 580908 211148 580960 211200
rect 680360 211148 680412 211200
rect 683120 211148 683172 211200
rect 633440 211012 633492 211064
rect 633808 211012 633860 211064
rect 635556 210128 635608 210180
rect 636568 210128 636620 210180
rect 35808 209788 35860 209840
rect 40224 209788 40276 209840
rect 579528 209788 579580 209840
rect 582288 209788 582340 209840
rect 581644 208564 581696 208616
rect 632152 209516 632204 209568
rect 652024 209516 652076 209568
rect 667572 209040 667624 209092
rect 35808 208496 35860 208548
rect 40500 208496 40552 208548
rect 35624 208360 35676 208412
rect 40040 208360 40092 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 35808 207136 35860 207188
rect 40776 207136 40828 207188
rect 580908 206864 580960 206916
rect 589464 206864 589516 206916
rect 35808 205776 35860 205828
rect 40960 205776 41012 205828
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 582288 205504 582340 205556
rect 589464 205504 589516 205556
rect 35808 204552 35860 204604
rect 40408 204552 40460 204604
rect 35624 204280 35676 204332
rect 41696 204348 41748 204400
rect 42064 204348 42116 204400
rect 43352 204348 43404 204400
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 42432 190136 42484 190188
rect 42984 190136 43036 190188
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 42432 187620 42484 187672
rect 43168 187620 43220 187672
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 582380 168376 582432 168428
rect 589464 168376 589516 168428
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579988 167016 580040 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589648 166268 589700 166320
rect 579344 165180 579396 165232
rect 582380 165180 582432 165232
rect 668216 165180 668268 165232
rect 669596 165180 669648 165232
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 578240 163616 578292 163668
rect 579988 163616 580040 163668
rect 668216 163276 668268 163328
rect 669780 163276 669832 163328
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 675852 162800 675904 162852
rect 678244 162800 678296 162852
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 668216 160012 668268 160064
rect 670332 160012 670384 160064
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 158720 585836 158772
rect 589464 158720 589516 158772
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 668308 155116 668360 155168
rect 670792 155116 670844 155168
rect 578332 154640 578384 154692
rect 580540 154640 580592 154692
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580264 151784 580316 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 585784 150560 585836 150612
rect 585140 149064 585192 149116
rect 589464 149064 589516 149116
rect 668216 148724 668268 148776
rect 670148 148724 670200 148776
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 578884 146276 578936 146328
rect 585140 146276 585192 146328
rect 584772 144916 584824 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 585784 143556 585836 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 580448 140768 580500 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580264 140700 580316 140752
rect 583024 139408 583076 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579528 138660 579580 138712
rect 588544 138660 588596 138712
rect 579068 137300 579120 137352
rect 584772 137300 584824 137352
rect 584588 136620 584640 136672
rect 589464 136620 589516 136672
rect 668216 136212 668268 136264
rect 669964 136212 670016 136264
rect 580264 134512 580316 134564
rect 589464 134512 589516 134564
rect 585968 132472 586020 132524
rect 589464 132472 589516 132524
rect 581828 131248 581880 131300
rect 589464 131248 589516 131300
rect 578884 131112 578936 131164
rect 585784 131112 585836 131164
rect 668584 129684 668636 129736
rect 670792 129684 670844 129736
rect 583392 129140 583444 129192
rect 590384 129140 590436 129192
rect 579528 129004 579580 129056
rect 587164 129004 587216 129056
rect 587808 126964 587860 127016
rect 589464 126964 589516 127016
rect 578332 125604 578384 125656
rect 580448 125604 580500 125656
rect 675944 125264 675996 125316
rect 676588 125264 676640 125316
rect 579068 124856 579120 124908
rect 587808 124856 587860 124908
rect 578700 124108 578752 124160
rect 583024 124108 583076 124160
rect 675852 123360 675904 123412
rect 676404 123360 676456 123412
rect 584404 122816 584456 122868
rect 589464 122816 589516 122868
rect 578884 122136 578936 122188
rect 584588 122136 584640 122188
rect 580632 122000 580684 122052
rect 590108 122000 590160 122052
rect 587348 121456 587400 121508
rect 589280 121456 589332 121508
rect 583208 120708 583260 120760
rect 590568 120708 590620 120760
rect 578516 118532 578568 118584
rect 580264 118532 580316 118584
rect 579528 116900 579580 116952
rect 583392 116900 583444 116952
rect 675852 116492 675904 116544
rect 676864 116492 676916 116544
rect 585784 115948 585836 116000
rect 589464 115948 589516 116000
rect 584588 115200 584640 115252
rect 589648 115200 589700 115252
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 583024 113160 583076 113212
rect 589464 113160 589516 113212
rect 579528 112820 579580 112872
rect 585968 112820 586020 112872
rect 586152 112412 586204 112464
rect 590108 112412 590160 112464
rect 668216 111460 668268 111512
rect 670700 111460 670752 111512
rect 581644 110440 581696 110492
rect 589464 110440 589516 110492
rect 579344 110236 579396 110288
rect 581828 110236 581880 110288
rect 580448 109080 580500 109132
rect 589464 109080 589516 109132
rect 578332 108944 578384 108996
rect 580632 108944 580684 108996
rect 667940 108808 667992 108860
rect 669964 108808 670016 108860
rect 582288 107652 582340 107704
rect 589464 107652 589516 107704
rect 580264 106292 580316 106344
rect 589464 106292 589516 106344
rect 579344 105612 579396 105664
rect 582288 105612 582340 105664
rect 587164 104864 587216 104916
rect 589832 104864 589884 104916
rect 578516 103368 578568 103420
rect 588728 103368 588780 103420
rect 579160 102076 579212 102128
rect 584404 102076 584456 102128
rect 584404 100104 584456 100156
rect 589464 100104 589516 100156
rect 578608 99968 578660 100020
rect 587348 99968 587400 100020
rect 592684 99968 592736 100020
rect 667940 99968 667992 100020
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 579528 99220 579580 99272
rect 583208 99220 583260 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 624608 99016 624660 99068
rect 635004 99016 635056 99068
rect 625068 98880 625120 98932
rect 636292 98880 636344 98932
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 647148 98744 647200 98796
rect 661960 98744 662012 98796
rect 630496 98608 630548 98660
rect 646596 98608 646648 98660
rect 631416 98268 631468 98320
rect 642180 98268 642232 98320
rect 633624 98132 633676 98184
rect 640708 98132 640760 98184
rect 618720 97928 618772 97980
rect 625804 97928 625856 97980
rect 629760 97928 629812 97980
rect 645308 97996 645360 98048
rect 659200 97928 659252 97980
rect 664168 97928 664220 97980
rect 620192 97792 620244 97844
rect 626356 97792 626408 97844
rect 628288 97792 628340 97844
rect 631416 97792 631468 97844
rect 632704 97792 632756 97844
rect 647700 97792 647752 97844
rect 653956 97792 654008 97844
rect 654324 97792 654376 97844
rect 655428 97792 655480 97844
rect 631232 97656 631284 97708
rect 647332 97656 647384 97708
rect 651840 97656 651892 97708
rect 659568 97656 659620 97708
rect 659936 97792 659988 97844
rect 665364 97792 665416 97844
rect 662512 97656 662564 97708
rect 627552 97520 627604 97572
rect 633624 97520 633676 97572
rect 633808 97520 633860 97572
rect 637764 97520 637816 97572
rect 643008 97520 643060 97572
rect 658004 97520 658056 97572
rect 658188 97520 658240 97572
rect 663064 97520 663116 97572
rect 605472 97384 605524 97436
rect 611912 97384 611964 97436
rect 612648 97384 612700 97436
rect 620284 97384 620336 97436
rect 621664 97384 621716 97436
rect 629300 97384 629352 97436
rect 631968 97384 632020 97436
rect 648620 97384 648672 97436
rect 650368 97384 650420 97436
rect 658280 97384 658332 97436
rect 623136 97248 623188 97300
rect 632060 97248 632112 97300
rect 633256 97248 633308 97300
rect 650552 97248 650604 97300
rect 656808 97180 656860 97232
rect 661408 97180 661460 97232
rect 626080 97112 626132 97164
rect 633808 97112 633860 97164
rect 634176 97112 634228 97164
rect 649080 97112 649132 97164
rect 658004 97044 658056 97096
rect 659844 97044 659896 97096
rect 634728 96976 634780 97028
rect 647148 96976 647200 97028
rect 597652 96908 597704 96960
rect 598204 96908 598256 96960
rect 598940 96908 598992 96960
rect 599676 96908 599728 96960
rect 606208 96908 606260 96960
rect 607128 96908 607180 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 654784 96908 654836 96960
rect 655428 96908 655480 96960
rect 656716 96908 656768 96960
rect 660120 96908 660172 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 626816 96840 626868 96892
rect 639236 96840 639288 96892
rect 644296 96772 644348 96824
rect 658832 96772 658884 96824
rect 609152 96704 609204 96756
rect 609704 96704 609756 96756
rect 640064 96568 640116 96620
rect 645124 96568 645176 96620
rect 646412 96568 646464 96620
rect 652208 96568 652260 96620
rect 652576 96568 652628 96620
rect 664352 96568 664404 96620
rect 638592 96432 638644 96484
rect 641352 96432 641404 96484
rect 641536 96432 641588 96484
rect 648436 96432 648488 96484
rect 648896 96432 648948 96484
rect 664536 96432 664588 96484
rect 637580 96296 637632 96348
rect 660672 96296 660724 96348
rect 644940 96160 644992 96212
rect 648068 96160 648120 96212
rect 648436 96160 648488 96212
rect 663800 96160 663852 96212
rect 591304 96024 591356 96076
rect 602620 96024 602672 96076
rect 610624 96024 610676 96076
rect 621664 96024 621716 96076
rect 640524 96024 640576 96076
rect 645584 96024 645636 96076
rect 647516 96024 647568 96076
rect 663984 96024 664036 96076
rect 594064 95888 594116 95940
rect 668032 95888 668084 95940
rect 639052 95752 639104 95804
rect 648620 95752 648672 95804
rect 653312 95752 653364 95804
rect 665180 95752 665232 95804
rect 645124 95616 645176 95668
rect 652024 95616 652076 95668
rect 652392 95616 652444 95668
rect 656348 95616 656400 95668
rect 648068 95480 648120 95532
rect 656164 95480 656216 95532
rect 641352 95412 641404 95464
rect 643468 95412 643520 95464
rect 647884 95412 647936 95464
rect 578332 95140 578384 95192
rect 584588 95140 584640 95192
rect 620928 95140 620980 95192
rect 625436 95140 625488 95192
rect 647516 95276 647568 95328
rect 652392 95276 652444 95328
rect 647516 95140 647568 95192
rect 647148 95004 647200 95056
rect 650276 95140 650328 95192
rect 616512 94936 616564 94988
rect 624976 94936 625028 94988
rect 607680 94460 607732 94512
rect 620836 94460 620888 94512
rect 619548 93780 619600 93832
rect 626172 93780 626224 93832
rect 651288 93576 651340 93628
rect 654692 93576 654744 93628
rect 579252 93372 579304 93424
rect 586152 93372 586204 93424
rect 609704 93100 609756 93152
rect 618628 93100 618680 93152
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 647516 92420 647568 92472
rect 655428 92420 655480 92472
rect 606944 91740 606996 91792
rect 622400 91740 622452 91792
rect 578608 91128 578660 91180
rect 585784 91128 585836 91180
rect 618168 91128 618220 91180
rect 611268 90992 611320 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 648620 90788 648672 90840
rect 655428 90788 655480 90840
rect 620836 89632 620888 89684
rect 626448 89632 626500 89684
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 664168 88748 664220 88800
rect 656348 88612 656400 88664
rect 657452 88612 657504 88664
rect 579252 88272 579304 88324
rect 589924 88272 589976 88324
rect 622400 88272 622452 88324
rect 626448 88272 626500 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 618168 88136 618220 88188
rect 626264 88136 626316 88188
rect 648252 86980 648304 87032
rect 662512 86980 662564 87032
rect 578332 86912 578384 86964
rect 580448 86912 580500 86964
rect 656716 86844 656768 86896
rect 659568 86844 659620 86896
rect 656164 86708 656216 86760
rect 660672 86708 660724 86760
rect 652024 86572 652076 86624
rect 660120 86572 660172 86624
rect 652208 86436 652260 86488
rect 657176 86436 657228 86488
rect 621664 86300 621716 86352
rect 626448 86300 626500 86352
rect 647884 86300 647936 86352
rect 661408 86300 661460 86352
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 618628 85348 618680 85400
rect 625252 85348 625304 85400
rect 608508 84124 608560 84176
rect 626448 84124 626500 84176
rect 579252 83988 579304 84040
rect 581644 83988 581696 84040
rect 578884 82764 578936 82816
rect 583024 82764 583076 82816
rect 579252 82084 579304 82136
rect 587164 82084 587216 82136
rect 628748 81064 628800 81116
rect 642456 81064 642508 81116
rect 615408 80928 615460 80980
rect 646320 80928 646372 80980
rect 613844 80792 613896 80844
rect 647332 80792 647384 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 614028 79432 614080 79484
rect 646044 79432 646096 79484
rect 583024 79296 583076 79348
rect 600504 79296 600556 79348
rect 612648 79296 612700 79348
rect 648620 79296 648672 79348
rect 578240 78072 578292 78124
rect 580264 78072 580316 78124
rect 633440 78072 633492 78124
rect 645308 78072 645360 78124
rect 631048 77936 631100 77988
rect 643100 77936 643152 77988
rect 628472 77664 628524 77716
rect 632796 77664 632848 77716
rect 624424 77392 624476 77444
rect 628472 77392 628524 77444
rect 625804 77256 625856 77308
rect 631048 77256 631100 77308
rect 620284 76780 620336 76832
rect 648988 76780 649040 76832
rect 612004 76644 612056 76696
rect 662420 76644 662472 76696
rect 587164 76508 587216 76560
rect 668216 76508 668268 76560
rect 616788 75420 616840 75472
rect 646688 75420 646740 75472
rect 607128 75284 607180 75336
rect 646504 75284 646556 75336
rect 578884 75148 578936 75200
rect 666560 75148 666612 75200
rect 579528 73108 579580 73160
rect 588544 73108 588596 73160
rect 578516 71544 578568 71596
rect 584404 71544 584456 71596
rect 579528 66852 579580 66904
rect 625988 66852 626040 66904
rect 579528 64812 579580 64864
rect 592684 64812 592736 64864
rect 579528 62024 579580 62076
rect 587164 62024 587216 62076
rect 578332 59984 578384 60036
rect 624424 59984 624476 60036
rect 577504 58760 577556 58812
rect 604460 58760 604512 58812
rect 576124 58624 576176 58676
rect 603080 58624 603132 58676
rect 579528 57876 579580 57928
rect 594064 57876 594116 57928
rect 574928 57196 574980 57248
rect 600320 57196 600372 57248
rect 574744 55972 574796 56024
rect 598940 55972 598992 56024
rect 574468 55836 574520 55888
rect 601884 55836 601936 55888
rect 596456 55156 596508 55208
rect 597836 55020 597888 55072
rect 463332 53592 463384 53644
rect 463516 53592 463568 53644
rect 463884 53592 463936 53644
rect 464068 53592 464120 53644
rect 460388 53456 460440 53508
rect 597652 54884 597704 54936
rect 599124 54748 599176 54800
rect 623044 54612 623096 54664
rect 625804 54476 625856 54528
rect 596272 54340 596324 54392
rect 465908 53592 465960 53644
rect 470324 53592 470376 53644
rect 470968 53592 471020 53644
rect 471152 53592 471204 53644
rect 471704 53592 471756 53644
rect 471980 53592 472032 53644
rect 476764 53592 476816 53644
rect 583024 54204 583076 54256
rect 580448 54068 580500 54120
rect 574744 53932 574796 53984
rect 464988 53456 465040 53508
rect 479616 53592 479668 53644
rect 479984 53592 480036 53644
rect 480168 53592 480220 53644
rect 50528 53320 50580 53372
rect 130384 53320 130436 53372
rect 462228 53320 462280 53372
rect 574928 53796 574980 53848
rect 48964 53184 49016 53236
rect 129004 53184 129056 53236
rect 463148 53184 463200 53236
rect 479616 53184 479668 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 47584 53048 47636 53100
rect 129188 53048 129240 53100
rect 461308 53048 461360 53100
rect 480168 53048 480220 53100
rect 463332 52912 463384 52964
rect 463792 52912 463844 52964
rect 459146 52776 459198 52828
rect 465126 52776 465178 52828
rect 479984 52776 480036 52828
rect 471704 52640 471756 52692
rect 50344 51824 50396 51876
rect 129372 51824 129424 51876
rect 46204 51688 46256 51740
rect 130568 51688 130620 51740
rect 145380 51688 145432 51740
rect 306012 51688 306064 51740
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 49148 50328 49200 50380
rect 131028 50328 131080 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 51724 49104 51776 49156
rect 129648 49104 129700 49156
rect 45468 48968 45520 49020
rect 128820 48968 128872 49020
rect 128820 47812 128872 47864
rect 130752 47812 130804 47864
rect 625988 46452 626040 46504
rect 661776 46452 661828 46504
rect 129004 46044 129056 46096
rect 131764 46044 131816 46096
rect 130568 45908 130620 45960
rect 132500 45908 132552 45960
rect 129648 45364 129700 45416
rect 43812 45160 43864 45212
rect 131120 45160 131172 45212
rect 131396 45296 131448 45348
rect 132960 45296 133012 45348
rect 131396 45160 131448 45212
rect 133144 45160 133196 45212
rect 129372 45024 129424 45076
rect 131580 44752 131632 44804
rect 131764 44644 131816 44696
rect 131948 44616 132000 44668
rect 129188 44480 129240 44532
rect 43628 44276 43680 44328
rect 129096 44276 129148 44328
rect 130752 44276 130804 44328
rect 132500 44344 132552 44396
rect 43444 44140 43496 44192
rect 131580 44140 131632 44192
rect 132960 44252 133012 44304
rect 130384 44004 130436 44056
rect 133144 44140 133196 44192
rect 440240 43596 440292 43648
rect 441068 43596 441120 43648
rect 187332 42712 187384 42764
rect 431224 42712 431276 42764
rect 441068 42712 441120 42764
rect 449164 42712 449216 42764
rect 459560 42440 459612 42492
rect 460112 42440 460164 42492
rect 454500 42304 454552 42356
rect 463056 42304 463108 42356
rect 661408 42129 661460 42181
rect 431224 41964 431276 42016
rect 441068 41964 441120 42016
rect 449164 41964 449216 42016
rect 459376 41964 459428 42016
rect 404636 41828 404688 41880
rect 420736 41692 420788 41744
rect 427084 41692 427136 41744
rect 459192 41692 459244 41744
rect 311072 41556 311124 41608
rect 454500 41556 454552 41608
rect 420736 41420 420788 41472
rect 427084 41420 427136 41472
<< metal2 >>
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676036 897096
rect 676088 897087 676090 897096
rect 676036 897058 676088 897064
rect 652024 897048 652076 897054
rect 652024 896990 652076 896996
rect 651472 868896 651524 868902
rect 651472 868838 651524 868844
rect 651484 868601 651512 868838
rect 651470 868592 651526 868601
rect 651470 868527 651526 868536
rect 652036 867649 652064 896990
rect 675850 896744 675906 896753
rect 675850 896679 675906 896688
rect 675864 895830 675892 896679
rect 676034 896336 676090 896345
rect 676034 896271 676090 896280
rect 654784 895824 654836 895830
rect 654784 895766 654836 895772
rect 675852 895824 675904 895830
rect 675852 895766 675904 895772
rect 653404 880524 653456 880530
rect 653404 880466 653456 880472
rect 652022 867640 652078 867649
rect 652022 867575 652078 867584
rect 651472 866652 651524 866658
rect 651472 866594 651524 866600
rect 651484 866289 651512 866594
rect 651470 866280 651526 866289
rect 651470 866215 651526 866224
rect 653416 865230 653444 880466
rect 654796 868902 654824 895766
rect 676048 895694 676076 896271
rect 672724 895688 672776 895694
rect 672724 895630 672776 895636
rect 676036 895688 676088 895694
rect 676036 895630 676088 895636
rect 672540 894464 672592 894470
rect 672540 894406 672592 894412
rect 671988 893036 672040 893042
rect 671988 892978 672040 892984
rect 670884 892900 670936 892906
rect 670884 892842 670936 892848
rect 657544 869440 657596 869446
rect 657544 869382 657596 869388
rect 654784 868896 654836 868902
rect 654784 868838 654836 868844
rect 654140 868080 654192 868086
rect 654140 868022 654192 868028
rect 651380 865224 651432 865230
rect 651378 865192 651380 865201
rect 653404 865224 653456 865230
rect 651432 865192 651434 865201
rect 653404 865166 653456 865172
rect 651378 865127 651434 865136
rect 651472 863864 651524 863870
rect 651470 863832 651472 863841
rect 651524 863832 651526 863841
rect 651470 863767 651526 863776
rect 654152 862510 654180 868022
rect 657556 863870 657584 869382
rect 657544 863864 657596 863870
rect 657544 863806 657596 863812
rect 651472 862504 651524 862510
rect 651472 862446 651524 862452
rect 654140 862504 654192 862510
rect 654140 862446 654192 862452
rect 651484 862345 651512 862446
rect 651470 862336 651526 862345
rect 651470 862271 651526 862280
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35622 818000 35678 818009
rect 35622 817935 35678 817944
rect 35636 817154 35664 817935
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817154 35848 817255
rect 35624 817148 35676 817154
rect 35624 817090 35676 817096
rect 35808 817148 35860 817154
rect 35808 817090 35860 817096
rect 46204 817148 46256 817154
rect 46204 817090 46256 817096
rect 35622 816912 35678 816921
rect 35622 816847 35678 816856
rect 35636 815794 35664 816847
rect 35806 816096 35862 816105
rect 35806 816031 35862 816040
rect 35624 815788 35676 815794
rect 35624 815730 35676 815736
rect 35820 815658 35848 816031
rect 44824 815788 44876 815794
rect 44824 815730 44876 815736
rect 35808 815652 35860 815658
rect 35808 815594 35860 815600
rect 35622 815280 35678 815289
rect 35622 815215 35678 815224
rect 35636 814434 35664 815215
rect 35806 814464 35862 814473
rect 35624 814428 35676 814434
rect 35806 814399 35862 814408
rect 44272 814428 44324 814434
rect 35624 814370 35676 814376
rect 35820 814298 35848 814399
rect 44272 814370 44324 814376
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41326 813648 41382 813657
rect 41326 813583 41382 813592
rect 41340 812870 41368 813583
rect 41328 812864 41380 812870
rect 41142 812832 41198 812841
rect 41328 812806 41380 812812
rect 43260 812864 43312 812870
rect 43260 812806 43312 812812
rect 41142 812767 41198 812776
rect 40498 812424 40554 812433
rect 40498 812359 40554 812368
rect 39302 811608 39358 811617
rect 39302 811543 39358 811552
rect 33046 811200 33102 811209
rect 33046 811135 33102 811144
rect 31022 809976 31078 809985
rect 31022 809911 31078 809920
rect 31036 801106 31064 809911
rect 31758 806712 31814 806721
rect 31758 806647 31760 806656
rect 31812 806647 31814 806656
rect 31760 806618 31812 806624
rect 33060 802466 33088 811135
rect 33782 809568 33838 809577
rect 33782 809503 33838 809512
rect 33048 802460 33100 802466
rect 33048 802402 33100 802408
rect 33796 801242 33824 809503
rect 35624 806676 35676 806682
rect 35624 806618 35676 806624
rect 35636 802602 35664 806618
rect 35624 802596 35676 802602
rect 35624 802538 35676 802544
rect 33784 801236 33836 801242
rect 33784 801178 33836 801184
rect 31024 801100 31076 801106
rect 31024 801042 31076 801048
rect 39316 800902 39344 811543
rect 40512 805633 40540 812359
rect 41156 810762 41184 812767
rect 41786 810792 41842 810801
rect 41144 810756 41196 810762
rect 41144 810698 41196 810704
rect 41616 810750 41786 810778
rect 40682 809160 40738 809169
rect 40682 809095 40738 809104
rect 40498 805624 40554 805633
rect 40498 805559 40554 805568
rect 40132 801236 40184 801242
rect 40132 801178 40184 801184
rect 39304 800896 39356 800902
rect 40144 800873 40172 801178
rect 39304 800838 39356 800844
rect 40130 800864 40186 800873
rect 40130 800799 40186 800808
rect 40696 800601 40724 809095
rect 40958 808344 41014 808353
rect 40958 808279 41014 808288
rect 40972 807362 41000 808279
rect 41142 807936 41198 807945
rect 41142 807871 41198 807880
rect 41156 807498 41184 807871
rect 41144 807492 41196 807498
rect 41144 807434 41196 807440
rect 40960 807356 41012 807362
rect 40960 807298 41012 807304
rect 41326 806304 41382 806313
rect 41326 806239 41382 806248
rect 41340 806002 41368 806239
rect 41328 805996 41380 806002
rect 41328 805938 41380 805944
rect 41616 804681 41644 810750
rect 41786 810727 41842 810736
rect 42524 810756 42576 810762
rect 42524 810698 42576 810704
rect 41970 810384 42026 810393
rect 41970 810319 42026 810328
rect 41786 808752 41842 808761
rect 41786 808687 41842 808696
rect 41800 805225 41828 808687
rect 41786 805216 41842 805225
rect 41786 805151 41842 805160
rect 41984 804953 42012 810319
rect 41970 804944 42026 804953
rect 41970 804879 42026 804888
rect 41602 804672 41658 804681
rect 41602 804607 41658 804616
rect 42156 802460 42208 802466
rect 42156 802402 42208 802408
rect 42340 802460 42392 802466
rect 42340 802402 42392 802408
rect 42168 801530 42196 802402
rect 42352 802346 42380 802402
rect 42352 802318 42472 802346
rect 42168 801502 42288 801530
rect 41972 800896 42024 800902
rect 41972 800838 42024 800844
rect 40682 800592 40738 800601
rect 40682 800527 40738 800536
rect 41984 800329 42012 800838
rect 41970 800320 42026 800329
rect 41970 800255 42026 800264
rect 42260 799898 42288 801502
rect 42168 799870 42288 799898
rect 42168 799445 42196 799870
rect 42444 799490 42472 802318
rect 42260 799462 42472 799490
rect 42260 798266 42288 799462
rect 42536 799218 42564 810698
rect 42890 807528 42946 807537
rect 42890 807463 42946 807472
rect 43076 807492 43128 807498
rect 42182 798238 42288 798266
rect 42352 799190 42564 799218
rect 42352 797994 42380 799190
rect 42260 797966 42380 797994
rect 42260 797619 42288 797966
rect 42524 797700 42576 797706
rect 42524 797642 42576 797648
rect 42182 797591 42288 797619
rect 42154 797328 42210 797337
rect 42154 797263 42210 797272
rect 42168 796960 42196 797263
rect 41786 796240 41842 796249
rect 41786 796175 41842 796184
rect 41800 795765 41828 796175
rect 42536 795138 42564 797642
rect 42904 796770 42932 807463
rect 43076 807434 43128 807440
rect 43088 804554 43116 807434
rect 43088 804526 43208 804554
rect 42904 796742 43116 796770
rect 42892 796544 42944 796550
rect 42812 796492 42892 796498
rect 42812 796486 42944 796492
rect 42812 796470 42932 796486
rect 42812 795546 42840 796470
rect 43088 796226 43116 796742
rect 42182 795110 42564 795138
rect 42720 795518 42840 795546
rect 42904 796198 43116 796226
rect 42432 795048 42484 795054
rect 42432 794990 42484 794996
rect 42444 794594 42472 794990
rect 42182 794566 42472 794594
rect 41786 794472 41842 794481
rect 41786 794407 41842 794416
rect 41800 793900 41828 794407
rect 42432 794096 42484 794102
rect 42432 794038 42484 794044
rect 42444 793302 42472 794038
rect 42182 793274 42472 793302
rect 42062 792976 42118 792985
rect 42062 792911 42118 792920
rect 42076 792744 42104 792911
rect 42720 791738 42748 795518
rect 42444 791710 42748 791738
rect 42246 791344 42302 791353
rect 42246 791279 42302 791288
rect 41786 790664 41842 790673
rect 41786 790599 41842 790608
rect 41800 790228 41828 790599
rect 42260 789750 42288 791279
rect 42248 789744 42300 789750
rect 42248 789686 42300 789692
rect 42444 789630 42472 791710
rect 42614 791616 42670 791625
rect 42614 791551 42670 791560
rect 42182 789602 42472 789630
rect 42248 789540 42300 789546
rect 42248 789482 42300 789488
rect 42260 789290 42288 789482
rect 42168 789262 42288 789290
rect 42168 788936 42196 789262
rect 42628 788746 42656 791551
rect 42168 788718 42656 788746
rect 42168 788392 42196 788718
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 41786 786856 41842 786865
rect 41786 786791 41842 786800
rect 41800 786556 41828 786791
rect 41786 786176 41842 786185
rect 41786 786111 41842 786120
rect 41800 785944 41828 786111
rect 42260 785278 42288 788151
rect 42616 786684 42668 786690
rect 42616 786626 42668 786632
rect 42182 785250 42288 785278
rect 42628 784734 42656 786626
rect 42182 784706 42656 784734
rect 40498 776656 40554 776665
rect 40498 776591 40554 776600
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774752 35862 774761
rect 35806 774687 35862 774696
rect 35820 774246 35848 774687
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 35162 773936 35218 773945
rect 35162 773871 35218 773880
rect 35176 772886 35204 773871
rect 35346 773528 35402 773537
rect 35346 773463 35402 773472
rect 35360 773022 35388 773463
rect 40512 773430 40540 776591
rect 41696 774240 41748 774246
rect 42064 774240 42116 774246
rect 41748 774188 42064 774194
rect 41696 774182 42116 774188
rect 41708 774166 42104 774182
rect 35808 773424 35860 773430
rect 35808 773366 35860 773372
rect 40500 773424 40552 773430
rect 40500 773366 40552 773372
rect 35532 773152 35584 773158
rect 35530 773120 35532 773129
rect 35820 773129 35848 773366
rect 40500 773152 40552 773158
rect 35584 773120 35586 773129
rect 35530 773055 35586 773064
rect 35806 773120 35862 773129
rect 35806 773055 35862 773064
rect 40498 773120 40500 773129
rect 40552 773120 40554 773129
rect 40498 773055 40554 773064
rect 35348 773016 35400 773022
rect 35348 772958 35400 772964
rect 41696 773016 41748 773022
rect 42064 773016 42116 773022
rect 41748 772964 42064 772970
rect 41696 772958 42116 772964
rect 41708 772942 42104 772958
rect 35164 772880 35216 772886
rect 35164 772822 35216 772828
rect 41696 772744 41748 772750
rect 42064 772744 42116 772750
rect 41748 772692 42064 772698
rect 41696 772686 42116 772692
rect 41708 772670 42104 772686
rect 35622 772304 35678 772313
rect 35622 772239 35678 772248
rect 41326 772304 41382 772313
rect 41326 772239 41382 772248
rect 35636 771594 35664 772239
rect 35806 771896 35862 771905
rect 35806 771831 35808 771840
rect 35860 771831 35862 771840
rect 39580 771860 39632 771866
rect 35808 771802 35860 771808
rect 39580 771802 39632 771808
rect 35624 771588 35676 771594
rect 35624 771530 35676 771536
rect 39592 771497 39620 771802
rect 41340 771662 41368 772239
rect 41328 771656 41380 771662
rect 41328 771598 41380 771604
rect 42064 771520 42116 771526
rect 35806 771488 35862 771497
rect 35806 771423 35808 771432
rect 35860 771423 35862 771432
rect 39578 771488 39634 771497
rect 41708 771468 42064 771474
rect 41708 771462 42116 771468
rect 41708 771458 42104 771462
rect 39578 771423 39634 771432
rect 41696 771452 42104 771458
rect 35808 771394 35860 771400
rect 41748 771446 42104 771452
rect 41696 771394 41748 771400
rect 35622 771080 35678 771089
rect 35622 771015 35678 771024
rect 35636 770234 35664 771015
rect 35806 770672 35862 770681
rect 35806 770607 35862 770616
rect 40038 770672 40094 770681
rect 40038 770607 40094 770616
rect 35820 770506 35848 770607
rect 40052 770506 40080 770607
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 40040 770500 40092 770506
rect 40040 770442 40092 770448
rect 35806 770264 35862 770273
rect 35624 770228 35676 770234
rect 35806 770199 35862 770208
rect 40316 770228 40368 770234
rect 35624 770170 35676 770176
rect 35820 770098 35848 770199
rect 40316 770170 40368 770176
rect 35808 770092 35860 770098
rect 35808 770034 35860 770040
rect 35346 769448 35402 769457
rect 35346 769383 35402 769392
rect 35360 768738 35388 769383
rect 35530 769040 35586 769049
rect 35530 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35808 768984
rect 35544 768874 35572 768975
rect 35860 768975 35862 768984
rect 39764 769004 39816 769010
rect 35808 768946 35860 768952
rect 39764 768946 39816 768952
rect 35532 768868 35584 768874
rect 35532 768810 35584 768816
rect 35348 768732 35400 768738
rect 35348 768674 35400 768680
rect 39776 768641 39804 768946
rect 39762 768632 39818 768641
rect 39762 768567 39818 768576
rect 35622 768224 35678 768233
rect 35622 768159 35678 768168
rect 33046 767816 33102 767825
rect 33046 767751 33102 767760
rect 33060 761054 33088 767751
rect 35636 767378 35664 768159
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 35820 767514 35848 767751
rect 35808 767508 35860 767514
rect 35808 767450 35860 767456
rect 36544 767508 36596 767514
rect 36544 767450 36596 767456
rect 35624 767372 35676 767378
rect 35624 767314 35676 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 33048 761048 33100 761054
rect 33048 760990 33100 760996
rect 35176 759626 35204 766935
rect 35806 766592 35862 766601
rect 35806 766527 35862 766536
rect 35820 766086 35848 766527
rect 35808 766080 35860 766086
rect 35808 766022 35860 766028
rect 35806 765776 35862 765785
rect 35806 765711 35862 765720
rect 35820 764862 35848 765711
rect 35808 764856 35860 764862
rect 35808 764798 35860 764804
rect 35808 764584 35860 764590
rect 35806 764552 35808 764561
rect 35860 764552 35862 764561
rect 35806 764487 35862 764496
rect 35806 764144 35862 764153
rect 35806 764079 35862 764088
rect 35820 763298 35848 764079
rect 35808 763292 35860 763298
rect 35808 763234 35860 763240
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761938 35848 762855
rect 35808 761932 35860 761938
rect 35808 761874 35860 761880
rect 35164 759620 35216 759626
rect 35164 759562 35216 759568
rect 36556 759121 36584 767450
rect 40328 767009 40356 770170
rect 41708 770098 42104 770114
rect 41696 770092 42116 770098
rect 41748 770086 42064 770092
rect 41696 770034 41748 770040
rect 42064 770034 42116 770040
rect 40684 768868 40736 768874
rect 40684 768810 40736 768816
rect 40314 767000 40370 767009
rect 40314 766935 40370 766944
rect 39304 766080 39356 766086
rect 39304 766022 39356 766028
rect 39316 764561 39344 766022
rect 40408 764856 40460 764862
rect 40408 764798 40460 764804
rect 39302 764552 39358 764561
rect 39302 764487 39358 764496
rect 40420 764153 40448 764798
rect 40406 764144 40462 764153
rect 40406 764079 40462 764088
rect 37094 763736 37150 763745
rect 37094 763671 37096 763680
rect 37148 763671 37150 763680
rect 39304 763700 39356 763706
rect 37096 763642 37148 763648
rect 39304 763642 39356 763648
rect 36542 759112 36598 759121
rect 36542 759047 36598 759056
rect 39316 757790 39344 763642
rect 39948 761932 40000 761938
rect 39948 761874 40000 761880
rect 39304 757784 39356 757790
rect 39304 757726 39356 757732
rect 39960 757489 39988 761874
rect 40500 759552 40552 759558
rect 40498 759520 40500 759529
rect 40552 759520 40554 759529
rect 40498 759455 40554 759464
rect 40696 757761 40724 768810
rect 41696 768732 41748 768738
rect 41696 768674 41748 768680
rect 41708 768618 41736 768674
rect 42706 768632 42762 768641
rect 41708 768590 42012 768618
rect 41696 767304 41748 767310
rect 41696 767246 41748 767252
rect 41708 765914 41736 767246
rect 41708 765886 41920 765914
rect 41696 764584 41748 764590
rect 41696 764526 41748 764532
rect 41708 763745 41736 764526
rect 41694 763736 41750 763745
rect 41694 763671 41750 763680
rect 41694 763328 41750 763337
rect 41694 763263 41696 763272
rect 41748 763263 41750 763272
rect 41696 763234 41748 763240
rect 41512 761048 41564 761054
rect 41512 760990 41564 760996
rect 41524 758690 41552 760990
rect 41892 758826 41920 765886
rect 41984 763154 42012 768590
rect 42706 768567 42762 768576
rect 41984 763126 42196 763154
rect 42168 758985 42196 763126
rect 42430 759520 42486 759529
rect 42486 759478 42656 759506
rect 42430 759455 42486 759464
rect 42154 758976 42210 758985
rect 42154 758911 42210 758920
rect 41892 758798 42564 758826
rect 41524 758662 42380 758690
rect 41604 757784 41656 757790
rect 40682 757752 40738 757761
rect 41656 757732 41828 757738
rect 41604 757726 41828 757732
rect 41616 757710 41828 757726
rect 40682 757687 40738 757696
rect 39946 757480 40002 757489
rect 39946 757415 40002 757424
rect 41800 757081 41828 757710
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 42352 756254 42380 758662
rect 42168 756226 42380 756254
rect 41878 755440 41934 755449
rect 41878 755375 41934 755384
rect 41892 755072 41920 755375
rect 42154 754896 42210 754905
rect 42154 754831 42210 754840
rect 42168 754392 42196 754831
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42340 753976 42392 753982
rect 42392 753924 42472 753930
rect 42340 753918 42472 753924
rect 42352 753902 42472 753918
rect 42248 753568 42300 753574
rect 42248 753510 42300 753516
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42076 751777 42104 751944
rect 42062 751768 42118 751777
rect 42062 751703 42118 751712
rect 42260 751383 42288 753510
rect 42182 751355 42288 751383
rect 42444 750938 42472 753902
rect 42168 750910 42472 750938
rect 42168 750720 42196 750910
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42536 749714 42564 758798
rect 42168 749686 42564 749714
rect 42168 749529 42196 749686
rect 42338 749592 42394 749601
rect 42338 749527 42394 749536
rect 42352 747062 42380 749527
rect 42182 747034 42380 747062
rect 41786 746736 41842 746745
rect 41786 746671 41842 746680
rect 41800 746401 41828 746671
rect 42628 746594 42656 759478
rect 42352 746566 42656 746594
rect 42352 746042 42380 746566
rect 42168 746014 42380 746042
rect 42168 745756 42196 746014
rect 42720 745498 42748 768567
rect 42168 745470 42748 745498
rect 42168 745212 42196 745470
rect 42522 745104 42578 745113
rect 42352 745062 42522 745090
rect 42062 744832 42118 744841
rect 42118 744790 42288 744818
rect 42062 744767 42118 744776
rect 41786 743744 41842 743753
rect 41786 743679 41842 743688
rect 41800 743376 41828 743679
rect 42260 743050 42288 744790
rect 42168 743022 42288 743050
rect 42168 742696 42196 743022
rect 42352 742098 42380 745062
rect 42522 745039 42578 745048
rect 42524 744048 42576 744054
rect 42524 743990 42576 743996
rect 42182 742070 42380 742098
rect 42536 741554 42564 743990
rect 42182 741526 42564 741554
rect 39578 732320 39634 732329
rect 39578 732255 39634 732264
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 35806 731368 35862 731377
rect 35806 731303 35862 731312
rect 35820 731134 35848 731303
rect 35808 731128 35860 731134
rect 35808 731070 35860 731076
rect 35622 730960 35678 730969
rect 35622 730895 35678 730904
rect 35438 730552 35494 730561
rect 35438 730487 35494 730496
rect 35254 729736 35310 729745
rect 35254 729671 35310 729680
rect 35268 728686 35296 729671
rect 35452 729434 35480 730487
rect 35636 730318 35664 730895
rect 35808 730584 35860 730590
rect 35808 730526 35860 730532
rect 35624 730312 35676 730318
rect 35624 730254 35676 730260
rect 35820 730153 35848 730526
rect 35806 730144 35862 730153
rect 35806 730079 35862 730088
rect 35440 729428 35492 729434
rect 35440 729370 35492 729376
rect 35622 729328 35678 729337
rect 35622 729263 35678 729272
rect 35636 728822 35664 729263
rect 35808 729088 35860 729094
rect 35808 729030 35860 729036
rect 35820 728929 35848 729030
rect 35806 728920 35862 728929
rect 35806 728855 35862 728864
rect 39592 728822 39620 732255
rect 39946 732048 40002 732057
rect 39946 731983 40002 731992
rect 39960 730590 39988 731983
rect 40406 731640 40462 731649
rect 40406 731575 40462 731584
rect 39948 730584 40000 730590
rect 39948 730526 40000 730532
rect 35624 728816 35676 728822
rect 35624 728758 35676 728764
rect 39580 728816 39632 728822
rect 39580 728758 39632 728764
rect 35256 728680 35308 728686
rect 35256 728622 35308 728628
rect 35622 728512 35678 728521
rect 35622 728447 35678 728456
rect 35636 727598 35664 728447
rect 35806 728104 35862 728113
rect 35806 728039 35862 728048
rect 35820 727870 35848 728039
rect 35808 727864 35860 727870
rect 35808 727806 35860 727812
rect 35806 727696 35862 727705
rect 35806 727631 35862 727640
rect 35624 727592 35676 727598
rect 35624 727534 35676 727540
rect 35820 727462 35848 727631
rect 40420 727598 40448 731575
rect 42064 731196 42116 731202
rect 42064 731138 42116 731144
rect 41696 731128 41748 731134
rect 42076 731082 42104 731138
rect 41748 731076 42104 731082
rect 41696 731070 42104 731076
rect 41708 731054 42104 731070
rect 41696 730312 41748 730318
rect 41694 730280 41696 730289
rect 41748 730280 41750 730289
rect 41694 730215 41750 730224
rect 41708 729434 42104 729450
rect 41696 729428 42104 729434
rect 41748 729422 42104 729428
rect 41696 729370 41748 729376
rect 42076 729366 42104 729422
rect 42064 729360 42116 729366
rect 42064 729302 42116 729308
rect 41696 729088 41748 729094
rect 41696 729030 41748 729036
rect 41708 728770 41736 729030
rect 41708 728742 42104 728770
rect 42076 728686 42104 728742
rect 41696 728680 41748 728686
rect 41694 728648 41696 728657
rect 42064 728680 42116 728686
rect 41748 728648 41750 728657
rect 42064 728622 42116 728628
rect 41694 728583 41750 728592
rect 42064 727932 42116 727938
rect 42064 727874 42116 727880
rect 41512 727864 41564 727870
rect 42076 727818 42104 727874
rect 41512 727806 41564 727812
rect 40408 727592 40460 727598
rect 40408 727534 40460 727540
rect 35808 727456 35860 727462
rect 35808 727398 35860 727404
rect 35808 727320 35860 727326
rect 35806 727288 35808 727297
rect 35860 727288 35862 727297
rect 35806 727223 35862 727232
rect 41524 727002 41552 727806
rect 41708 727790 42104 727818
rect 41708 727462 41736 727790
rect 41696 727456 41748 727462
rect 41696 727398 41748 727404
rect 41696 727320 41748 727326
rect 42064 727320 42116 727326
rect 41748 727268 42064 727274
rect 41696 727262 42116 727268
rect 41708 727246 42104 727262
rect 41694 727016 41750 727025
rect 41524 726974 41694 727002
rect 41694 726951 41750 726960
rect 41142 726880 41198 726889
rect 41142 726815 41198 726824
rect 39302 726234 39358 726243
rect 39302 726169 39358 726178
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 31666 724432 31722 724441
rect 31666 724367 31722 724376
rect 31680 718321 31708 724367
rect 33046 724024 33102 724033
rect 33046 723959 33102 723968
rect 31666 718312 31722 718321
rect 31666 718247 31722 718256
rect 33060 715562 33088 723959
rect 33782 723208 33838 723217
rect 33782 723143 33838 723152
rect 33796 715698 33824 723143
rect 35176 715834 35204 724775
rect 39316 716145 39344 726169
rect 41156 725966 41184 726815
rect 41326 726234 41382 726243
rect 41326 726169 41382 726178
rect 41696 726232 41748 726238
rect 41748 726180 42196 726186
rect 41696 726174 42196 726180
rect 41708 726158 42196 726174
rect 41144 725960 41196 725966
rect 41144 725902 41196 725908
rect 41604 725960 41656 725966
rect 41604 725902 41656 725908
rect 41616 725778 41644 725902
rect 41786 725792 41842 725801
rect 41616 725750 41786 725778
rect 41786 725727 41842 725736
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41142 725248 41198 725257
rect 41142 725183 41198 725192
rect 41156 719273 41184 725183
rect 41340 724514 41368 725591
rect 42168 724514 42196 726158
rect 41340 724486 41552 724514
rect 42168 724486 42288 724514
rect 41326 720352 41382 720361
rect 41326 720287 41382 720296
rect 41142 719264 41198 719273
rect 41142 719199 41198 719208
rect 41340 717614 41368 720287
rect 41524 719001 41552 724486
rect 41970 722392 42026 722401
rect 41970 722327 42026 722336
rect 41786 721984 41842 721993
rect 41786 721919 41842 721928
rect 41510 718992 41566 719001
rect 41510 718927 41566 718936
rect 41800 718593 41828 721919
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 41984 718049 42012 722327
rect 41970 718040 42026 718049
rect 41970 717975 42026 717984
rect 41248 717586 41368 717614
rect 39302 716136 39358 716145
rect 39302 716071 39358 716080
rect 35164 715828 35216 715834
rect 35164 715770 35216 715776
rect 33784 715692 33836 715698
rect 33784 715634 33836 715640
rect 37740 715692 37792 715698
rect 37740 715634 37792 715640
rect 33048 715556 33100 715562
rect 33048 715498 33100 715504
rect 37752 714513 37780 715634
rect 39854 715592 39910 715601
rect 39854 715527 39856 715536
rect 39908 715527 39910 715536
rect 39856 715498 39908 715504
rect 37738 714504 37794 714513
rect 37738 714439 37794 714448
rect 41248 714241 41276 717586
rect 41696 715828 41748 715834
rect 41696 715770 41748 715776
rect 41708 714354 41736 715770
rect 42260 715442 42288 724486
rect 42614 719264 42670 719273
rect 42670 719222 42840 719250
rect 42614 719199 42670 719208
rect 42614 718992 42670 719001
rect 42614 718927 42670 718936
rect 42430 715592 42486 715601
rect 42430 715527 42486 715536
rect 42444 715442 42472 715527
rect 42260 715414 42380 715442
rect 42444 715414 42564 715442
rect 42352 714898 42380 715414
rect 42536 715034 42564 715414
rect 42628 715170 42656 718927
rect 42628 715142 42748 715170
rect 42536 715006 42656 715034
rect 42352 714870 42472 714898
rect 42062 714504 42118 714513
rect 42118 714462 42380 714490
rect 42062 714439 42118 714448
rect 41708 714326 42288 714354
rect 41234 714232 41290 714241
rect 41234 714167 41290 714176
rect 42260 713062 42288 714326
rect 42182 713034 42288 713062
rect 42352 712858 42380 714462
rect 42260 712830 42380 712858
rect 41786 712192 41842 712201
rect 41786 712127 41842 712136
rect 41800 711824 41828 712127
rect 42260 711754 42288 712830
rect 42248 711748 42300 711754
rect 42248 711690 42300 711696
rect 42444 711634 42472 714870
rect 42628 713474 42656 715006
rect 42352 711606 42472 711634
rect 42536 713446 42656 713474
rect 42352 711498 42380 711606
rect 42168 711470 42380 711498
rect 42168 711212 42196 711470
rect 42248 711136 42300 711142
rect 42300 711084 42380 711090
rect 42248 711078 42380 711084
rect 42260 711062 42380 711078
rect 42154 710832 42210 710841
rect 42154 710767 42210 710776
rect 42168 710561 42196 710767
rect 42352 709390 42380 711062
rect 42182 709362 42380 709390
rect 42248 709232 42300 709238
rect 42248 709174 42300 709180
rect 42076 708529 42104 708696
rect 42062 708520 42118 708529
rect 42062 708455 42118 708464
rect 42260 708234 42288 709174
rect 42168 708206 42288 708234
rect 42168 708152 42196 708206
rect 42062 707704 42118 707713
rect 42536 707690 42564 713446
rect 42720 710002 42748 715142
rect 42062 707639 42118 707648
rect 42444 707662 42564 707690
rect 42628 709974 42748 710002
rect 42076 707540 42104 707639
rect 41786 707432 41842 707441
rect 41786 707367 41842 707376
rect 41800 706860 41828 707367
rect 42444 707130 42472 707662
rect 42628 707470 42656 709974
rect 42616 707464 42668 707470
rect 42616 707406 42668 707412
rect 42432 707124 42484 707130
rect 42432 707066 42484 707072
rect 42812 707010 42840 719222
rect 42536 706982 42840 707010
rect 42536 706874 42564 706982
rect 42260 706846 42564 706874
rect 42260 706738 42288 706846
rect 42168 706710 42288 706738
rect 42616 706716 42668 706722
rect 42168 706602 42196 706710
rect 42616 706658 42668 706664
rect 42076 706574 42196 706602
rect 42432 706648 42484 706654
rect 42432 706590 42484 706596
rect 42076 706316 42104 706574
rect 42246 706208 42302 706217
rect 42246 706143 42302 706152
rect 42260 704290 42288 706143
rect 42444 705194 42472 706590
rect 42628 706330 42656 706658
rect 42536 706302 42656 706330
rect 42536 706058 42564 706302
rect 42536 706030 42656 706058
rect 42444 705166 42564 705194
rect 42076 704262 42288 704290
rect 42076 703868 42104 704262
rect 42062 703488 42118 703497
rect 42062 703423 42118 703432
rect 42076 703188 42104 703423
rect 42536 702658 42564 705166
rect 42352 702630 42564 702658
rect 42352 702590 42380 702630
rect 42168 702522 42196 702576
rect 42260 702562 42380 702590
rect 42260 702522 42288 702562
rect 42168 702494 42288 702522
rect 42628 702250 42656 706030
rect 42444 702222 42656 702250
rect 42444 702046 42472 702222
rect 42706 702128 42762 702137
rect 42168 701978 42196 702032
rect 42260 702018 42472 702046
rect 42536 702086 42706 702114
rect 42260 701978 42288 702018
rect 42168 701950 42288 701978
rect 42338 701856 42394 701865
rect 42338 701791 42394 701800
rect 41786 700496 41842 700505
rect 41786 700431 41842 700440
rect 41800 700165 41828 700431
rect 42352 699530 42380 701791
rect 42182 699502 42380 699530
rect 42536 698918 42564 702086
rect 42706 702063 42762 702072
rect 42708 701072 42760 701078
rect 42708 701014 42760 701020
rect 42168 698850 42196 698904
rect 42260 698890 42564 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 42720 698339 42748 701014
rect 42182 698311 42748 698339
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 42706 688120 42762 688129
rect 42706 688055 42762 688064
rect 42720 687342 42748 688055
rect 42708 687336 42760 687342
rect 42708 687278 42760 687284
rect 40866 686896 40922 686905
rect 40866 686831 40922 686840
rect 40880 685914 40908 686831
rect 41142 686488 41198 686497
rect 41142 686423 41198 686432
rect 41156 686050 41184 686423
rect 41144 686044 41196 686050
rect 41144 685986 41196 685992
rect 41696 686044 41748 686050
rect 42064 686044 42116 686050
rect 41748 686004 42064 686032
rect 41696 685986 41748 685992
rect 42064 685986 42116 685992
rect 40868 685908 40920 685914
rect 40868 685850 40920 685856
rect 41050 685910 41106 685919
rect 41050 685845 41106 685854
rect 41696 685908 41748 685914
rect 42064 685908 42116 685914
rect 41748 685868 42064 685896
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 40866 684856 40922 684865
rect 40866 684791 40922 684800
rect 40880 684622 40908 684791
rect 41064 684758 41092 685845
rect 41052 684752 41104 684758
rect 41696 684752 41748 684758
rect 41052 684694 41104 684700
rect 41694 684720 41696 684729
rect 41748 684720 41750 684729
rect 41694 684655 41750 684664
rect 40868 684616 40920 684622
rect 40868 684558 40920 684564
rect 41708 684554 42104 684570
rect 41696 684548 42116 684554
rect 41748 684542 42064 684548
rect 41696 684490 41748 684496
rect 42064 684490 42116 684496
rect 41326 683462 41382 683471
rect 41326 683397 41382 683406
rect 41696 683460 41748 683466
rect 41696 683402 41748 683408
rect 40958 682816 41014 682825
rect 40958 682751 41014 682760
rect 35162 682000 35218 682009
rect 35162 681935 35218 681944
rect 32402 681184 32458 681193
rect 32402 681119 32458 681128
rect 32416 672761 32444 681119
rect 33782 680776 33838 680785
rect 33782 680711 33838 680720
rect 33796 672790 33824 680711
rect 35176 672926 35204 681935
rect 40972 679182 41000 682751
rect 41708 681850 41736 683402
rect 42522 682408 42578 682417
rect 42522 682343 42578 682352
rect 41708 681822 42472 681850
rect 42246 681592 42302 681601
rect 42246 681527 42302 681536
rect 41142 679960 41198 679969
rect 41142 679895 41198 679904
rect 40960 679176 41012 679182
rect 40960 679118 41012 679124
rect 41156 679046 41184 679895
rect 41328 679176 41380 679182
rect 41328 679118 41380 679124
rect 41144 679040 41196 679046
rect 41144 678982 41196 678988
rect 41340 678858 41368 679118
rect 41696 679040 41748 679046
rect 42064 679040 42116 679046
rect 41748 679000 42064 679028
rect 41696 678982 41748 678988
rect 42064 678982 42116 678988
rect 41786 678872 41842 678881
rect 41340 678830 41786 678858
rect 41786 678807 41842 678816
rect 41786 678328 41842 678337
rect 41616 678286 41786 678314
rect 40958 677750 41014 677759
rect 41616 677754 41644 678286
rect 41786 678263 41842 678272
rect 40958 677685 41014 677694
rect 41604 677748 41656 677754
rect 41604 677690 41656 677696
rect 39946 677104 40002 677113
rect 39946 677039 40002 677048
rect 39960 673033 39988 677039
rect 42260 674370 42288 681527
rect 42444 676214 42472 681822
rect 42076 674342 42288 674370
rect 42352 676186 42472 676214
rect 42536 676214 42564 682343
rect 42904 676214 42932 796198
rect 43180 795138 43208 804526
rect 43088 795110 43208 795138
rect 43088 795054 43116 795110
rect 43076 795048 43128 795054
rect 43076 794990 43128 794996
rect 43076 794912 43128 794918
rect 43076 794854 43128 794860
rect 43088 794102 43116 794854
rect 43076 794096 43128 794102
rect 43076 794038 43128 794044
rect 43074 771488 43130 771497
rect 43074 771423 43130 771432
rect 43088 732329 43116 771423
rect 43272 770681 43300 812806
rect 43812 805996 43864 806002
rect 43812 805938 43864 805944
rect 43628 801100 43680 801106
rect 43628 801042 43680 801048
rect 43444 799060 43496 799066
rect 43444 799002 43496 799008
rect 43456 797337 43484 799002
rect 43442 797328 43498 797337
rect 43442 797263 43498 797272
rect 43640 796550 43668 801042
rect 43628 796544 43680 796550
rect 43628 796486 43680 796492
rect 43258 770672 43314 770681
rect 43258 770607 43314 770616
rect 43626 764144 43682 764153
rect 43626 764079 43682 764088
rect 43258 757480 43314 757489
rect 43258 757415 43314 757424
rect 43074 732320 43130 732329
rect 43074 732255 43130 732264
rect 43076 728680 43128 728686
rect 43076 728622 43128 728628
rect 43088 686089 43116 728622
rect 43074 686080 43130 686089
rect 43074 686015 43130 686024
rect 43074 677920 43130 677929
rect 43074 677855 43130 677864
rect 42536 676186 42656 676214
rect 39946 673024 40002 673033
rect 39946 672959 40002 672968
rect 35164 672920 35216 672926
rect 35164 672862 35216 672868
rect 38936 672920 38988 672926
rect 38936 672862 38988 672868
rect 33784 672784 33836 672790
rect 32402 672752 32458 672761
rect 33784 672726 33836 672732
rect 38200 672784 38252 672790
rect 38200 672726 38252 672732
rect 32402 672687 32458 672696
rect 38212 670993 38240 672726
rect 38948 671265 38976 672862
rect 38934 671256 38990 671265
rect 38934 671191 38990 671200
rect 38198 670984 38254 670993
rect 38198 670919 38254 670928
rect 42076 670834 42104 674342
rect 42076 670806 42288 670834
rect 42168 669746 42196 669868
rect 42260 669746 42288 670806
rect 42168 669718 42288 669746
rect 41786 669080 41842 669089
rect 41786 669015 41842 669024
rect 41800 668644 41828 669015
rect 42352 668522 42380 676186
rect 42260 668494 42380 668522
rect 42260 668386 42288 668494
rect 41984 668358 42288 668386
rect 41984 668032 42012 668358
rect 42248 667480 42300 667486
rect 42248 667422 42300 667428
rect 42260 667366 42288 667422
rect 42182 667338 42288 667366
rect 42628 666652 42656 676186
rect 42812 676186 42932 676214
rect 42812 671514 42840 676186
rect 43088 671650 43116 677855
rect 43272 671945 43300 757415
rect 43444 754928 43496 754934
rect 43444 754870 43496 754876
rect 43456 753001 43484 754870
rect 43640 753982 43668 764079
rect 43628 753976 43680 753982
rect 43628 753918 43680 753924
rect 43442 752992 43498 753001
rect 43442 752927 43498 752936
rect 43442 723616 43498 723625
rect 43442 723551 43498 723560
rect 43456 703497 43484 723551
rect 43628 712156 43680 712162
rect 43628 712098 43680 712104
rect 43640 710841 43668 712098
rect 43626 710832 43682 710841
rect 43626 710767 43682 710776
rect 43628 709368 43680 709374
rect 43628 709310 43680 709316
rect 43640 707713 43668 709310
rect 43626 707704 43682 707713
rect 43626 707639 43682 707648
rect 43442 703488 43498 703497
rect 43442 703423 43498 703432
rect 43442 687304 43498 687313
rect 43442 687239 43498 687248
rect 43456 686526 43484 687239
rect 43444 686520 43496 686526
rect 43444 686462 43496 686468
rect 43626 680368 43682 680377
rect 43626 680303 43682 680312
rect 43442 676696 43498 676705
rect 43442 676631 43498 676640
rect 43456 676214 43484 676631
rect 43456 676186 43576 676214
rect 43258 671936 43314 671945
rect 43258 671871 43314 671880
rect 43088 671622 43300 671650
rect 42812 671486 43208 671514
rect 42798 671256 42854 671265
rect 42798 671191 42854 671200
rect 42154 666632 42210 666641
rect 42154 666567 42210 666576
rect 42536 666624 42656 666652
rect 42168 666165 42196 666567
rect 42536 666482 42564 666624
rect 42536 666454 42656 666482
rect 42062 665952 42118 665961
rect 42062 665887 42118 665896
rect 42076 665516 42104 665887
rect 42430 665544 42486 665553
rect 42430 665479 42486 665488
rect 42246 665272 42302 665281
rect 42246 665207 42302 665216
rect 42260 664986 42288 665207
rect 42444 665174 42472 665479
rect 42444 665146 42564 665174
rect 42182 664958 42288 664986
rect 42248 664896 42300 664902
rect 42248 664838 42300 664844
rect 42260 664339 42288 664838
rect 42536 664714 42564 665146
rect 42352 664686 42564 664714
rect 42352 664442 42380 664686
rect 42628 664442 42656 666454
rect 42812 665174 42840 671191
rect 43180 666924 43208 671486
rect 42352 664414 42472 664442
rect 42182 664311 42288 664339
rect 42248 664216 42300 664222
rect 42248 664158 42300 664164
rect 41786 664048 41842 664057
rect 41786 663983 41842 663992
rect 41800 663680 41828 663983
rect 42260 663150 42288 664158
rect 42182 663122 42288 663150
rect 42248 663060 42300 663066
rect 42248 663002 42300 663008
rect 42062 662824 42118 662833
rect 42260 662810 42288 663002
rect 42260 662782 42380 662810
rect 42062 662759 42118 662768
rect 42076 662674 42104 662759
rect 42076 662646 42288 662674
rect 42260 661042 42288 662646
rect 42168 661014 42288 661042
rect 42168 660620 42196 661014
rect 42352 660022 42380 662782
rect 42182 659994 42380 660022
rect 42444 659371 42472 664414
rect 42536 664414 42656 664442
rect 42720 665146 42840 665174
rect 42904 666896 43208 666924
rect 42536 659954 42564 664414
rect 42720 664222 42748 665146
rect 42708 664216 42760 664222
rect 42708 664158 42760 664164
rect 42706 660920 42762 660929
rect 42706 660855 42762 660864
rect 42536 659926 42656 659954
rect 42628 659654 42656 659926
rect 42182 659343 42472 659371
rect 42536 659626 42656 659654
rect 42536 659002 42564 659626
rect 42168 658974 42564 659002
rect 42168 658784 42196 658974
rect 42522 658608 42578 658617
rect 42352 658566 42522 658594
rect 41800 658430 42288 658458
rect 41800 658345 41828 658430
rect 41786 658336 41842 658345
rect 41786 658271 41842 658280
rect 42064 657416 42116 657422
rect 42064 657358 42116 657364
rect 42076 656948 42104 657358
rect 42260 656350 42288 658430
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42352 655670 42380 658566
rect 42522 658543 42578 658552
rect 42524 657552 42576 657558
rect 42524 657494 42576 657500
rect 42260 655642 42380 655670
rect 42536 655126 42564 657494
rect 42720 657422 42748 660855
rect 42708 657416 42760 657422
rect 42708 657358 42760 657364
rect 42182 655098 42564 655126
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 40130 644736 40186 644745
rect 40130 644671 40186 644680
rect 35820 644502 35848 644671
rect 35808 644496 35860 644502
rect 35808 644438 35860 644444
rect 38566 644328 38622 644337
rect 38566 644263 38622 644272
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 35622 642696 35678 642705
rect 35622 642631 35678 642640
rect 35636 642054 35664 642631
rect 38580 642530 38608 644263
rect 39948 643544 40000 643550
rect 39948 643486 40000 643492
rect 39960 643113 39988 643486
rect 39946 643104 40002 643113
rect 39946 643039 40002 643048
rect 38568 642524 38620 642530
rect 38568 642466 38620 642472
rect 35806 642288 35862 642297
rect 35806 642223 35862 642232
rect 35624 642048 35676 642054
rect 35624 641990 35676 641996
rect 35820 641782 35848 642223
rect 40144 642054 40172 644671
rect 41696 644496 41748 644502
rect 42064 644496 42116 644502
rect 41748 644446 42064 644474
rect 41696 644438 41748 644444
rect 42064 644438 42116 644444
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 41696 642524 41748 642530
rect 41748 642484 42104 642512
rect 41696 642466 41748 642472
rect 42076 642394 42104 642484
rect 42064 642388 42116 642394
rect 42064 642330 42116 642336
rect 40132 642048 40184 642054
rect 40132 641990 40184 641996
rect 35808 641776 35860 641782
rect 35808 641718 35860 641724
rect 41696 641776 41748 641782
rect 42064 641776 42116 641782
rect 41748 641724 42064 641730
rect 41696 641718 42116 641724
rect 41708 641702 42104 641718
rect 35438 641472 35494 641481
rect 35438 641407 35494 641416
rect 35452 640490 35480 641407
rect 35806 641064 35862 641073
rect 35806 640999 35862 641008
rect 39762 641064 39818 641073
rect 39762 640999 39818 641008
rect 35820 640762 35848 640999
rect 39776 640762 39804 640999
rect 35808 640756 35860 640762
rect 35808 640698 35860 640704
rect 39764 640756 39816 640762
rect 39764 640698 39816 640704
rect 35622 640656 35678 640665
rect 35622 640591 35678 640600
rect 35440 640484 35492 640490
rect 35440 640426 35492 640432
rect 35636 640354 35664 640591
rect 40040 640484 40092 640490
rect 40040 640426 40092 640432
rect 35624 640348 35676 640354
rect 35624 640290 35676 640296
rect 40052 640257 40080 640426
rect 41696 640348 41748 640354
rect 42064 640348 42116 640354
rect 41748 640306 42064 640334
rect 41696 640290 41748 640296
rect 42064 640290 42116 640296
rect 40038 640248 40094 640257
rect 40038 640183 40094 640192
rect 35806 639840 35862 639849
rect 35806 639775 35862 639784
rect 35820 639198 35848 639775
rect 35808 639192 35860 639198
rect 35808 639134 35860 639140
rect 37924 639124 37976 639130
rect 37924 639066 37976 639072
rect 35806 639024 35862 639033
rect 35806 638959 35808 638968
rect 35860 638959 35862 638968
rect 35808 638930 35860 638936
rect 35622 638616 35678 638625
rect 35622 638551 35678 638560
rect 35162 637800 35218 637809
rect 35162 637735 35218 637744
rect 31942 636984 31998 636993
rect 31942 636919 31998 636928
rect 31956 629950 31984 636919
rect 31944 629944 31996 629950
rect 35176 629921 35204 637735
rect 35636 636954 35664 638551
rect 35806 638208 35862 638217
rect 35806 638143 35862 638152
rect 35820 637770 35848 638143
rect 35808 637764 35860 637770
rect 35808 637706 35860 637712
rect 36544 637764 36596 637770
rect 36544 637706 36596 637712
rect 35624 636948 35676 636954
rect 35624 636890 35676 636896
rect 35530 636576 35586 636585
rect 35530 636511 35532 636520
rect 35584 636511 35586 636520
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35532 636482 35584 636488
rect 35820 636274 35848 636511
rect 35808 636268 35860 636274
rect 35808 636210 35860 636216
rect 35806 635760 35862 635769
rect 35806 635695 35862 635704
rect 35820 634982 35848 635695
rect 35808 634976 35860 634982
rect 35808 634918 35860 634924
rect 35622 634536 35678 634545
rect 35622 634471 35678 634480
rect 35636 633486 35664 634471
rect 35808 633752 35860 633758
rect 35806 633720 35808 633729
rect 35860 633720 35862 633729
rect 35806 633655 35862 633664
rect 35624 633480 35676 633486
rect 35624 633422 35676 633428
rect 36556 630766 36584 637706
rect 37936 631417 37964 639066
rect 41420 638920 41472 638926
rect 41420 638862 41472 638868
rect 40684 636948 40736 636954
rect 40684 636890 40736 636896
rect 40696 636585 40724 636890
rect 40682 636576 40738 636585
rect 40682 636511 40738 636520
rect 39856 636472 39908 636478
rect 39856 636414 39908 636420
rect 39868 636177 39896 636414
rect 39854 636168 39910 636177
rect 39854 636103 39910 636112
rect 38566 633720 38622 633729
rect 38566 633655 38622 633664
rect 39580 633684 39632 633690
rect 37922 631408 37978 631417
rect 37922 631343 37978 631352
rect 36544 630760 36596 630766
rect 36544 630702 36596 630708
rect 31944 629886 31996 629892
rect 35162 629912 35218 629921
rect 35162 629847 35218 629856
rect 38580 628318 38608 633655
rect 39580 633626 39632 633632
rect 39592 630737 39620 633626
rect 40132 633480 40184 633486
rect 40132 633422 40184 633428
rect 40144 631961 40172 633422
rect 41432 632913 41460 638862
rect 42706 636576 42762 636585
rect 42706 636511 42762 636520
rect 42720 636426 42748 636511
rect 42720 636398 42840 636426
rect 41708 636274 42104 636290
rect 41696 636268 42116 636274
rect 41748 636262 42064 636268
rect 41696 636210 41748 636216
rect 42064 636210 42116 636216
rect 41604 634976 41656 634982
rect 41602 634944 41604 634953
rect 41656 634944 41658 634953
rect 41602 634879 41658 634888
rect 41418 632904 41474 632913
rect 41418 632839 41474 632848
rect 40130 631952 40186 631961
rect 40130 631887 40186 631896
rect 42614 631408 42670 631417
rect 42614 631343 42670 631352
rect 41604 630760 41656 630766
rect 39578 630728 39634 630737
rect 41604 630702 41656 630708
rect 39578 630663 39634 630672
rect 40224 629944 40276 629950
rect 40224 629886 40276 629892
rect 40236 629241 40264 629886
rect 40222 629232 40278 629241
rect 40222 629167 40278 629176
rect 38568 628312 38620 628318
rect 40500 628312 40552 628318
rect 38568 628254 38620 628260
rect 40498 628280 40500 628289
rect 40552 628280 40554 628289
rect 40498 628215 40554 628224
rect 41616 627722 41644 630702
rect 42154 629232 42210 629241
rect 42154 629167 42210 629176
rect 42168 628130 42196 629167
rect 42338 628314 42394 628323
rect 42394 628258 42472 628266
rect 42338 628249 42472 628258
rect 42352 628238 42472 628249
rect 42168 628102 42380 628130
rect 41616 627694 42288 627722
rect 42260 627178 42288 627694
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 627042 42380 628102
rect 42260 627014 42380 627042
rect 42260 625705 42288 627014
rect 42246 625696 42302 625705
rect 42246 625631 42302 625640
rect 42444 625478 42472 628238
rect 42628 626534 42656 631343
rect 42182 625450 42472 625478
rect 42536 626506 42656 626534
rect 42536 625394 42564 626506
rect 42248 625388 42300 625394
rect 42248 625330 42300 625336
rect 42524 625388 42576 625394
rect 42524 625330 42576 625336
rect 42260 624866 42288 625330
rect 42812 625138 42840 636398
rect 42720 625122 42840 625138
rect 42524 625116 42576 625122
rect 42524 625058 42576 625064
rect 42708 625116 42840 625122
rect 42760 625110 42840 625116
rect 42708 625058 42760 625064
rect 42168 624838 42288 624866
rect 42168 624784 42196 624838
rect 42340 624436 42392 624442
rect 42340 624378 42392 624384
rect 42352 624186 42380 624378
rect 42182 624158 42380 624186
rect 42248 624096 42300 624102
rect 42248 624038 42300 624044
rect 42260 623914 42288 624038
rect 42260 623886 42380 623914
rect 42062 623792 42118 623801
rect 42118 623750 42288 623778
rect 42062 623727 42118 623736
rect 42062 623384 42118 623393
rect 42062 623319 42118 623328
rect 42076 622948 42104 623319
rect 42076 622169 42104 622336
rect 42062 622160 42118 622169
rect 42062 622095 42118 622104
rect 42168 621738 42196 621792
rect 42260 621738 42288 623750
rect 42168 621710 42288 621738
rect 42352 621126 42380 623886
rect 42182 621098 42380 621126
rect 41786 620936 41842 620945
rect 41786 620871 41842 620880
rect 41800 620500 41828 620871
rect 42536 619970 42564 625058
rect 42706 624608 42762 624617
rect 42706 624543 42762 624552
rect 42168 619834 42196 619956
rect 42260 619942 42564 619970
rect 42260 619834 42288 619942
rect 42168 619806 42288 619834
rect 42522 619848 42578 619857
rect 42522 619783 42578 619792
rect 42248 619676 42300 619682
rect 42248 619618 42300 619624
rect 42260 617454 42288 619618
rect 42182 617426 42288 617454
rect 42536 617114 42564 619783
rect 42352 617086 42564 617114
rect 42352 616842 42380 617086
rect 42168 616706 42196 616828
rect 42260 616814 42380 616842
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 41786 616448 41842 616457
rect 41786 616383 41842 616392
rect 41800 616148 41828 616383
rect 42720 616298 42748 624543
rect 42260 616270 42748 616298
rect 42260 616026 42288 616270
rect 42614 616176 42670 616185
rect 42614 616111 42670 616120
rect 42168 615998 42288 616026
rect 42168 615604 42196 615998
rect 42338 615768 42394 615777
rect 42338 615703 42394 615712
rect 42352 615482 42380 615703
rect 42260 615454 42380 615482
rect 42260 613782 42288 615454
rect 42628 615346 42656 616111
rect 42182 613754 42288 613782
rect 42352 615318 42656 615346
rect 42352 613135 42380 615318
rect 42614 615224 42670 615233
rect 42182 613107 42380 613135
rect 42444 615182 42614 615210
rect 42444 612490 42472 615182
rect 42614 615159 42670 615168
rect 42616 614168 42668 614174
rect 42616 614110 42668 614116
rect 42182 612462 42472 612490
rect 42628 611946 42656 614110
rect 42904 613873 42932 666896
rect 43272 666754 43300 671622
rect 43088 666726 43300 666754
rect 43548 666754 43576 676186
rect 43640 669314 43668 680303
rect 43640 669286 43760 669314
rect 43548 666726 43668 666754
rect 43088 615466 43116 666726
rect 43258 666568 43314 666577
rect 43640 666554 43668 666726
rect 43258 666503 43314 666512
rect 43456 666526 43668 666554
rect 43076 615460 43128 615466
rect 43076 615402 43128 615408
rect 42890 613864 42946 613873
rect 42890 613799 42946 613808
rect 43272 612241 43300 666503
rect 43258 612232 43314 612241
rect 43258 612167 43314 612176
rect 42182 611918 42656 611946
rect 43456 611402 43484 666526
rect 43732 663082 43760 669286
rect 43640 663066 43760 663082
rect 43628 663060 43760 663066
rect 43680 663054 43760 663060
rect 43628 663002 43680 663008
rect 43626 631952 43682 631961
rect 43626 631887 43682 631896
rect 43640 612354 43668 631887
rect 43824 612610 43852 805938
rect 44284 772313 44312 814370
rect 44548 814292 44600 814298
rect 44548 814234 44600 814240
rect 44270 772304 44326 772313
rect 44270 772239 44326 772248
rect 44560 771526 44588 814234
rect 44836 806614 44864 815730
rect 45008 815652 45060 815658
rect 45008 815594 45060 815600
rect 44824 806608 44876 806614
rect 44824 806550 44876 806556
rect 45020 776665 45048 815594
rect 45192 807356 45244 807362
rect 45192 807298 45244 807304
rect 45204 794918 45232 807298
rect 45192 794912 45244 794918
rect 45192 794854 45244 794860
rect 46216 785194 46244 817090
rect 61384 817012 61436 817018
rect 61384 816954 61436 816960
rect 53104 799060 53156 799066
rect 53104 799002 53156 799008
rect 53116 790770 53144 799002
rect 57244 797700 57296 797706
rect 57244 797642 57296 797648
rect 53104 790764 53156 790770
rect 53104 790706 53156 790712
rect 57256 789206 57284 797642
rect 57244 789200 57296 789206
rect 57244 789142 57296 789148
rect 61396 786185 61424 816954
rect 62764 806608 62816 806614
rect 62764 806550 62816 806556
rect 62212 790764 62264 790770
rect 62212 790706 62264 790712
rect 62224 790537 62252 790706
rect 62210 790528 62266 790537
rect 62210 790463 62266 790472
rect 62120 789200 62172 789206
rect 62118 789168 62120 789177
rect 62172 789168 62174 789177
rect 62118 789103 62174 789112
rect 62118 787400 62174 787409
rect 62118 787335 62174 787344
rect 62132 786690 62160 787335
rect 62776 787137 62804 806550
rect 669228 790968 669280 790974
rect 669228 790910 669280 790916
rect 653404 790832 653456 790838
rect 653404 790774 653456 790780
rect 62762 787128 62818 787137
rect 62762 787063 62818 787072
rect 62120 786684 62172 786690
rect 62120 786626 62172 786632
rect 61382 786176 61438 786185
rect 61382 786111 61438 786120
rect 46204 785188 46256 785194
rect 46204 785130 46256 785136
rect 62120 785188 62172 785194
rect 62120 785130 62172 785136
rect 62132 784961 62160 785130
rect 62118 784952 62174 784961
rect 62118 784887 62174 784896
rect 651470 778424 651526 778433
rect 651470 778359 651526 778368
rect 651484 777646 651512 778359
rect 651472 777640 651524 777646
rect 651472 777582 651524 777588
rect 652022 777064 652078 777073
rect 652022 776999 652078 777008
rect 45006 776656 45062 776665
rect 45006 776591 45062 776600
rect 651470 776112 651526 776121
rect 651470 776047 651526 776056
rect 651484 775742 651512 776047
rect 651472 775736 651524 775742
rect 651472 775678 651524 775684
rect 651380 775328 651432 775334
rect 651378 775296 651380 775305
rect 651432 775296 651434 775305
rect 651378 775231 651434 775240
rect 60004 774240 60056 774246
rect 60004 774182 60056 774188
rect 651470 774208 651526 774217
rect 44914 773120 44970 773129
rect 44914 773055 44970 773064
rect 44548 771520 44600 771526
rect 44548 771462 44600 771468
rect 44272 770092 44324 770098
rect 44272 770034 44324 770040
rect 44284 727938 44312 770034
rect 44546 767000 44602 767009
rect 44546 766935 44602 766944
rect 44560 731649 44588 766935
rect 44732 755540 44784 755546
rect 44732 755482 44784 755488
rect 44744 754089 44772 755482
rect 44730 754080 44786 754089
rect 44730 754015 44786 754024
rect 44928 732057 44956 773055
rect 46204 773016 46256 773022
rect 46204 772958 46256 772964
rect 45098 764552 45154 764561
rect 45098 764487 45154 764496
rect 45112 754934 45140 764487
rect 45282 763736 45338 763745
rect 45282 763671 45338 763680
rect 45100 754928 45152 754934
rect 45100 754870 45152 754876
rect 45296 753574 45324 763671
rect 45558 763328 45614 763337
rect 45558 763263 45614 763272
rect 45284 753568 45336 753574
rect 45284 753510 45336 753516
rect 45098 751768 45154 751777
rect 45098 751703 45154 751712
rect 45112 746570 45140 751703
rect 45100 746564 45152 746570
rect 45100 746506 45152 746512
rect 44914 732048 44970 732057
rect 44914 731983 44970 731992
rect 44546 731640 44602 731649
rect 44546 731575 44602 731584
rect 45190 728648 45246 728657
rect 45190 728583 45246 728592
rect 44272 727932 44324 727938
rect 44272 727874 44324 727880
rect 45008 727320 45060 727326
rect 45008 727262 45060 727268
rect 44270 727016 44326 727025
rect 44270 726951 44326 726960
rect 44284 685273 44312 726951
rect 44454 722800 44510 722809
rect 44454 722735 44510 722744
rect 44468 709374 44496 722735
rect 44638 721576 44694 721585
rect 44638 721511 44694 721520
rect 44456 709368 44508 709374
rect 44456 709310 44508 709316
rect 44652 709238 44680 721511
rect 44640 709232 44692 709238
rect 44640 709174 44692 709180
rect 44454 708520 44510 708529
rect 44454 708455 44510 708464
rect 44468 703798 44496 708455
rect 44456 703792 44508 703798
rect 44456 703734 44508 703740
rect 44822 687712 44878 687721
rect 44822 687647 44878 687656
rect 44640 686044 44692 686050
rect 44640 685986 44692 685992
rect 44270 685264 44326 685273
rect 44270 685199 44326 685208
rect 44454 684720 44510 684729
rect 44454 684655 44510 684664
rect 44270 684040 44326 684049
rect 44270 683975 44326 683984
rect 43994 679552 44050 679561
rect 43994 679487 44050 679496
rect 44008 664902 44036 679487
rect 43996 664896 44048 664902
rect 43996 664838 44048 664844
rect 44284 641073 44312 683975
rect 44468 644745 44496 684655
rect 44454 644736 44510 644745
rect 44454 644671 44510 644680
rect 44652 643346 44680 685986
rect 44836 655518 44864 687647
rect 45020 684457 45048 727262
rect 45204 685914 45232 728583
rect 45192 685908 45244 685914
rect 45192 685850 45244 685856
rect 45192 684548 45244 684554
rect 45192 684490 45244 684496
rect 45006 684448 45062 684457
rect 45006 684383 45062 684392
rect 45008 679040 45060 679046
rect 45008 678982 45060 678988
rect 45020 667457 45048 678982
rect 45006 667448 45062 667457
rect 45006 667383 45062 667392
rect 44824 655512 44876 655518
rect 44824 655454 44876 655460
rect 44640 643340 44692 643346
rect 44640 643282 44692 643288
rect 44730 643104 44786 643113
rect 44730 643039 44786 643048
rect 44270 641064 44326 641073
rect 44270 640999 44326 641008
rect 44548 636268 44600 636274
rect 44548 636210 44600 636216
rect 43994 636168 44050 636177
rect 43994 636103 44050 636112
rect 44008 623393 44036 636103
rect 44362 634944 44418 634953
rect 44362 634879 44418 634888
rect 44180 625864 44232 625870
rect 44180 625806 44232 625812
rect 44192 624442 44220 625806
rect 44180 624436 44232 624442
rect 44180 624378 44232 624384
rect 44376 624322 44404 634879
rect 44560 634794 44588 636210
rect 44744 635474 44772 643039
rect 45204 641782 45232 684490
rect 45376 669384 45428 669390
rect 45376 669326 45428 669332
rect 45388 667486 45416 669326
rect 45376 667480 45428 667486
rect 45376 667422 45428 667428
rect 45192 641776 45244 641782
rect 45192 641718 45244 641724
rect 45284 640348 45336 640354
rect 45284 640290 45336 640296
rect 45098 640248 45154 640257
rect 45098 640183 45154 640192
rect 44192 624294 44404 624322
rect 44468 634766 44588 634794
rect 44652 635446 44772 635474
rect 44192 623914 44220 624294
rect 44468 624102 44496 634766
rect 44456 624096 44508 624102
rect 44456 624038 44508 624044
rect 44192 623886 44404 623914
rect 43994 623384 44050 623393
rect 43994 623319 44050 623328
rect 44178 622160 44234 622169
rect 44178 622095 44234 622104
rect 44192 616826 44220 622095
rect 44376 619682 44404 623886
rect 44364 619676 44416 619682
rect 44364 619618 44416 619624
rect 44180 616820 44232 616826
rect 44180 616762 44232 616768
rect 44088 615460 44140 615466
rect 44088 615402 44140 615408
rect 44100 614122 44128 615402
rect 44100 614094 44220 614122
rect 44192 613986 44220 614094
rect 44192 613958 44312 613986
rect 44086 613864 44142 613873
rect 44086 613799 44142 613808
rect 43812 612604 43864 612610
rect 43812 612546 43864 612552
rect 44100 612406 44128 613799
rect 44088 612400 44140 612406
rect 43640 612326 43944 612354
rect 44088 612342 44140 612348
rect 43916 612270 43944 612326
rect 43904 612264 43956 612270
rect 43764 612232 43820 612241
rect 43904 612206 43956 612212
rect 43764 612167 43766 612176
rect 43818 612167 43820 612176
rect 43766 612138 43818 612144
rect 44086 612096 44142 612105
rect 44086 612031 44088 612040
rect 44140 612031 44142 612040
rect 44088 612002 44140 612008
rect 43994 611824 44050 611833
rect 43994 611759 43996 611768
rect 44048 611759 44050 611768
rect 43996 611730 44048 611736
rect 44088 611584 44140 611590
rect 44086 611552 44088 611561
rect 44140 611552 44142 611561
rect 44284 611538 44312 613958
rect 44456 612264 44508 612270
rect 44456 612206 44508 612212
rect 44284 611510 44358 611538
rect 44086 611487 44142 611496
rect 43456 611386 44251 611402
rect 43456 611380 44263 611386
rect 43456 611374 44211 611380
rect 44211 611322 44263 611328
rect 44330 611182 44358 611510
rect 44468 611454 44496 612206
rect 44456 611448 44508 611454
rect 44456 611390 44508 611396
rect 44318 611176 44370 611182
rect 44318 611118 44370 611124
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 35806 601760 35862 601769
rect 35806 601695 35808 601704
rect 35860 601695 35862 601704
rect 36544 601724 36596 601730
rect 35808 601666 35860 601672
rect 36544 601666 36596 601672
rect 33046 595402 33102 595411
rect 33046 595337 33102 595346
rect 35438 595402 35494 595411
rect 35438 595337 35494 595346
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585818 31064 594351
rect 33060 587178 33088 595337
rect 33782 593600 33838 593609
rect 33782 593535 33838 593544
rect 33048 587172 33100 587178
rect 33048 587114 33100 587120
rect 33796 585954 33824 593535
rect 35452 587314 35480 595337
rect 36556 592958 36584 601666
rect 38566 601352 38622 601361
rect 38566 601287 38622 601296
rect 38580 594318 38608 601287
rect 39946 600944 40002 600953
rect 39946 600879 40002 600888
rect 39960 595814 39988 600879
rect 44652 600545 44680 635446
rect 44914 630728 44970 630737
rect 44914 630663 44970 630672
rect 44928 611182 44956 630663
rect 44916 611176 44968 611182
rect 44916 611118 44968 611124
rect 44638 600536 44694 600545
rect 44638 600471 44694 600480
rect 44914 600128 44970 600137
rect 44914 600063 44970 600072
rect 42982 597680 43038 597689
rect 42982 597615 43038 597624
rect 42996 597446 43024 597615
rect 42984 597440 43036 597446
rect 42984 597382 43036 597388
rect 42984 597032 43036 597038
rect 42984 596974 43036 596980
rect 43166 597000 43222 597009
rect 42614 596864 42670 596873
rect 42614 596799 42670 596808
rect 42338 596048 42394 596057
rect 42338 595983 42394 595992
rect 39948 595808 40000 595814
rect 41696 595808 41748 595814
rect 39948 595750 40000 595756
rect 41694 595776 41696 595785
rect 41748 595776 41750 595785
rect 41694 595711 41750 595720
rect 39302 594824 39358 594833
rect 39302 594759 39358 594768
rect 38568 594312 38620 594318
rect 38568 594254 38620 594260
rect 36544 592952 36596 592958
rect 36544 592894 36596 592900
rect 35440 587308 35492 587314
rect 35440 587250 35492 587256
rect 33784 585948 33836 585954
rect 33784 585890 33836 585896
rect 31024 585812 31076 585818
rect 31024 585754 31076 585760
rect 39316 585177 39344 594759
rect 41604 594312 41656 594318
rect 41786 594280 41842 594289
rect 41656 594260 41786 594266
rect 41604 594254 41786 594260
rect 41616 594238 41786 594254
rect 41786 594215 41842 594224
rect 41696 592952 41748 592958
rect 41694 592920 41696 592929
rect 41748 592920 41750 592929
rect 41694 592855 41750 592864
rect 42352 592034 42380 595983
rect 42352 592006 42472 592034
rect 41234 589656 41290 589665
rect 41234 589591 41290 589600
rect 40682 587344 40738 587353
rect 40682 587279 40684 587288
rect 40736 587279 40738 587288
rect 40684 587250 40736 587256
rect 40130 585984 40186 585993
rect 40130 585919 40132 585928
rect 40184 585919 40186 585928
rect 40132 585890 40184 585896
rect 41248 585857 41276 589591
rect 41512 587172 41564 587178
rect 41512 587114 41564 587120
rect 41234 585848 41290 585857
rect 40592 585812 40644 585818
rect 41234 585783 41290 585792
rect 40592 585754 40644 585760
rect 39302 585168 39358 585177
rect 39302 585103 39358 585112
rect 40604 584633 40632 585754
rect 40590 584624 40646 584633
rect 40590 584559 40646 584568
rect 41524 584474 41552 587114
rect 42154 585848 42210 585857
rect 42210 585806 42380 585834
rect 42154 585783 42210 585792
rect 41524 584446 42288 584474
rect 42260 583454 42288 584446
rect 42182 583426 42288 583454
rect 42352 582706 42380 585806
rect 42168 582678 42380 582706
rect 42168 582249 42196 582678
rect 42444 582298 42472 592006
rect 42628 587625 42656 596799
rect 42614 587616 42670 587625
rect 42614 587551 42670 587560
rect 42706 587344 42762 587353
rect 42762 587302 42932 587330
rect 42706 587279 42762 587288
rect 42706 584624 42762 584633
rect 42706 584559 42762 584568
rect 42720 584474 42748 584559
rect 42352 582270 42472 582298
rect 42628 584446 42748 584474
rect 42154 581904 42210 581913
rect 42154 581839 42210 581848
rect 42168 581604 42196 581839
rect 42168 580689 42196 580961
rect 42154 580680 42210 580689
rect 42154 580615 42210 580624
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42352 579614 42380 582270
rect 42352 579586 42472 579614
rect 42182 579107 42288 579135
rect 42062 578776 42118 578785
rect 42062 578711 42118 578720
rect 42076 578544 42104 578711
rect 42260 578513 42288 579107
rect 42246 578504 42302 578513
rect 42246 578439 42302 578448
rect 42062 578096 42118 578105
rect 42062 578031 42118 578040
rect 42076 577932 42104 578031
rect 42248 577856 42300 577862
rect 41786 577824 41842 577833
rect 42248 577798 42300 577804
rect 41786 577759 41842 577768
rect 41800 577281 41828 577759
rect 42260 576858 42288 577798
rect 42168 576830 42288 576858
rect 42168 576708 42196 576830
rect 42246 575648 42302 575657
rect 42246 575583 42302 575592
rect 41786 574696 41842 574705
rect 41786 574631 41842 574640
rect 41800 574260 41828 574631
rect 42260 573866 42288 575583
rect 42168 573838 42288 573866
rect 42168 573580 42196 573838
rect 42156 573504 42208 573510
rect 42156 573446 42208 573452
rect 42168 572968 42196 573446
rect 42444 573322 42472 579586
rect 42628 577946 42656 584446
rect 42904 579614 42932 587302
rect 42536 577918 42656 577946
rect 42720 579586 42932 579614
rect 42536 573594 42564 577918
rect 42720 577862 42748 579586
rect 42708 577856 42760 577862
rect 42708 577798 42760 577804
rect 42536 573566 42656 573594
rect 42628 573510 42656 573566
rect 42616 573504 42668 573510
rect 42616 573446 42668 573452
rect 42352 573294 42472 573322
rect 42352 572438 42380 573294
rect 42614 572792 42670 572801
rect 42614 572727 42670 572736
rect 42168 572370 42196 572424
rect 42260 572410 42380 572438
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42062 571568 42118 571577
rect 42062 571503 42118 571512
rect 42076 571282 42104 571503
rect 42430 571432 42486 571441
rect 42430 571367 42486 571376
rect 42076 571254 42380 571282
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42352 569310 42380 571254
rect 42168 569242 42196 569296
rect 42260 569282 42380 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42444 568766 42472 571367
rect 42628 570994 42656 572727
rect 42616 570988 42668 570994
rect 42616 570930 42668 570936
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 42996 567194 43024 596974
rect 43166 596935 43222 596944
rect 43180 582374 43208 596935
rect 44362 593192 44418 593201
rect 44362 593127 44418 593136
rect 44178 591968 44234 591977
rect 44178 591903 44234 591912
rect 43350 591560 43406 591569
rect 43350 591495 43406 591504
rect 42812 567166 43024 567194
rect 43088 582346 43208 582374
rect 43364 582374 43392 591495
rect 43626 590336 43682 590345
rect 43626 590271 43682 590280
rect 43364 582346 43484 582374
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 42338 558104 42394 558113
rect 42338 558039 42394 558048
rect 40038 553408 40094 553417
rect 40038 553343 40094 553352
rect 40958 553408 41014 553417
rect 40958 553343 41014 553352
rect 34426 551984 34482 551993
rect 34426 551919 34482 551928
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 31760 547402 31812 547408
rect 34440 544406 34468 551919
rect 40052 551002 40080 553343
rect 40040 550996 40092 551002
rect 40040 550938 40092 550944
rect 40972 549794 41000 553343
rect 42352 552673 42380 558039
rect 42812 554849 42840 567166
rect 43088 556481 43116 582346
rect 43074 556472 43130 556481
rect 43074 556407 43130 556416
rect 42798 554840 42854 554849
rect 42798 554775 42854 554784
rect 42338 552664 42394 552673
rect 42338 552599 42394 552608
rect 42982 552392 43038 552401
rect 42982 552327 43038 552336
rect 42798 551168 42854 551177
rect 42798 551103 42854 551112
rect 41696 550996 41748 551002
rect 41748 550956 42380 550984
rect 41696 550938 41748 550944
rect 41878 550352 41934 550361
rect 41878 550287 41934 550296
rect 40972 549766 41184 549794
rect 41156 547346 41184 549766
rect 41696 547460 41748 547466
rect 41696 547402 41748 547408
rect 41156 547318 41368 547346
rect 41340 546417 41368 547318
rect 41326 546408 41382 546417
rect 41326 546343 41382 546352
rect 34428 544400 34480 544406
rect 34428 544342 34480 544348
rect 41328 544400 41380 544406
rect 41328 544342 41380 544348
rect 41340 541385 41368 544342
rect 41708 543538 41736 547402
rect 41892 545737 41920 550287
rect 42062 549944 42118 549953
rect 42062 549879 42118 549888
rect 41878 545728 41934 545737
rect 41878 545663 41934 545672
rect 42076 545465 42104 549879
rect 42352 549254 42380 550956
rect 42352 549226 42656 549254
rect 42062 545456 42118 545465
rect 42062 545391 42118 545400
rect 41708 543510 42380 543538
rect 41326 541376 41382 541385
rect 41326 541311 41382 541320
rect 42352 540818 42380 543510
rect 42260 540790 42380 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 41800 540260 41828 540631
rect 42260 539050 42288 540790
rect 42628 540682 42656 549226
rect 42182 539022 42288 539050
rect 42352 540654 42656 540682
rect 42352 538438 42380 540654
rect 42522 539608 42578 539617
rect 42522 539543 42578 539552
rect 42168 538370 42196 538424
rect 42260 538410 42380 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42536 538234 42564 539543
rect 42352 538206 42564 538234
rect 42168 537798 42288 537826
rect 42168 537744 42196 537798
rect 42260 537758 42288 537798
rect 42352 537758 42380 538206
rect 42614 538112 42670 538121
rect 42812 538098 42840 551103
rect 42996 550634 43024 552327
rect 42904 550606 43024 550634
rect 42904 540974 42932 550606
rect 43166 549536 43222 549545
rect 43166 549471 43222 549480
rect 42904 540946 43024 540974
rect 42996 538218 43024 540946
rect 42984 538212 43036 538218
rect 42984 538154 43036 538160
rect 42812 538070 43024 538098
rect 42614 538047 42670 538056
rect 42260 537730 42380 537758
rect 42430 537432 42486 537441
rect 42430 537367 42486 537376
rect 41786 537024 41842 537033
rect 41786 536959 41842 536968
rect 41800 536588 41828 536959
rect 42246 536480 42302 536489
rect 42246 536415 42302 536424
rect 42076 535673 42104 535908
rect 42062 535664 42118 535673
rect 42062 535599 42118 535608
rect 42260 535514 42288 536415
rect 42168 535486 42288 535514
rect 42168 535364 42196 535486
rect 42444 534766 42472 537367
rect 42628 536874 42656 538047
rect 42800 537940 42852 537946
rect 42800 537882 42852 537888
rect 42812 537758 42840 537882
rect 42168 534698 42196 534752
rect 42260 534738 42472 534766
rect 42536 536846 42656 536874
rect 42720 537730 42840 537758
rect 42260 534698 42288 534738
rect 42168 534670 42288 534698
rect 42536 534290 42564 536846
rect 42444 534262 42564 534290
rect 42444 534086 42472 534262
rect 42182 534058 42472 534086
rect 42720 533610 42748 537730
rect 42536 533582 42748 533610
rect 42536 533542 42564 533582
rect 42182 533514 42564 533542
rect 42706 532808 42762 532817
rect 42432 532772 42484 532778
rect 42706 532743 42762 532752
rect 42432 532714 42484 532720
rect 42444 531059 42472 532714
rect 42182 531031 42472 531059
rect 42720 530890 42748 532743
rect 42444 530862 42748 530890
rect 42444 530414 42472 530862
rect 42614 530768 42670 530777
rect 42614 530703 42670 530712
rect 42168 530346 42196 530400
rect 42352 530386 42472 530414
rect 42352 530346 42380 530386
rect 42168 530318 42380 530346
rect 42156 530120 42208 530126
rect 42156 530062 42208 530068
rect 42168 529757 42196 530062
rect 42430 529544 42486 529553
rect 42430 529479 42486 529488
rect 41800 529009 41828 529205
rect 41786 529000 41842 529009
rect 41786 528935 41842 528944
rect 42246 528864 42302 528873
rect 42246 528799 42302 528808
rect 42064 527808 42116 527814
rect 42064 527750 42116 527756
rect 42076 527340 42104 527750
rect 42260 526810 42288 528799
rect 42168 526782 42288 526810
rect 42168 526728 42196 526782
rect 42444 526091 42472 529479
rect 42628 527814 42656 530703
rect 42996 530126 43024 538070
rect 43180 532778 43208 549471
rect 43168 532772 43220 532778
rect 43168 532714 43220 532720
rect 42984 530120 43036 530126
rect 42984 530062 43036 530068
rect 42616 527808 42668 527814
rect 42616 527750 42668 527756
rect 42614 527232 42670 527241
rect 42614 527167 42670 527176
rect 42182 526063 42472 526091
rect 42168 525558 42288 525586
rect 42168 525504 42196 525558
rect 42260 525518 42288 525558
rect 42628 525518 42656 527167
rect 42260 525490 42656 525518
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 35806 430128 35862 430137
rect 35806 430063 35862 430072
rect 35820 429214 35848 430063
rect 35808 429208 35860 429214
rect 35808 429150 35860 429156
rect 41696 429208 41748 429214
rect 41696 429150 41748 429156
rect 41708 427122 41736 429150
rect 41970 427136 42026 427145
rect 41708 427094 41970 427122
rect 41970 427071 42026 427080
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 41142 425640 41198 425649
rect 41142 425575 41198 425584
rect 40958 425232 41014 425241
rect 40958 425167 41014 425176
rect 32034 424416 32090 424425
rect 32034 424351 32090 424360
rect 32048 416226 32076 424351
rect 40972 424318 41000 425167
rect 40960 424312 41012 424318
rect 40960 424254 41012 424260
rect 41156 418849 41184 425575
rect 41340 425134 41368 425983
rect 41328 425128 41380 425134
rect 41328 425070 41380 425076
rect 41696 425128 41748 425134
rect 41748 425076 42104 425082
rect 41696 425070 42104 425076
rect 41708 425054 42104 425070
rect 41512 424312 41564 424318
rect 41878 424280 41934 424289
rect 41564 424260 41878 424266
rect 41512 424254 41878 424260
rect 41524 424238 41878 424254
rect 41878 424215 41934 424224
rect 41142 418840 41198 418849
rect 41142 418775 41198 418784
rect 42076 418154 42104 425054
rect 42798 423600 42854 423609
rect 42798 423535 42854 423544
rect 42522 419928 42578 419937
rect 42522 419863 42578 419872
rect 42076 418126 42380 418154
rect 32036 416220 32088 416226
rect 32036 416162 32088 416168
rect 41696 416220 41748 416226
rect 41696 416162 41748 416168
rect 41708 416106 41736 416162
rect 41708 416078 42288 416106
rect 42260 413114 42288 416078
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42352 411074 42380 418126
rect 42536 411913 42564 419863
rect 42522 411904 42578 411913
rect 42522 411839 42578 411848
rect 42168 411046 42380 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 41970 408096 42026 408105
rect 41970 408031 42026 408040
rect 41984 407796 42012 408031
rect 42168 407946 42196 408340
rect 42168 407918 42288 407946
rect 42260 407674 42288 407918
rect 42444 407833 42472 410162
rect 42430 407824 42486 407833
rect 42430 407759 42486 407768
rect 42260 407646 42472 407674
rect 42246 407552 42302 407561
rect 42246 407487 42302 407496
rect 42260 407130 42288 407487
rect 42182 407102 42288 407130
rect 42062 406736 42118 406745
rect 42062 406671 42118 406680
rect 42076 406504 42104 406671
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 42444 405657 42472 407646
rect 42246 405648 42302 405657
rect 42246 405583 42302 405592
rect 42430 405648 42486 405657
rect 42430 405583 42486 405592
rect 42260 403458 42288 405583
rect 42182 403430 42288 403458
rect 42812 402974 42840 423535
rect 43258 420744 43314 420753
rect 43258 420679 43314 420688
rect 43074 419520 43130 419529
rect 43074 419455 43130 419464
rect 42536 402946 42840 402974
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42536 402166 42564 402946
rect 42182 402138 42564 402166
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 42430 400208 42486 400217
rect 42430 400143 42486 400152
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 42444 399135 42472 400143
rect 42182 399107 42472 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 42168 395729 42196 397936
rect 42154 395720 42210 395729
rect 42154 395655 42210 395664
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41142 387152 41198 387161
rect 41142 387087 41198 387096
rect 40774 385928 40830 385937
rect 40774 385863 40830 385872
rect 40788 381449 40816 385863
rect 41156 381857 41184 387087
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41340 385937 41368 386679
rect 41326 385928 41382 385937
rect 41326 385863 41382 385872
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382294 41368 382599
rect 41328 382288 41380 382294
rect 41328 382230 41380 382236
rect 41696 382288 41748 382294
rect 41696 382230 41748 382236
rect 40958 381848 41014 381857
rect 40958 381783 41014 381792
rect 41142 381848 41198 381857
rect 41142 381783 41198 381792
rect 40222 381440 40278 381449
rect 40222 381375 40278 381384
rect 40774 381440 40830 381449
rect 40774 381375 40830 381384
rect 35162 381032 35218 381041
rect 35162 380967 35218 380976
rect 33782 379808 33838 379817
rect 33782 379743 33838 379752
rect 33796 371929 33824 379743
rect 33782 371920 33838 371929
rect 35176 371890 35204 380967
rect 37922 380216 37978 380225
rect 37922 380151 37978 380160
rect 35808 379704 35860 379710
rect 35808 379646 35860 379652
rect 35820 379409 35848 379646
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 35820 374649 35848 376479
rect 35806 374640 35862 374649
rect 35806 374575 35862 374584
rect 37936 372745 37964 380151
rect 40236 378078 40264 381375
rect 40972 379817 41000 381783
rect 40958 379808 41014 379817
rect 40958 379743 41014 379752
rect 40592 379704 40644 379710
rect 40592 379646 40644 379652
rect 40604 379409 40632 379646
rect 41708 379514 41736 382230
rect 41708 379486 42380 379514
rect 40590 379400 40646 379409
rect 40590 379335 40646 379344
rect 40224 378072 40276 378078
rect 40224 378014 40276 378020
rect 41696 378072 41748 378078
rect 41748 378020 42104 378026
rect 41696 378014 42104 378020
rect 41708 378010 42104 378014
rect 41708 378004 42116 378010
rect 41708 377998 42064 378004
rect 42064 377946 42116 377952
rect 37922 372736 37978 372745
rect 37922 372671 37978 372680
rect 33782 371855 33838 371864
rect 35164 371884 35216 371890
rect 35164 371826 35216 371832
rect 41696 371884 41748 371890
rect 41696 371826 41748 371832
rect 41708 371770 41736 371826
rect 41708 371742 42288 371770
rect 42260 369458 42288 371742
rect 42182 369430 42288 369458
rect 41786 368520 41842 368529
rect 41786 368455 41842 368464
rect 41800 368249 41828 368455
rect 42352 367622 42380 379486
rect 42890 379400 42946 379409
rect 42890 379335 42946 379344
rect 42708 378004 42760 378010
rect 42708 377946 42760 377952
rect 42182 367594 42380 367622
rect 42182 366947 42288 366975
rect 42062 366208 42118 366217
rect 42062 366143 42118 366152
rect 42076 365772 42104 366143
rect 42260 365294 42288 366947
rect 42248 365288 42300 365294
rect 42248 365230 42300 365236
rect 42182 365107 42472 365135
rect 42248 364948 42300 364954
rect 42248 364890 42300 364896
rect 42062 364848 42118 364857
rect 42062 364783 42118 364792
rect 42076 364548 42104 364783
rect 42260 364342 42288 364890
rect 42248 364336 42300 364342
rect 42248 364278 42300 364284
rect 42246 364168 42302 364177
rect 42246 364103 42302 364112
rect 42260 363950 42288 364103
rect 42182 363922 42288 363950
rect 41786 363760 41842 363769
rect 41786 363695 41842 363704
rect 41800 363256 41828 363695
rect 42444 363066 42472 365107
rect 42720 364334 42748 377946
rect 42904 366217 42932 379335
rect 42890 366208 42946 366217
rect 42890 366143 42946 366152
rect 42260 363038 42472 363066
rect 42536 364306 42748 364334
rect 42260 362953 42288 363038
rect 42246 362944 42302 362953
rect 42246 362879 42302 362888
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362726 42564 364306
rect 42708 364200 42760 364206
rect 42708 364142 42760 364148
rect 42720 363225 42748 364142
rect 42706 363216 42762 363225
rect 42706 363151 42762 363160
rect 42260 362698 42564 362726
rect 42430 361584 42486 361593
rect 42430 361519 42486 361528
rect 42444 360278 42472 361519
rect 42168 360210 42196 360264
rect 42260 360250 42472 360278
rect 42260 360210 42288 360250
rect 42168 360182 42288 360210
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 41800 359584 41828 360023
rect 41786 359272 41842 359281
rect 41786 359207 41842 359216
rect 41800 358972 41828 359207
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 42168 356538 42196 356592
rect 42260 356578 42472 356606
rect 42260 356538 42288 356578
rect 42168 356510 42288 356538
rect 41786 356144 41842 356153
rect 41786 356079 41842 356088
rect 41800 355912 41828 356079
rect 42168 355042 42196 355300
rect 42168 355014 42288 355042
rect 42168 353297 42196 354725
rect 42260 353920 42288 355014
rect 42444 354385 42472 356578
rect 42430 354376 42486 354385
rect 42430 354311 42486 354320
rect 43088 353977 43116 419455
rect 43074 353968 43130 353977
rect 42260 353892 42380 353920
rect 43074 353903 43130 353912
rect 42154 353288 42210 353297
rect 42154 353223 42210 353232
rect 42352 353025 42380 353892
rect 43272 353705 43300 420679
rect 43456 354674 43484 582346
rect 43640 354929 43668 590271
rect 44192 578785 44220 591903
rect 44178 578776 44234 578785
rect 44178 578711 44234 578720
rect 44376 578105 44404 593127
rect 44638 580680 44694 580689
rect 44638 580615 44694 580624
rect 44362 578096 44418 578105
rect 44362 578031 44418 578040
rect 44652 575482 44680 580615
rect 44640 575476 44692 575482
rect 44640 575418 44692 575424
rect 44928 558793 44956 600063
rect 45112 598913 45140 640183
rect 45098 598904 45154 598913
rect 45098 598839 45154 598848
rect 45098 598496 45154 598505
rect 45098 598431 45154 598440
rect 44914 558784 44970 558793
rect 44914 558719 44970 558728
rect 44546 556880 44602 556889
rect 44546 556815 44602 556824
rect 44270 556064 44326 556073
rect 44270 555999 44326 556008
rect 43810 548312 43866 548321
rect 43810 548247 43866 548256
rect 43824 355201 43852 548247
rect 43994 547088 44050 547097
rect 43994 547023 44050 547032
rect 43810 355192 43866 355201
rect 43810 355127 43866 355136
rect 43626 354920 43682 354929
rect 43626 354855 43682 354864
rect 43456 354646 43760 354674
rect 43732 354634 43760 354646
rect 44008 354634 44036 547023
rect 44284 428913 44312 555999
rect 44560 429729 44588 556815
rect 45112 555665 45140 598431
rect 45296 598097 45324 640290
rect 45572 612105 45600 763263
rect 46216 743782 46244 772958
rect 46204 743776 46256 743782
rect 46204 743718 46256 743724
rect 60016 742422 60044 774182
rect 651470 774143 651472 774152
rect 651524 774143 651526 774152
rect 651472 774114 651524 774120
rect 651472 773832 651524 773838
rect 651472 773774 651524 773780
rect 651484 773401 651512 773774
rect 651470 773392 651526 773401
rect 651470 773327 651526 773336
rect 61384 772880 61436 772886
rect 61384 772822 61436 772828
rect 61396 747046 61424 772822
rect 62764 755540 62816 755546
rect 62764 755482 62816 755488
rect 62776 747697 62804 755482
rect 62762 747688 62818 747697
rect 62762 747623 62818 747632
rect 61384 747040 61436 747046
rect 61384 746982 61436 746988
rect 62396 747040 62448 747046
rect 62396 746982 62448 746988
rect 62120 746564 62172 746570
rect 62120 746506 62172 746512
rect 62132 746201 62160 746506
rect 62118 746192 62174 746201
rect 62118 746127 62174 746136
rect 62118 744152 62174 744161
rect 62118 744087 62174 744096
rect 62132 743918 62160 744087
rect 62120 743912 62172 743918
rect 62120 743854 62172 743860
rect 62120 743776 62172 743782
rect 62118 743744 62120 743753
rect 62172 743744 62174 743753
rect 62118 743679 62174 743688
rect 60004 742416 60056 742422
rect 62120 742416 62172 742422
rect 60004 742358 60056 742364
rect 62118 742384 62120 742393
rect 62172 742384 62174 742393
rect 62118 742319 62174 742328
rect 62408 741849 62436 746982
rect 62394 741840 62450 741849
rect 62394 741775 62450 741784
rect 652036 736234 652064 776999
rect 653416 775334 653444 790774
rect 655520 781108 655572 781114
rect 655520 781050 655572 781056
rect 655152 778524 655204 778530
rect 655152 778466 655204 778472
rect 653404 775328 653456 775334
rect 653404 775270 653456 775276
rect 655164 773838 655192 778466
rect 655532 774178 655560 781050
rect 660304 777640 660356 777646
rect 660304 777582 660356 777588
rect 655520 774172 655572 774178
rect 655520 774114 655572 774120
rect 655152 773832 655204 773838
rect 655152 773774 655204 773780
rect 652024 736228 652076 736234
rect 652024 736170 652076 736176
rect 653404 736228 653456 736234
rect 653404 736170 653456 736176
rect 651470 734224 651526 734233
rect 651470 734159 651526 734168
rect 651484 733446 651512 734159
rect 651472 733440 651524 733446
rect 651472 733382 651524 733388
rect 651470 733000 651526 733009
rect 651470 732935 651526 732944
rect 651484 732834 651512 732935
rect 651472 732828 651524 732834
rect 651472 732770 651524 732776
rect 651470 731776 651526 731785
rect 651470 731711 651526 731720
rect 651484 731474 651512 731711
rect 651472 731468 651524 731474
rect 651472 731410 651524 731416
rect 651472 731332 651524 731338
rect 651472 731274 651524 731280
rect 61384 731196 61436 731202
rect 61384 731138 61436 731144
rect 46202 730280 46258 730289
rect 46202 730215 46258 730224
rect 46216 698222 46244 730215
rect 47214 721168 47270 721177
rect 47214 721103 47270 721112
rect 47030 719944 47086 719953
rect 47030 719879 47086 719888
rect 46204 698216 46256 698222
rect 46204 698158 46256 698164
rect 45744 667956 45796 667962
rect 45744 667898 45796 667904
rect 45756 665961 45784 667898
rect 45742 665952 45798 665961
rect 45742 665887 45798 665896
rect 45558 612096 45614 612105
rect 45558 612031 45614 612040
rect 47044 611833 47072 719879
rect 47030 611824 47086 611833
rect 47030 611759 47086 611768
rect 47228 611561 47256 721103
rect 50344 712156 50396 712162
rect 50344 712098 50396 712104
rect 50356 705158 50384 712098
rect 50344 705152 50396 705158
rect 50344 705094 50396 705100
rect 61396 699689 61424 731138
rect 651484 731105 651512 731274
rect 651470 731096 651526 731105
rect 651470 731031 651526 731040
rect 651472 730040 651524 730046
rect 651472 729982 651524 729988
rect 651484 729881 651512 729982
rect 651470 729872 651526 729881
rect 651470 729807 651526 729816
rect 62764 729360 62816 729366
rect 62764 729302 62816 729308
rect 62120 705152 62172 705158
rect 62120 705094 62172 705100
rect 62132 704449 62160 705094
rect 62118 704440 62174 704449
rect 62118 704375 62174 704384
rect 62120 703792 62172 703798
rect 62120 703734 62172 703740
rect 62132 703361 62160 703734
rect 62118 703352 62174 703361
rect 62118 703287 62174 703296
rect 62210 701312 62266 701321
rect 62210 701247 62266 701256
rect 62224 701078 62252 701247
rect 62212 701072 62264 701078
rect 62212 701014 62264 701020
rect 62776 700913 62804 729302
rect 651472 728544 651524 728550
rect 651470 728512 651472 728521
rect 651524 728512 651526 728521
rect 651470 728447 651526 728456
rect 653416 716310 653444 736170
rect 657544 735616 657596 735622
rect 657544 735558 657596 735564
rect 654784 734188 654836 734194
rect 654784 734130 654836 734136
rect 654796 728550 654824 734130
rect 657556 730046 657584 735558
rect 658924 731468 658976 731474
rect 658924 731410 658976 731416
rect 657544 730040 657596 730046
rect 657544 729982 657596 729988
rect 654784 728544 654836 728550
rect 654784 728486 654836 728492
rect 653404 716304 653456 716310
rect 653404 716246 653456 716252
rect 654784 701072 654836 701078
rect 654784 701014 654836 701020
rect 62762 700904 62818 700913
rect 62762 700839 62818 700848
rect 61382 699680 61438 699689
rect 61382 699615 61438 699624
rect 62120 698216 62172 698222
rect 62118 698184 62120 698193
rect 62172 698184 62174 698193
rect 62118 698119 62174 698128
rect 651654 689480 651710 689489
rect 651654 689415 651710 689424
rect 651470 688800 651526 688809
rect 651470 688735 651526 688744
rect 651484 687954 651512 688735
rect 651668 688702 651696 689415
rect 652760 688832 652812 688838
rect 652760 688774 652812 688780
rect 651656 688696 651708 688702
rect 651656 688638 651708 688644
rect 651472 687948 651524 687954
rect 651472 687890 651524 687896
rect 652022 687304 652078 687313
rect 61384 687268 61436 687274
rect 652022 687239 652078 687248
rect 61384 687210 61436 687216
rect 53104 669384 53156 669390
rect 53104 669326 53156 669332
rect 53116 660958 53144 669326
rect 57244 667956 57296 667962
rect 57244 667898 57296 667904
rect 53104 660952 53156 660958
rect 53104 660894 53156 660900
rect 57256 659598 57284 667898
rect 57244 659592 57296 659598
rect 57244 659534 57296 659540
rect 61396 656577 61424 687210
rect 651472 687200 651524 687206
rect 651472 687142 651524 687148
rect 651484 686905 651512 687142
rect 651470 686896 651526 686905
rect 651470 686831 651526 686840
rect 62764 686520 62816 686526
rect 62764 686462 62816 686468
rect 62120 660952 62172 660958
rect 62118 660920 62120 660929
rect 62172 660920 62174 660929
rect 62118 660855 62174 660864
rect 62120 659592 62172 659598
rect 62118 659560 62120 659569
rect 62172 659560 62174 659569
rect 62118 659495 62174 659504
rect 62118 658336 62174 658345
rect 62118 658271 62174 658280
rect 62132 657558 62160 658271
rect 62776 657665 62804 686462
rect 651472 685568 651524 685574
rect 651472 685510 651524 685516
rect 651484 685273 651512 685510
rect 651470 685264 651526 685273
rect 651470 685199 651526 685208
rect 62762 657656 62818 657665
rect 62762 657591 62818 657600
rect 62120 657552 62172 657558
rect 62120 657494 62172 657500
rect 61382 656568 61438 656577
rect 61382 656503 61438 656512
rect 62120 655512 62172 655518
rect 62120 655454 62172 655460
rect 62132 655353 62160 655454
rect 62118 655344 62174 655353
rect 62118 655279 62174 655288
rect 652036 645182 652064 687239
rect 652574 684448 652630 684457
rect 652772 684434 652800 688774
rect 654796 687206 654824 701014
rect 656808 690056 656860 690062
rect 656808 689998 656860 690004
rect 654784 687200 654836 687206
rect 654784 687142 654836 687148
rect 656820 685574 656848 689998
rect 656808 685568 656860 685574
rect 656808 685510 656860 685516
rect 652630 684406 652800 684434
rect 652574 684383 652630 684392
rect 658936 669526 658964 731410
rect 660316 714882 660344 777582
rect 668400 775600 668452 775606
rect 668400 775542 668452 775548
rect 661684 732828 661736 732834
rect 661684 732770 661736 732776
rect 660304 714876 660356 714882
rect 660304 714818 660356 714824
rect 660304 688696 660356 688702
rect 660304 688638 660356 688644
rect 658924 669520 658976 669526
rect 658924 669462 658976 669468
rect 653404 655580 653456 655586
rect 653404 655522 653456 655528
rect 652024 645176 652076 645182
rect 652024 645118 652076 645124
rect 60004 644496 60056 644502
rect 60004 644438 60056 644444
rect 60016 612678 60044 644438
rect 651470 643240 651526 643249
rect 651470 643175 651526 643184
rect 61384 643136 61436 643142
rect 61384 643078 61436 643084
rect 61396 613873 61424 643078
rect 651484 642394 651512 643175
rect 62764 642388 62816 642394
rect 62764 642330 62816 642336
rect 651472 642388 651524 642394
rect 651472 642330 651524 642336
rect 62120 616820 62172 616826
rect 62120 616762 62172 616768
rect 62132 616593 62160 616762
rect 62118 616584 62174 616593
rect 62118 616519 62174 616528
rect 62118 614680 62174 614689
rect 62118 614615 62174 614624
rect 62132 614174 62160 614615
rect 62120 614168 62172 614174
rect 62120 614110 62172 614116
rect 61382 613864 61438 613873
rect 61382 613799 61438 613808
rect 60004 612672 60056 612678
rect 62120 612672 62172 612678
rect 60004 612614 60056 612620
rect 62118 612640 62120 612649
rect 62172 612640 62174 612649
rect 62118 612575 62174 612584
rect 62776 612105 62804 642330
rect 652022 641880 652078 641889
rect 652022 641815 652078 641824
rect 651470 640792 651526 640801
rect 651470 640727 651526 640736
rect 651484 640354 651512 640727
rect 651472 640348 651524 640354
rect 651472 640290 651524 640296
rect 651380 640144 651432 640150
rect 651378 640112 651380 640121
rect 651432 640112 651434 640121
rect 651378 640047 651434 640056
rect 651656 638920 651708 638926
rect 651656 638862 651708 638868
rect 651472 638784 651524 638790
rect 651472 638726 651524 638732
rect 651484 638625 651512 638726
rect 651470 638616 651526 638625
rect 651470 638551 651526 638560
rect 651668 638217 651696 638862
rect 651654 638208 651710 638217
rect 651654 638143 651710 638152
rect 62948 625864 63000 625870
rect 62948 625806 63000 625812
rect 62960 618089 62988 625806
rect 62946 618080 63002 618089
rect 62946 618015 63002 618024
rect 62762 612096 62818 612105
rect 62762 612031 62818 612040
rect 47214 611552 47270 611561
rect 47214 611487 47270 611496
rect 45282 598088 45338 598097
rect 45282 598023 45338 598032
rect 651470 597952 651526 597961
rect 651470 597887 651526 597896
rect 651484 597582 651512 597887
rect 651472 597576 651524 597582
rect 651472 597518 651524 597524
rect 651470 596728 651526 596737
rect 651470 596663 651526 596672
rect 651484 596222 651512 596663
rect 651472 596216 651524 596222
rect 651472 596158 651524 596164
rect 62946 595776 63002 595785
rect 62946 595711 63002 595720
rect 62762 594144 62818 594153
rect 62762 594079 62818 594088
rect 45558 578504 45614 578513
rect 45558 578439 45614 578448
rect 45572 574054 45600 578439
rect 62120 575476 62172 575482
rect 62120 575418 62172 575424
rect 62132 574841 62160 575418
rect 62118 574832 62174 574841
rect 62118 574767 62174 574776
rect 45560 574048 45612 574054
rect 45560 573990 45612 573996
rect 62120 574048 62172 574054
rect 62120 573990 62172 573996
rect 62132 573617 62160 573990
rect 62118 573608 62174 573617
rect 62118 573543 62174 573552
rect 62776 568585 62804 594079
rect 62960 571169 62988 595711
rect 651470 595504 651526 595513
rect 651470 595439 651526 595448
rect 651656 595468 651708 595474
rect 651484 594930 651512 595439
rect 651656 595410 651708 595416
rect 651668 595241 651696 595410
rect 651654 595232 651710 595241
rect 651654 595167 651710 595176
rect 651472 594924 651524 594930
rect 651472 594866 651524 594872
rect 651472 594720 651524 594726
rect 651472 594662 651524 594668
rect 651484 594153 651512 594662
rect 651470 594144 651526 594153
rect 651470 594079 651526 594088
rect 651472 593088 651524 593094
rect 651472 593030 651524 593036
rect 63130 592920 63186 592929
rect 63130 592855 63186 592864
rect 62946 571160 63002 571169
rect 62946 571095 63002 571104
rect 63144 569945 63172 592855
rect 651484 592793 651512 593030
rect 651470 592784 651526 592793
rect 651470 592719 651526 592728
rect 652036 581058 652064 641815
rect 653416 640150 653444 655522
rect 655520 645924 655572 645930
rect 655520 645866 655572 645872
rect 655336 643136 655388 643142
rect 655336 643078 655388 643084
rect 653404 640144 653456 640150
rect 653404 640086 653456 640092
rect 655348 638926 655376 643078
rect 655336 638920 655388 638926
rect 655336 638862 655388 638868
rect 655532 638790 655560 645866
rect 658924 642388 658976 642394
rect 658924 642330 658976 642336
rect 655520 638784 655572 638790
rect 655520 638726 655572 638732
rect 653404 611380 653456 611386
rect 653404 611322 653456 611328
rect 653416 595474 653444 611322
rect 657544 600500 657596 600506
rect 657544 600442 657596 600448
rect 654784 599004 654836 599010
rect 654784 598946 654836 598952
rect 653404 595468 653456 595474
rect 653404 595410 653456 595416
rect 654796 593094 654824 598946
rect 656164 594924 656216 594930
rect 656164 594866 656216 594872
rect 654784 593088 654836 593094
rect 654784 593030 654836 593036
rect 652024 581052 652076 581058
rect 652024 580994 652076 581000
rect 63130 569936 63186 569945
rect 63130 569871 63186 569880
rect 62762 568576 62818 568585
rect 62762 568511 62818 568520
rect 653404 565888 653456 565894
rect 653404 565830 653456 565836
rect 61382 557560 61438 557569
rect 61382 557495 61438 557504
rect 45098 555656 45154 555665
rect 45098 555591 45154 555600
rect 45650 555248 45706 555257
rect 45650 555183 45706 555192
rect 45190 551576 45246 551585
rect 45190 551511 45246 551520
rect 45006 549128 45062 549137
rect 45006 549063 45062 549072
rect 44730 548720 44786 548729
rect 44730 548655 44786 548664
rect 44744 536897 44772 548655
rect 45020 538121 45048 549063
rect 45006 538112 45062 538121
rect 45006 538047 45062 538056
rect 44730 536888 44786 536897
rect 44730 536823 44786 536832
rect 44730 535664 44786 535673
rect 44730 535599 44786 535608
rect 44744 531146 44772 535599
rect 44732 531140 44784 531146
rect 44732 531082 44784 531088
rect 45204 528873 45232 551511
rect 45374 550760 45430 550769
rect 45374 550695 45430 550704
rect 45388 532817 45416 550695
rect 45374 532808 45430 532817
rect 45374 532743 45430 532752
rect 45190 528864 45246 528873
rect 45190 528799 45246 528808
rect 45100 528624 45152 528630
rect 45100 528566 45152 528572
rect 45112 527241 45140 528566
rect 45098 527232 45154 527241
rect 45098 527167 45154 527176
rect 44546 429720 44602 429729
rect 44546 429655 44602 429664
rect 44638 429312 44694 429321
rect 44638 429247 44694 429256
rect 44270 428904 44326 428913
rect 44270 428839 44326 428848
rect 44270 428496 44326 428505
rect 44270 428431 44326 428440
rect 44284 385665 44312 428431
rect 44454 422376 44510 422385
rect 44454 422311 44510 422320
rect 44468 407561 44496 422311
rect 44454 407552 44510 407561
rect 44454 407487 44510 407496
rect 44652 386481 44680 429247
rect 45664 428097 45692 555183
rect 45834 554432 45890 554441
rect 45834 554367 45890 554376
rect 45650 428088 45706 428097
rect 45650 428023 45706 428032
rect 45558 427680 45614 427689
rect 45558 427615 45614 427624
rect 45006 423192 45062 423201
rect 45006 423127 45062 423136
rect 44822 405648 44878 405657
rect 44822 405583 44878 405592
rect 44836 402966 44864 405583
rect 44824 402960 44876 402966
rect 45020 402937 45048 423127
rect 45374 421560 45430 421569
rect 45374 421495 45430 421504
rect 45190 421152 45246 421161
rect 45190 421087 45246 421096
rect 45204 408105 45232 421087
rect 45190 408096 45246 408105
rect 45190 408031 45246 408040
rect 45388 406745 45416 421495
rect 45374 406736 45430 406745
rect 45374 406671 45430 406680
rect 44824 402902 44876 402908
rect 45006 402928 45062 402937
rect 45006 402863 45062 402872
rect 44638 386472 44694 386481
rect 44638 386407 44694 386416
rect 44270 385656 44326 385665
rect 44270 385591 44326 385600
rect 45098 385248 45154 385257
rect 45098 385183 45154 385192
rect 44362 379128 44418 379137
rect 44362 379063 44418 379072
rect 44178 376272 44234 376281
rect 44178 376207 44234 376216
rect 44192 359666 44220 376207
rect 44376 364177 44404 379063
rect 44546 378720 44602 378729
rect 44546 378655 44602 378664
rect 44362 364168 44418 364177
rect 44362 364103 44418 364112
rect 44560 361593 44588 378655
rect 44730 377904 44786 377913
rect 44730 377839 44786 377848
rect 44744 364857 44772 377839
rect 44914 377496 44970 377505
rect 44914 377431 44970 377440
rect 44730 364848 44786 364857
rect 44730 364783 44786 364792
rect 44928 364334 44956 377431
rect 45112 369854 45140 385183
rect 45572 384849 45600 427615
rect 45848 427417 45876 554367
rect 60002 539608 60058 539617
rect 60002 539543 60058 539552
rect 60016 531282 60044 539543
rect 60004 531276 60056 531282
rect 60004 531218 60056 531224
rect 61396 527105 61424 557495
rect 63406 556744 63462 556753
rect 63406 556679 63462 556688
rect 62946 552664 63002 552673
rect 62946 552599 63002 552608
rect 62118 531312 62174 531321
rect 62118 531247 62120 531256
rect 62172 531247 62174 531256
rect 62120 531218 62172 531224
rect 62120 531140 62172 531146
rect 62120 531082 62172 531088
rect 62132 530641 62160 531082
rect 62118 530632 62174 530641
rect 62118 530567 62174 530576
rect 62120 528624 62172 528630
rect 62118 528592 62120 528601
rect 62172 528592 62174 528601
rect 62118 528527 62174 528536
rect 61382 527096 61438 527105
rect 61382 527031 61438 527040
rect 62960 525745 62988 552599
rect 63420 528057 63448 556679
rect 651470 553480 651526 553489
rect 651470 553415 651526 553424
rect 651484 552702 651512 553415
rect 651472 552696 651524 552702
rect 651472 552638 651524 552644
rect 651470 552392 651526 552401
rect 651470 552327 651526 552336
rect 651484 552090 651512 552327
rect 651472 552084 651524 552090
rect 651472 552026 651524 552032
rect 652022 551032 652078 551041
rect 652022 550967 652078 550976
rect 651380 550384 651432 550390
rect 651378 550352 651380 550361
rect 651432 550352 651434 550361
rect 651378 550287 651434 550296
rect 651470 549128 651526 549137
rect 651470 549063 651472 549072
rect 651524 549063 651526 549072
rect 651472 549034 651524 549040
rect 651472 548820 651524 548826
rect 651472 548762 651524 548768
rect 651484 548457 651512 548762
rect 651470 548448 651526 548457
rect 651470 548383 651526 548392
rect 63406 528048 63462 528057
rect 63406 527983 63462 527992
rect 62946 525736 63002 525745
rect 62946 525671 63002 525680
rect 652036 493338 652064 550967
rect 653416 550390 653444 565830
rect 655152 553444 655204 553450
rect 655152 553386 655204 553392
rect 653404 550384 653456 550390
rect 653404 550326 653456 550332
rect 655164 548826 655192 553386
rect 655152 548820 655204 548826
rect 655152 548762 655204 548768
rect 656176 534274 656204 594866
rect 657556 594726 657584 600442
rect 657544 594720 657596 594726
rect 657544 594662 657596 594668
rect 658936 579698 658964 642330
rect 660316 625190 660344 688638
rect 661696 670750 661724 732770
rect 668412 710054 668440 775542
rect 668768 741124 668820 741130
rect 668768 741066 668820 741072
rect 668584 733440 668636 733446
rect 668584 733382 668636 733388
rect 668400 710048 668452 710054
rect 668400 709990 668452 709996
rect 666468 697128 666520 697134
rect 666468 697070 666520 697076
rect 661684 670744 661736 670750
rect 661684 670686 661736 670692
rect 660304 625184 660356 625190
rect 660304 625126 660356 625132
rect 666480 619682 666508 697070
rect 667204 687948 667256 687954
rect 667204 687890 667256 687896
rect 667216 625870 667244 687890
rect 668398 685536 668454 685545
rect 668398 685471 668454 685480
rect 667848 661156 667900 661162
rect 667848 661098 667900 661104
rect 667388 647284 667440 647290
rect 667388 647226 667440 647232
rect 667204 625864 667256 625870
rect 667204 625806 667256 625812
rect 666468 619676 666520 619682
rect 666468 619618 666520 619624
rect 667204 596216 667256 596222
rect 667204 596158 667256 596164
rect 658924 579692 658976 579698
rect 658924 579634 658976 579640
rect 657820 554804 657872 554810
rect 657820 554746 657872 554752
rect 657832 549098 657860 554746
rect 665824 552696 665876 552702
rect 665824 552638 665876 552644
rect 660304 552084 660356 552090
rect 660304 552026 660356 552032
rect 657820 549092 657872 549098
rect 657820 549034 657872 549040
rect 656164 534268 656216 534274
rect 656164 534210 656216 534216
rect 652024 493332 652076 493338
rect 652024 493274 652076 493280
rect 660316 491366 660344 552026
rect 665836 491502 665864 552638
rect 667216 535498 667244 596158
rect 667400 571742 667428 647226
rect 667570 595504 667626 595513
rect 667570 595439 667626 595448
rect 667388 571736 667440 571742
rect 667388 571678 667440 571684
rect 667204 535492 667256 535498
rect 667204 535434 667256 535440
rect 667584 529990 667612 595439
rect 667572 529984 667624 529990
rect 667572 529926 667624 529932
rect 665824 491496 665876 491502
rect 665824 491438 665876 491444
rect 660304 491360 660356 491366
rect 660304 491302 660356 491308
rect 667860 455666 667888 661098
rect 668216 654152 668268 654158
rect 668216 654094 668268 654100
rect 668228 574462 668256 654094
rect 668412 616865 668440 685471
rect 668596 671158 668624 733382
rect 668584 671152 668636 671158
rect 668584 671094 668636 671100
rect 668780 662998 668808 741066
rect 669042 733816 669098 733825
rect 669042 733751 669098 733760
rect 668768 662992 668820 662998
rect 668768 662934 668820 662940
rect 669056 661638 669084 733751
rect 669240 710734 669268 790910
rect 670608 789404 670660 789410
rect 670608 789346 670660 789352
rect 670424 782536 670476 782542
rect 670424 782478 670476 782484
rect 670240 777028 670292 777034
rect 670240 776970 670292 776976
rect 669964 775736 670016 775742
rect 669964 775678 670016 775684
rect 669780 739968 669832 739974
rect 669780 739910 669832 739916
rect 669596 734460 669648 734466
rect 669596 734402 669648 734408
rect 669228 710728 669280 710734
rect 669228 710670 669280 710676
rect 669410 698320 669466 698329
rect 669410 698255 669466 698264
rect 669226 697368 669282 697377
rect 669226 697303 669282 697312
rect 669044 661632 669096 661638
rect 669044 661574 669096 661580
rect 669042 647864 669098 647873
rect 669042 647799 669098 647808
rect 668584 645176 668636 645182
rect 668584 645118 668636 645124
rect 668596 625598 668624 645118
rect 668858 638752 668914 638761
rect 668858 638687 668914 638696
rect 668584 625592 668636 625598
rect 668584 625534 668636 625540
rect 668398 616856 668454 616865
rect 668398 616791 668454 616800
rect 668584 597576 668636 597582
rect 668584 597518 668636 597524
rect 668216 574456 668268 574462
rect 668216 574398 668268 574404
rect 668398 555248 668454 555257
rect 668398 555183 668454 555192
rect 668412 485858 668440 555183
rect 668596 535702 668624 597518
rect 668872 574190 668900 638687
rect 668860 574184 668912 574190
rect 668860 574126 668912 574132
rect 669056 571470 669084 647799
rect 669240 619070 669268 697303
rect 669424 621246 669452 698255
rect 669608 662590 669636 734402
rect 669792 665650 669820 739910
rect 669976 715766 670004 775678
rect 669964 715760 670016 715766
rect 669964 715702 670016 715708
rect 670252 705362 670280 776970
rect 670436 710462 670464 782478
rect 670424 710456 670476 710462
rect 670424 710398 670476 710404
rect 670620 709646 670648 789346
rect 670896 713726 670924 892842
rect 671804 885692 671856 885698
rect 671804 885634 671856 885640
rect 671618 779376 671674 779385
rect 671618 779311 671674 779320
rect 671068 745272 671120 745278
rect 671068 745214 671120 745220
rect 670884 713720 670936 713726
rect 670884 713662 670936 713668
rect 670608 709640 670660 709646
rect 670608 709582 670660 709588
rect 670240 705356 670292 705362
rect 670240 705298 670292 705304
rect 670608 703860 670660 703866
rect 670608 703802 670660 703808
rect 670240 685976 670292 685982
rect 670240 685918 670292 685924
rect 669780 665644 669832 665650
rect 669780 665586 669832 665592
rect 669596 662584 669648 662590
rect 669596 662526 669648 662532
rect 669964 640348 670016 640354
rect 669964 640290 670016 640296
rect 669596 623076 669648 623082
rect 669596 623018 669648 623024
rect 669412 621240 669464 621246
rect 669412 621182 669464 621188
rect 669228 619064 669280 619070
rect 669228 619006 669280 619012
rect 669412 614916 669464 614922
rect 669412 614858 669464 614864
rect 669226 608016 669282 608025
rect 669226 607951 669282 607960
rect 669044 571464 669096 571470
rect 669044 571406 669096 571412
rect 669042 562320 669098 562329
rect 669042 562255 669098 562264
rect 668860 550656 668912 550662
rect 668860 550598 668912 550604
rect 668584 535696 668636 535702
rect 668584 535638 668636 535644
rect 668400 485852 668452 485858
rect 668400 485794 668452 485800
rect 668872 484430 668900 550598
rect 669056 484566 669084 562255
rect 669240 528630 669268 607951
rect 669228 528624 669280 528630
rect 669228 528566 669280 528572
rect 669044 484560 669096 484566
rect 669044 484502 669096 484508
rect 668860 484424 668912 484430
rect 668860 484366 668912 484372
rect 667848 455660 667900 455666
rect 667848 455602 667900 455608
rect 669424 455433 669452 614858
rect 669608 577182 669636 623018
rect 669780 622260 669832 622266
rect 669780 622202 669832 622208
rect 669792 577454 669820 622202
rect 669976 580310 670004 640290
rect 670252 619886 670280 685918
rect 670424 669384 670476 669390
rect 670424 669326 670476 669332
rect 670436 625122 670464 669326
rect 670424 625116 670476 625122
rect 670424 625058 670476 625064
rect 670240 619880 670292 619886
rect 670240 619822 670292 619828
rect 670422 600400 670478 600409
rect 670422 600335 670478 600344
rect 669964 580304 670016 580310
rect 669964 580246 670016 580252
rect 670148 578400 670200 578406
rect 670148 578342 670200 578348
rect 669964 578264 670016 578270
rect 669964 578206 670016 578212
rect 669780 577448 669832 577454
rect 669780 577390 669832 577396
rect 669596 577176 669648 577182
rect 669596 577118 669648 577124
rect 669976 534546 670004 578206
rect 670160 577130 670188 578342
rect 670068 577102 670188 577130
rect 670068 563054 670096 577102
rect 670240 577040 670292 577046
rect 670240 576982 670292 576988
rect 670252 563054 670280 576982
rect 670068 563026 670188 563054
rect 670252 563026 670372 563054
rect 669964 534540 670016 534546
rect 669964 534482 670016 534488
rect 670160 534410 670188 563026
rect 670148 534404 670200 534410
rect 670148 534346 670200 534352
rect 670344 534290 670372 563026
rect 670252 534262 670372 534290
rect 670252 533390 670280 534262
rect 670240 533384 670292 533390
rect 670240 533326 670292 533332
rect 670436 530126 670464 600335
rect 670424 530120 670476 530126
rect 670424 530062 670476 530068
rect 670620 456414 670648 703802
rect 670790 688528 670846 688537
rect 670790 688463 670846 688472
rect 670804 616622 670832 688463
rect 671080 673454 671108 745214
rect 671344 743776 671396 743782
rect 671344 743718 671396 743724
rect 671356 731338 671384 743718
rect 671344 731332 671396 731338
rect 671344 731274 671396 731280
rect 671252 730108 671304 730114
rect 671252 730050 671304 730056
rect 671264 717614 671292 730050
rect 670988 673426 671108 673454
rect 671172 717586 671292 717614
rect 670988 669254 671016 673426
rect 670976 669248 671028 669254
rect 670976 669190 671028 669196
rect 670976 666596 671028 666602
rect 670976 666538 671028 666544
rect 670988 622742 671016 666538
rect 671172 660142 671200 717586
rect 671344 713244 671396 713250
rect 671344 713186 671396 713192
rect 671356 668574 671384 713186
rect 671632 708014 671660 779311
rect 671816 728346 671844 885634
rect 671804 728340 671856 728346
rect 671804 728282 671856 728288
rect 671802 714912 671858 714921
rect 671802 714847 671858 714856
rect 672000 714854 672028 892978
rect 672356 742484 672408 742490
rect 672356 742426 672408 742432
rect 672172 735752 672224 735758
rect 672172 735694 672224 735700
rect 672184 734602 672212 735694
rect 672172 734596 672224 734602
rect 672172 734538 672224 734544
rect 671620 708008 671672 708014
rect 671620 707950 671672 707956
rect 671816 670138 671844 714847
rect 672000 714826 672212 714854
rect 671988 712428 672040 712434
rect 671988 712370 672040 712376
rect 671804 670132 671856 670138
rect 671804 670074 671856 670080
rect 671804 669248 671856 669254
rect 671804 669190 671856 669196
rect 671344 668568 671396 668574
rect 671344 668510 671396 668516
rect 671620 668228 671672 668234
rect 671620 668170 671672 668176
rect 671344 667956 671396 667962
rect 671344 667898 671396 667904
rect 671160 660136 671212 660142
rect 671160 660078 671212 660084
rect 671160 645924 671212 645930
rect 671160 645866 671212 645872
rect 671172 643657 671200 645866
rect 671158 643648 671214 643657
rect 671158 643583 671214 643592
rect 671160 624708 671212 624714
rect 671160 624650 671212 624656
rect 670976 622736 671028 622742
rect 670976 622678 671028 622684
rect 670792 616616 670844 616622
rect 670792 616558 670844 616564
rect 670974 593600 671030 593609
rect 670974 593535 671030 593544
rect 670792 534132 670844 534138
rect 670792 534074 670844 534080
rect 670804 490958 670832 534074
rect 670988 529718 671016 593535
rect 671172 580038 671200 624650
rect 671356 623558 671384 667898
rect 671632 624374 671660 668170
rect 671816 665310 671844 669190
rect 672000 666942 672028 712370
rect 672184 712201 672212 714826
rect 672170 712192 672226 712201
rect 672170 712127 672226 712136
rect 672170 690568 672226 690577
rect 672170 690503 672226 690512
rect 671988 666936 672040 666942
rect 671988 666878 672040 666884
rect 671804 665304 671856 665310
rect 671804 665246 671856 665252
rect 671986 652896 672042 652905
rect 671986 652831 672042 652840
rect 671802 641744 671858 641753
rect 671802 641679 671858 641688
rect 671620 624368 671672 624374
rect 671620 624310 671672 624316
rect 671620 623892 671672 623898
rect 671620 623834 671672 623840
rect 671344 623552 671396 623558
rect 671344 623494 671396 623500
rect 671342 594824 671398 594833
rect 671342 594759 671398 594768
rect 671160 580032 671212 580038
rect 671160 579974 671212 579980
rect 671160 576904 671212 576910
rect 671160 576846 671212 576852
rect 671172 532574 671200 576846
rect 671160 532568 671212 532574
rect 671160 532510 671212 532516
rect 670976 529712 671028 529718
rect 670976 529654 671028 529660
rect 671356 524686 671384 594759
rect 671632 578814 671660 623834
rect 671620 578808 671672 578814
rect 671620 578750 671672 578756
rect 671816 572898 671844 641679
rect 672000 575958 672028 652831
rect 672184 620634 672212 690503
rect 672368 665174 672396 742426
rect 672552 715329 672580 894406
rect 672736 866658 672764 895630
rect 675850 895520 675906 895529
rect 675850 895455 675906 895464
rect 675864 894470 675892 895455
rect 676034 894704 676090 894713
rect 676034 894639 676090 894648
rect 675852 894464 675904 894470
rect 675852 894406 675904 894412
rect 676048 894334 676076 894639
rect 673368 894328 673420 894334
rect 673368 894270 673420 894276
rect 676036 894328 676088 894334
rect 676036 894270 676088 894276
rect 673184 886916 673236 886922
rect 673184 886858 673236 886864
rect 672724 866652 672776 866658
rect 672724 866594 672776 866600
rect 673000 783896 673052 783902
rect 673000 783838 673052 783844
rect 672724 728680 672776 728686
rect 672724 728622 672776 728628
rect 672538 715320 672594 715329
rect 672538 715255 672594 715264
rect 672538 694648 672594 694657
rect 672538 694583 672594 694592
rect 672356 665168 672408 665174
rect 672356 665110 672408 665116
rect 672172 620628 672224 620634
rect 672172 620570 672224 620576
rect 672552 619041 672580 694583
rect 672736 663921 672764 728622
rect 673012 717614 673040 783838
rect 673196 728142 673224 886858
rect 673184 728136 673236 728142
rect 673184 728078 673236 728084
rect 673380 717614 673408 894270
rect 675850 893888 675906 893897
rect 675850 893823 675906 893832
rect 675864 892906 675892 893823
rect 676034 893072 676090 893081
rect 676034 893007 676036 893016
rect 676088 893007 676090 893016
rect 676036 892978 676088 892984
rect 675852 892900 675904 892906
rect 675852 892842 675904 892848
rect 676034 892664 676090 892673
rect 676090 892622 676444 892650
rect 676034 892599 676090 892608
rect 676034 891440 676090 891449
rect 676034 891375 676090 891384
rect 675206 891032 675262 891041
rect 675206 890967 675262 890976
rect 674932 890384 674984 890390
rect 674932 890326 674984 890332
rect 674472 888956 674524 888962
rect 674472 888898 674524 888904
rect 674288 887324 674340 887330
rect 674288 887266 674340 887272
rect 674300 868601 674328 887266
rect 674484 869666 674512 888898
rect 674746 888584 674802 888593
rect 674746 888519 674802 888528
rect 674760 881834 674788 888519
rect 674668 881806 674788 881834
rect 674668 870890 674696 881806
rect 674794 878688 674846 878694
rect 674846 878636 674880 878642
rect 674794 878630 674880 878636
rect 674806 878614 674880 878630
rect 674852 877690 674880 878614
rect 674806 877662 674880 877690
rect 674806 877554 674834 877662
rect 674806 877526 674880 877554
rect 674852 877418 674880 877526
rect 674760 877390 674880 877418
rect 674760 876602 674788 877390
rect 674760 876574 674834 876602
rect 674806 876466 674834 876574
rect 674806 876438 674880 876466
rect 674852 873730 674880 876438
rect 674944 874290 674972 890326
rect 675220 887354 675248 890967
rect 676048 890390 676076 891375
rect 676036 890384 676088 890390
rect 676036 890326 676088 890332
rect 676034 890216 676090 890225
rect 676090 890186 676260 890202
rect 676090 890180 676272 890186
rect 676090 890174 676220 890180
rect 676034 890151 676090 890160
rect 676220 890122 676272 890128
rect 676034 889400 676090 889409
rect 676090 889358 676260 889386
rect 676034 889335 676090 889344
rect 676034 888992 676090 889001
rect 676034 888927 676036 888936
rect 676088 888927 676090 888936
rect 676036 888898 676088 888904
rect 676232 888758 676260 889358
rect 676220 888752 676272 888758
rect 676220 888694 676272 888700
rect 675128 887326 675248 887354
rect 676034 887360 676090 887369
rect 675128 879458 675156 887326
rect 676034 887295 676036 887304
rect 676088 887295 676090 887304
rect 676036 887266 676088 887272
rect 676034 886952 676090 886961
rect 676034 886887 676036 886896
rect 676088 886887 676090 886896
rect 676036 886858 676088 886864
rect 676034 885728 676090 885737
rect 676034 885663 676036 885672
rect 676088 885663 676090 885672
rect 676036 885634 676088 885640
rect 675576 880524 675628 880530
rect 675576 880466 675628 880472
rect 675036 879430 675156 879458
rect 675036 874562 675064 879430
rect 675392 879368 675444 879374
rect 675392 879310 675444 879316
rect 675208 879096 675260 879102
rect 675208 879038 675260 879044
rect 675220 877010 675248 879038
rect 675404 878642 675432 879310
rect 675312 878614 675432 878642
rect 675312 877146 675340 878614
rect 675588 878084 675616 880466
rect 675944 880456 675996 880462
rect 675944 880398 675996 880404
rect 675760 879232 675812 879238
rect 675760 879174 675812 879180
rect 675772 878529 675800 879174
rect 675758 878520 675814 878529
rect 675956 878490 675984 880398
rect 676416 879102 676444 892622
rect 679622 891848 679678 891857
rect 679622 891783 679678 891792
rect 676864 890180 676916 890186
rect 676864 890122 676916 890128
rect 676876 879374 676904 890122
rect 678242 889808 678298 889817
rect 678242 889743 678298 889752
rect 677048 888752 677100 888758
rect 677048 888694 677100 888700
rect 676864 879368 676916 879374
rect 676864 879310 676916 879316
rect 676404 879096 676456 879102
rect 676404 879038 676456 879044
rect 677060 878694 677088 888694
rect 678256 879238 678284 889743
rect 679636 880462 679664 891783
rect 681002 890624 681058 890633
rect 681002 890559 681058 890568
rect 681016 880705 681044 890559
rect 683118 888176 683174 888185
rect 683118 888111 683174 888120
rect 681002 880696 681058 880705
rect 681002 880631 681058 880640
rect 679624 880456 679676 880462
rect 683132 880433 683160 888111
rect 679624 880398 679676 880404
rect 683118 880424 683174 880433
rect 683118 880359 683174 880368
rect 678244 879232 678296 879238
rect 678244 879174 678296 879180
rect 677048 878688 677100 878694
rect 677048 878630 677100 878636
rect 675758 878455 675814 878464
rect 675944 878484 675996 878490
rect 675944 878426 675996 878432
rect 675484 877804 675536 877810
rect 675484 877746 675536 877752
rect 675496 877540 675524 877746
rect 675312 877118 675432 877146
rect 675220 876982 675340 877010
rect 675312 876262 675340 876982
rect 675404 876860 675432 877118
rect 675312 876234 675418 876262
rect 675036 874534 675248 874562
rect 675220 874342 675248 874534
rect 675208 874336 675260 874342
rect 674944 874262 675064 874290
rect 675208 874278 675260 874284
rect 675036 874070 675064 874262
rect 675208 874200 675260 874206
rect 675208 874142 675260 874148
rect 675024 874064 675076 874070
rect 675024 874006 675076 874012
rect 674840 873724 674892 873730
rect 674840 873666 674892 873672
rect 675220 873610 675248 874142
rect 675404 874070 675432 874412
rect 675574 874168 675630 874177
rect 675574 874103 675630 874112
rect 675392 874064 675444 874070
rect 675392 874006 675444 874012
rect 675588 873868 675616 874103
rect 675392 873724 675444 873730
rect 675392 873666 675444 873672
rect 675220 873582 675340 873610
rect 675022 873080 675078 873089
rect 675022 873015 675078 873024
rect 674668 870862 674880 870890
rect 674484 869638 674696 869666
rect 674668 869122 674696 869638
rect 674852 869310 674880 870862
rect 675036 869530 675064 873015
rect 675312 870074 675340 873582
rect 675404 873188 675432 873666
rect 675758 872808 675814 872817
rect 675758 872743 675814 872752
rect 675772 872576 675800 872743
rect 675312 870046 675418 870074
rect 675036 869502 675418 869530
rect 675024 869440 675076 869446
rect 675022 869408 675024 869417
rect 675076 869408 675078 869417
rect 675022 869343 675078 869352
rect 674840 869304 674892 869310
rect 674840 869246 674892 869252
rect 675300 869304 675352 869310
rect 675300 869246 675352 869252
rect 674668 869094 674880 869122
rect 674286 868592 674342 868601
rect 674286 868527 674342 868536
rect 674852 867610 674880 869094
rect 675022 869000 675078 869009
rect 675022 868935 675078 868944
rect 675036 868578 675064 868935
rect 675312 868889 675340 869246
rect 675312 868861 675418 868889
rect 675390 868592 675446 868601
rect 675036 868550 675248 868578
rect 675024 868080 675076 868086
rect 675024 868022 675076 868028
rect 674840 867604 674892 867610
rect 674840 867546 674892 867552
rect 675036 865858 675064 868022
rect 675220 867694 675248 868550
rect 675390 868527 675446 868536
rect 675404 868224 675432 868527
rect 675220 867666 675418 867694
rect 675208 867604 675260 867610
rect 675208 867546 675260 867552
rect 675220 867049 675248 867546
rect 675220 867021 675418 867049
rect 675036 865830 675418 865858
rect 675298 865736 675354 865745
rect 675298 865671 675354 865680
rect 675312 863818 675340 865671
rect 675758 865464 675814 865473
rect 675758 865399 675814 865408
rect 675772 865195 675800 865399
rect 675666 865056 675722 865065
rect 675666 864991 675722 865000
rect 675680 864552 675708 864991
rect 675312 863790 675432 863818
rect 675404 863328 675432 863790
rect 675208 790968 675260 790974
rect 675208 790910 675260 790916
rect 675220 790650 675248 790910
rect 675392 790832 675444 790838
rect 675392 790774 675444 790780
rect 675220 790622 675340 790650
rect 675116 789404 675168 789410
rect 675116 789346 675168 789352
rect 675128 787693 675156 789346
rect 675312 788338 675340 790622
rect 675404 788868 675432 790774
rect 675312 788310 675418 788338
rect 675128 787665 675418 787693
rect 675772 786729 675800 787032
rect 675758 786720 675814 786729
rect 675758 786655 675814 786664
rect 674852 785182 675418 785210
rect 673552 780020 673604 780026
rect 673552 779962 673604 779968
rect 673564 717614 673592 779962
rect 673734 778832 673790 778841
rect 673734 778767 673790 778776
rect 673748 760394 673776 778767
rect 674470 777472 674526 777481
rect 674470 777407 674526 777416
rect 674102 775704 674158 775713
rect 674102 775639 674158 775648
rect 672920 717586 673040 717614
rect 673104 717586 673408 717614
rect 673472 717586 673592 717614
rect 673656 760366 673776 760394
rect 672920 709209 672948 717586
rect 673104 714513 673132 717586
rect 673276 715760 673328 715766
rect 673274 715728 673276 715737
rect 673328 715728 673330 715737
rect 673274 715663 673330 715672
rect 673090 714504 673146 714513
rect 673090 714439 673146 714448
rect 673274 714096 673330 714105
rect 673274 714031 673330 714040
rect 672906 709200 672962 709209
rect 672906 709135 672962 709144
rect 673288 707954 673316 714031
rect 673472 713017 673500 717586
rect 673458 713008 673514 713017
rect 673458 712943 673514 712952
rect 673656 712858 673684 760366
rect 674116 746594 674144 775639
rect 674484 746594 674512 777407
rect 674852 770054 674880 785182
rect 675128 784638 675418 784666
rect 675128 783902 675156 784638
rect 675116 783896 675168 783902
rect 675496 783873 675524 783972
rect 675116 783838 675168 783844
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675128 783346 675418 783374
rect 675128 782513 675156 783346
rect 675300 782536 675352 782542
rect 675114 782504 675170 782513
rect 675300 782478 675352 782484
rect 675114 782439 675170 782448
rect 675312 781402 675340 782478
rect 675312 781374 675432 781402
rect 675024 781108 675076 781114
rect 675024 781050 675076 781056
rect 675036 780994 675064 781050
rect 674944 780966 675064 780994
rect 674944 779714 674972 780966
rect 675404 780844 675432 781374
rect 675312 780422 675432 780450
rect 675312 780314 675340 780422
rect 675128 780286 675340 780314
rect 675404 780300 675432 780422
rect 675128 780026 675156 780286
rect 675116 780020 675168 780026
rect 675116 779962 675168 779968
rect 674944 779686 675340 779714
rect 675024 778524 675076 778530
rect 675024 778466 675076 778472
rect 675312 778478 675340 779686
rect 675496 779385 675524 779688
rect 675482 779376 675538 779385
rect 675482 779311 675538 779320
rect 675496 778841 675524 779008
rect 675482 778832 675538 778841
rect 675482 778767 675538 778776
rect 675036 778274 675064 778466
rect 675312 778450 675418 778478
rect 675036 778246 675340 778274
rect 675312 777050 675340 778246
rect 675496 777481 675524 777852
rect 675482 777472 675538 777481
rect 675482 777407 675538 777416
rect 675024 777028 675076 777034
rect 675312 777022 675432 777050
rect 675024 776970 675076 776976
rect 675036 776914 675064 776970
rect 675036 776886 675340 776914
rect 675024 775600 675076 775606
rect 675024 775542 675076 775548
rect 675036 774194 675064 775542
rect 675312 775350 675340 776886
rect 675404 776628 675432 777022
rect 675496 775713 675524 776016
rect 675482 775704 675538 775713
rect 675482 775639 675538 775648
rect 675312 775322 675418 775350
rect 675036 774166 675340 774194
rect 675312 774058 675340 774166
rect 675404 774058 675432 774180
rect 675312 774030 675432 774058
rect 674852 770026 675248 770054
rect 675220 746594 675248 770026
rect 674116 746566 674328 746594
rect 674484 746566 674696 746594
rect 673826 735720 673882 735729
rect 673826 735655 673882 735664
rect 673840 727410 673868 735655
rect 674102 735040 674158 735049
rect 674102 734975 674158 734984
rect 674116 727954 674144 734975
rect 674300 728113 674328 746566
rect 674472 731876 674524 731882
rect 674472 731818 674524 731824
rect 674286 728104 674342 728113
rect 674286 728039 674342 728048
rect 674116 727926 674236 727954
rect 673564 712830 673684 712858
rect 673748 727382 673868 727410
rect 673564 712745 673592 712830
rect 673550 712736 673606 712745
rect 673550 712671 673606 712680
rect 673288 707926 673408 707954
rect 672998 695600 673054 695609
rect 672998 695535 673054 695544
rect 672722 663912 672778 663921
rect 672722 663847 672778 663856
rect 672722 651400 672778 651409
rect 672722 651335 672778 651344
rect 672538 619032 672594 619041
rect 672538 618967 672594 618976
rect 672538 606520 672594 606529
rect 672538 606455 672594 606464
rect 672262 603528 672318 603537
rect 672262 603463 672318 603472
rect 671988 575952 672040 575958
rect 671988 575894 672040 575900
rect 671804 572892 671856 572898
rect 671804 572834 671856 572840
rect 671986 553480 672042 553489
rect 671986 553415 672042 553424
rect 671620 533588 671672 533594
rect 671620 533530 671672 533536
rect 671344 524680 671396 524686
rect 671344 524622 671396 524628
rect 670792 490952 670844 490958
rect 670792 490894 670844 490900
rect 671632 490142 671660 533530
rect 671804 532772 671856 532778
rect 671804 532714 671856 532720
rect 671620 490136 671672 490142
rect 671620 490078 671672 490084
rect 671816 489326 671844 532714
rect 671804 489320 671856 489326
rect 671804 489262 671856 489268
rect 672000 482390 672028 553415
rect 672276 528494 672304 603463
rect 672552 538214 672580 606455
rect 672736 576473 672764 651335
rect 673012 621014 673040 695535
rect 673184 685976 673236 685982
rect 673184 685918 673236 685924
rect 673196 685817 673224 685918
rect 673182 685808 673238 685817
rect 673182 685743 673238 685752
rect 673380 669497 673408 707926
rect 673552 701072 673604 701078
rect 673550 701040 673552 701049
rect 673604 701040 673606 701049
rect 673550 700975 673606 700984
rect 673552 697128 673604 697134
rect 673550 697096 673552 697105
rect 673604 697096 673606 697105
rect 673550 697031 673606 697040
rect 673552 690056 673604 690062
rect 673550 690024 673552 690033
rect 673604 690024 673606 690033
rect 673550 689959 673606 689968
rect 673552 688832 673604 688838
rect 673552 688774 673604 688780
rect 673564 687721 673592 688774
rect 673550 687712 673606 687721
rect 673550 687647 673606 687656
rect 673748 683114 673776 727382
rect 673918 727288 673974 727297
rect 673918 727223 673974 727232
rect 673932 717614 673960 727223
rect 674208 724514 674236 727926
rect 674484 727297 674512 731818
rect 674668 727841 674696 746566
rect 674852 746566 675248 746594
rect 674852 731134 674880 746566
rect 675116 745272 675168 745278
rect 675116 745214 675168 745220
rect 675128 743322 675156 745214
rect 675496 743782 675524 743852
rect 675484 743776 675536 743782
rect 675484 743718 675536 743724
rect 675128 743294 675418 743322
rect 675404 742490 675432 742696
rect 675392 742484 675444 742490
rect 675392 742426 675444 742432
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 674944 742002 675340 742030
rect 675404 742016 675432 742070
rect 674944 732034 674972 742002
rect 675300 741124 675352 741130
rect 675300 741066 675352 741072
rect 675312 741010 675340 741066
rect 675220 740982 675340 741010
rect 675220 739038 675248 740982
rect 675404 739974 675432 740180
rect 675392 739968 675444 739974
rect 675392 739910 675444 739916
rect 675758 739800 675814 739809
rect 675758 739735 675814 739744
rect 675772 739636 675800 739735
rect 675220 739010 675340 739038
rect 675312 738970 675340 739010
rect 675404 738970 675432 739024
rect 675312 738942 675432 738970
rect 675312 738330 675418 738358
rect 675312 738177 675340 738330
rect 675298 738168 675354 738177
rect 675298 738103 675354 738112
rect 675496 735729 675524 735896
rect 675482 735720 675538 735729
rect 675482 735655 675538 735664
rect 675496 735049 675524 735319
rect 675482 735040 675538 735049
rect 675482 734975 675538 734984
rect 675128 734658 675418 734686
rect 675128 734466 675156 734658
rect 675300 734596 675352 734602
rect 675300 734538 675352 734544
rect 675116 734460 675168 734466
rect 675116 734402 675168 734408
rect 675116 734324 675168 734330
rect 675116 734266 675168 734272
rect 674944 732006 675064 732034
rect 674840 731128 674892 731134
rect 674840 731070 674892 731076
rect 674840 730516 674892 730522
rect 674840 730458 674892 730464
rect 674654 727832 674710 727841
rect 674654 727767 674710 727776
rect 674470 727288 674526 727297
rect 674470 727223 674526 727232
rect 674208 724486 674420 724514
rect 674392 721750 674420 724486
rect 674852 722265 674880 730458
rect 674838 722256 674894 722265
rect 674838 722191 674894 722200
rect 674654 721984 674710 721993
rect 675036 721970 675064 732006
rect 675128 731626 675156 734266
rect 675312 734174 675340 734538
rect 675220 734146 675340 734174
rect 675220 733493 675248 734146
rect 675588 733825 675616 734031
rect 675574 733816 675630 733825
rect 675574 733751 675630 733760
rect 675220 733465 675418 733493
rect 675312 732822 675418 732850
rect 675312 731882 675340 732822
rect 675300 731876 675352 731882
rect 675300 731818 675352 731824
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 675128 731598 675340 731626
rect 675404 731612 675432 731734
rect 675208 730924 675260 730930
rect 675208 730866 675260 730872
rect 675220 730810 675248 730866
rect 674710 721942 675064 721970
rect 675128 730782 675248 730810
rect 674654 721919 674710 721928
rect 675128 721750 675156 730782
rect 675404 730674 675432 731000
rect 675312 730646 675432 730674
rect 675312 730522 675340 730646
rect 675300 730516 675352 730522
rect 675300 730458 675352 730464
rect 675312 730337 675418 730365
rect 675312 730114 675340 730337
rect 675300 730108 675352 730114
rect 675300 730050 675352 730056
rect 675312 729150 675418 729178
rect 675312 728686 675340 729150
rect 675300 728680 675352 728686
rect 675300 728622 675352 728628
rect 675850 728104 675906 728113
rect 675850 728039 675906 728048
rect 675864 727938 675892 728039
rect 675852 727932 675904 727938
rect 675852 727874 675904 727880
rect 683304 727932 683356 727938
rect 683304 727874 683356 727880
rect 676034 727832 676090 727841
rect 676034 727767 676090 727776
rect 676048 726578 676076 727767
rect 681002 726880 681058 726889
rect 681002 726815 681058 726824
rect 676036 726572 676088 726578
rect 676036 726514 676088 726520
rect 674380 721744 674432 721750
rect 674380 721686 674432 721692
rect 675116 721744 675168 721750
rect 675116 721686 675168 721692
rect 674380 721268 674432 721274
rect 674380 721210 674432 721216
rect 675116 721268 675168 721274
rect 675116 721210 675168 721216
rect 674392 720866 674420 721210
rect 675128 720866 675156 721210
rect 674380 720860 674432 720866
rect 674380 720802 674432 720808
rect 675116 720860 675168 720866
rect 675116 720802 675168 720808
rect 674380 720520 674432 720526
rect 674380 720462 674432 720468
rect 675392 720520 675444 720526
rect 675392 720462 675444 720468
rect 673656 683086 673776 683114
rect 673840 717586 673960 717614
rect 673656 682553 673684 683086
rect 673642 682544 673698 682553
rect 673642 682479 673698 682488
rect 673840 682394 673868 717586
rect 674010 716544 674066 716553
rect 674010 716479 674066 716488
rect 674024 716310 674052 716479
rect 674012 716304 674064 716310
rect 674012 716246 674064 716252
rect 674010 716136 674066 716145
rect 674010 716071 674066 716080
rect 674024 714950 674052 716071
rect 674012 714944 674064 714950
rect 674012 714886 674064 714892
rect 674392 714854 674420 720462
rect 674208 714826 674420 714854
rect 674012 713720 674064 713726
rect 674010 713688 674012 713697
rect 674064 713688 674066 713697
rect 674010 713623 674066 713632
rect 674010 713280 674066 713289
rect 674010 713215 674012 713224
rect 674064 713215 674066 713224
rect 674012 713186 674064 713192
rect 674010 712464 674066 712473
rect 674010 712399 674012 712408
rect 674064 712399 674066 712408
rect 674012 712370 674064 712376
rect 674010 711240 674066 711249
rect 674010 711175 674066 711184
rect 674024 710734 674052 711175
rect 674012 710728 674064 710734
rect 674012 710670 674064 710676
rect 674012 710456 674064 710462
rect 674010 710424 674012 710433
rect 674064 710424 674066 710433
rect 674010 710359 674066 710368
rect 674012 710048 674064 710054
rect 674010 710016 674012 710025
rect 674064 710016 674066 710025
rect 674010 709951 674066 709960
rect 674012 709640 674064 709646
rect 674010 709608 674012 709617
rect 674064 709608 674066 709617
rect 674010 709543 674066 709552
rect 674012 708008 674064 708014
rect 674010 707976 674012 707985
rect 674064 707976 674066 707985
rect 674010 707911 674066 707920
rect 674010 705392 674066 705401
rect 674010 705327 674012 705336
rect 674064 705327 674066 705336
rect 674012 705298 674064 705304
rect 674010 705120 674066 705129
rect 674010 705055 674066 705064
rect 674024 703866 674052 705055
rect 674012 703860 674064 703866
rect 674012 703802 674064 703808
rect 674208 702434 674236 714826
rect 674746 713008 674802 713017
rect 674746 712943 674802 712952
rect 674378 712736 674434 712745
rect 674378 712671 674434 712680
rect 674392 706761 674420 712671
rect 674760 707169 674788 712943
rect 674930 712872 674986 712881
rect 674930 712807 674986 712816
rect 674944 712201 674972 712807
rect 674930 712192 674986 712201
rect 674930 712127 674986 712136
rect 675404 710841 675432 720462
rect 681016 712065 681044 726815
rect 683118 726472 683174 726481
rect 683118 726407 683174 726416
rect 681002 712056 681058 712065
rect 681002 711991 681058 712000
rect 675390 710832 675446 710841
rect 675390 710767 675446 710776
rect 683132 708801 683160 726407
rect 683316 711657 683344 727874
rect 683488 726572 683540 726578
rect 683488 726514 683540 726520
rect 683302 711648 683358 711657
rect 683302 711583 683358 711592
rect 683118 708792 683174 708801
rect 683118 708727 683174 708736
rect 683500 708393 683528 726514
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683486 708384 683542 708393
rect 683486 708319 683542 708328
rect 674746 707160 674802 707169
rect 674746 707095 674802 707104
rect 674378 706752 674434 706761
rect 674378 706687 674434 706696
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 675850 705392 675906 705401
rect 675850 705327 675906 705336
rect 675864 705226 675892 705327
rect 683132 705226 683160 705463
rect 675852 705220 675904 705226
rect 675852 705162 675904 705168
rect 683120 705220 683172 705226
rect 683120 705162 683172 705168
rect 673656 682366 673868 682394
rect 673932 702406 674236 702434
rect 673656 682281 673684 682366
rect 673642 682272 673698 682281
rect 673642 682207 673698 682216
rect 673932 673454 673960 702406
rect 675114 701040 675170 701049
rect 675114 700975 675170 700984
rect 675128 698889 675156 700975
rect 675128 698861 675418 698889
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 675128 697666 675418 697694
rect 675128 697377 675156 697666
rect 675114 697368 675170 697377
rect 675114 697303 675170 697312
rect 675114 697096 675170 697105
rect 675114 697031 675170 697040
rect 674930 695600 674986 695609
rect 674930 695535 674986 695544
rect 674944 694022 674972 695535
rect 675128 695209 675156 697031
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695181 675418 695209
rect 675312 694742 675432 694770
rect 675114 694648 675170 694657
rect 675312 694634 675340 694742
rect 675170 694606 675340 694634
rect 675404 694620 675432 694742
rect 675114 694583 675170 694592
rect 674944 693994 675418 694022
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 674760 693314 675340 693342
rect 675404 693328 675432 693382
rect 674288 690056 674340 690062
rect 674288 689998 674340 690004
rect 674102 689208 674158 689217
rect 674102 689143 674158 689152
rect 674116 683114 674144 689143
rect 674300 683114 674328 689998
rect 674472 687268 674524 687274
rect 674472 687210 674524 687216
rect 674116 683086 674236 683114
rect 674300 683086 674420 683114
rect 673840 673426 673960 673454
rect 673642 671392 673698 671401
rect 673642 671327 673698 671336
rect 673656 670750 673684 671327
rect 673644 670744 673696 670750
rect 673644 670686 673696 670692
rect 673642 670576 673698 670585
rect 673642 670511 673698 670520
rect 673656 669526 673684 670511
rect 673644 669520 673696 669526
rect 673366 669488 673422 669497
rect 673644 669462 673696 669468
rect 673366 669423 673422 669432
rect 673642 668944 673698 668953
rect 673642 668879 673698 668888
rect 673656 668234 673684 668879
rect 673644 668228 673696 668234
rect 673644 668170 673696 668176
rect 673642 667312 673698 667321
rect 673642 667247 673698 667256
rect 673656 666602 673684 667247
rect 673644 666596 673696 666602
rect 673644 666538 673696 666544
rect 673642 666088 673698 666097
rect 673642 666023 673698 666032
rect 673656 665310 673684 666023
rect 673644 665304 673696 665310
rect 673644 665246 673696 665252
rect 673368 665168 673420 665174
rect 673368 665110 673420 665116
rect 673380 664193 673408 665110
rect 673642 664864 673698 664873
rect 673642 664799 673698 664808
rect 673366 664184 673422 664193
rect 673366 664119 673422 664128
rect 673656 663921 673684 664799
rect 673642 663912 673698 663921
rect 673642 663847 673698 663856
rect 673840 662017 673868 673426
rect 674012 671152 674064 671158
rect 674012 671094 674064 671100
rect 674024 670993 674052 671094
rect 674010 670984 674066 670993
rect 674010 670919 674066 670928
rect 674010 670168 674066 670177
rect 674010 670103 674012 670112
rect 674064 670103 674066 670112
rect 674012 670074 674064 670080
rect 674010 669760 674066 669769
rect 674010 669695 674066 669704
rect 674024 669390 674052 669695
rect 674012 669384 674064 669390
rect 674012 669326 674064 669332
rect 674012 668568 674064 668574
rect 674010 668536 674012 668545
rect 674064 668536 674066 668545
rect 674010 668471 674066 668480
rect 674010 668128 674066 668137
rect 674010 668063 674066 668072
rect 674024 667962 674052 668063
rect 674012 667956 674064 667962
rect 674012 667898 674064 667904
rect 674010 667720 674066 667729
rect 674010 667655 674066 667664
rect 674024 666942 674052 667655
rect 674012 666936 674064 666942
rect 674012 666878 674064 666884
rect 674010 665680 674066 665689
rect 674010 665615 674012 665624
rect 674064 665615 674066 665624
rect 674012 665586 674064 665592
rect 674010 663640 674066 663649
rect 674010 663575 674066 663584
rect 674024 662998 674052 663575
rect 674012 662992 674064 662998
rect 674012 662934 674064 662940
rect 674010 662824 674066 662833
rect 674010 662759 674066 662768
rect 674024 662590 674052 662759
rect 674012 662584 674064 662590
rect 674012 662526 674064 662532
rect 673826 662008 673882 662017
rect 673826 661943 673882 661952
rect 674012 661632 674064 661638
rect 674010 661600 674012 661609
rect 674064 661600 674066 661609
rect 674010 661535 674066 661544
rect 674010 661192 674066 661201
rect 674010 661127 674012 661136
rect 674064 661127 674066 661136
rect 674012 661098 674064 661104
rect 674012 660136 674064 660142
rect 674010 660104 674012 660113
rect 674064 660104 674066 660113
rect 674010 660039 674066 660048
rect 673274 659696 673330 659705
rect 673274 659631 673330 659640
rect 672920 620986 673040 621014
rect 672920 618633 672948 620986
rect 673092 620628 673144 620634
rect 673092 620570 673144 620576
rect 673104 620265 673132 620570
rect 673090 620256 673146 620265
rect 673090 620191 673146 620200
rect 673092 619880 673144 619886
rect 673090 619848 673092 619857
rect 673144 619848 673146 619857
rect 673090 619783 673146 619792
rect 672906 618624 672962 618633
rect 672906 618559 672962 618568
rect 673090 604344 673146 604353
rect 673090 604279 673146 604288
rect 672906 599720 672962 599729
rect 672906 599655 672962 599664
rect 672722 576464 672778 576473
rect 672722 576399 672778 576408
rect 672724 557864 672776 557870
rect 672724 557806 672776 557812
rect 672736 555490 672764 557806
rect 672724 555484 672776 555490
rect 672724 555426 672776 555432
rect 672920 549254 672948 599655
rect 673104 596174 673132 604279
rect 673104 596146 673224 596174
rect 673196 567194 673224 596146
rect 672828 549226 672948 549254
rect 673012 567166 673224 567194
rect 672828 539594 672856 549226
rect 673012 548842 673040 567166
rect 673288 557870 673316 659631
rect 674010 655616 674066 655625
rect 674010 655551 674012 655560
rect 674064 655551 674066 655560
rect 674012 655522 674064 655528
rect 674012 654152 674064 654158
rect 674010 654120 674012 654129
rect 674064 654120 674066 654129
rect 674010 654055 674066 654064
rect 673642 649224 673698 649233
rect 673642 649159 673698 649168
rect 673458 625968 673514 625977
rect 673458 625903 673514 625912
rect 673472 625258 673500 625903
rect 673460 625252 673512 625258
rect 673460 625194 673512 625200
rect 673458 620664 673514 620673
rect 673458 620599 673514 620608
rect 673472 619682 673500 620599
rect 673460 619676 673512 619682
rect 673460 619618 673512 619624
rect 673458 619440 673514 619449
rect 673458 619375 673514 619384
rect 673472 619070 673500 619375
rect 673460 619064 673512 619070
rect 673460 619006 673512 619012
rect 673460 616616 673512 616622
rect 673458 616584 673460 616593
rect 673512 616584 673514 616593
rect 673458 616519 673514 616528
rect 673458 614952 673514 614961
rect 673458 614887 673460 614896
rect 673512 614887 673514 614896
rect 673460 614858 673512 614864
rect 673458 611416 673514 611425
rect 673458 611351 673460 611360
rect 673512 611351 673514 611360
rect 673460 611322 673512 611328
rect 673460 600500 673512 600506
rect 673460 600442 673512 600448
rect 673472 600137 673500 600442
rect 673458 600128 673514 600137
rect 673458 600063 673514 600072
rect 673458 599040 673514 599049
rect 673458 598975 673460 598984
rect 673512 598975 673514 598984
rect 673460 598946 673512 598952
rect 673656 596174 673684 649159
rect 674010 647320 674066 647329
rect 674010 647255 674012 647264
rect 674064 647255 674066 647264
rect 674012 647226 674064 647232
rect 674208 647234 674236 683086
rect 674208 647206 674328 647234
rect 673826 644736 673882 644745
rect 673826 644671 673882 644680
rect 673840 640334 673868 644671
rect 674012 643136 674064 643142
rect 674010 643104 674012 643113
rect 674064 643104 674066 643113
rect 674010 643039 674066 643048
rect 674300 642649 674328 647206
rect 674392 643838 674420 683086
rect 674484 649994 674512 687210
rect 674760 683114 674788 693314
rect 675128 690866 675418 690894
rect 675128 690577 675156 690866
rect 675114 690568 675170 690577
rect 675114 690503 675170 690512
rect 675128 690322 675340 690350
rect 675128 690062 675156 690322
rect 675312 690282 675340 690322
rect 675404 690282 675432 690336
rect 675312 690254 675432 690282
rect 675116 690056 675168 690062
rect 674930 690024 674986 690033
rect 675116 689998 675168 690004
rect 674930 689959 674986 689968
rect 674944 688378 674972 689959
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 675128 689642 675340 689670
rect 675404 689656 675432 689710
rect 675128 689217 675156 689642
rect 675114 689208 675170 689217
rect 675114 689143 675170 689152
rect 675128 689030 675418 689058
rect 675128 688537 675156 689030
rect 675114 688528 675170 688537
rect 675114 688463 675170 688472
rect 675404 688378 675432 688500
rect 674944 688350 675432 688378
rect 675128 687806 675418 687834
rect 675128 687274 675156 687806
rect 675298 687712 675354 687721
rect 675298 687647 675354 687656
rect 675116 687268 675168 687274
rect 675116 687210 675168 687216
rect 674930 687168 674986 687177
rect 674930 687103 674986 687112
rect 674668 683086 674788 683114
rect 674944 683114 674972 687103
rect 675312 686610 675340 687647
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675758 686216 675814 686225
rect 675758 686151 675814 686160
rect 675772 685984 675800 686151
rect 675114 685808 675170 685817
rect 675114 685743 675170 685752
rect 675128 685658 675156 685743
rect 675036 685630 675156 685658
rect 675036 684162 675064 685630
rect 675482 685536 675538 685545
rect 675482 685471 675538 685480
rect 675496 685372 675524 685471
rect 675036 684134 675418 684162
rect 674944 683086 675340 683114
rect 674668 649994 674696 683086
rect 675312 676433 675340 683086
rect 675852 682576 675904 682582
rect 675850 682544 675852 682553
rect 683212 682576 683264 682582
rect 675904 682544 675906 682553
rect 683212 682518 683264 682524
rect 675850 682479 675906 682488
rect 675852 682304 675904 682310
rect 675666 682272 675722 682281
rect 675722 682252 675852 682258
rect 675722 682246 675904 682252
rect 675722 682230 675892 682246
rect 675666 682207 675722 682216
rect 682382 682136 682438 682145
rect 682382 682071 682438 682080
rect 678242 681864 678298 681873
rect 678242 681799 678298 681808
rect 675298 676424 675354 676433
rect 675298 676359 675354 676368
rect 678256 667049 678284 681799
rect 678242 667040 678298 667049
rect 678242 666975 678298 666984
rect 682396 666641 682424 682071
rect 682382 666632 682438 666641
rect 682382 666567 682438 666576
rect 683224 665417 683252 682518
rect 683396 682440 683448 682446
rect 683396 682382 683448 682388
rect 683210 665408 683266 665417
rect 683210 665343 683266 665352
rect 683408 663377 683436 682382
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683394 663368 683450 663377
rect 683394 663303 683450 663312
rect 675850 660104 675906 660113
rect 675850 660039 675906 660048
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 675864 659870 675892 660039
rect 683132 659870 683160 660039
rect 675852 659864 675904 659870
rect 675852 659806 675904 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675114 655616 675170 655625
rect 675114 655551 675170 655560
rect 674930 654120 674986 654129
rect 674930 654055 674986 654064
rect 674944 652474 674972 654055
rect 675128 653698 675156 655551
rect 675128 653670 675418 653698
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675312 652582 675432 652610
rect 675312 652474 675340 652582
rect 674944 652446 675340 652474
rect 675404 652460 675432 652582
rect 675128 651834 675418 651862
rect 675128 651409 675156 651834
rect 675114 651400 675170 651409
rect 675114 651335 675170 651344
rect 674484 649966 674604 649994
rect 674668 649966 674788 649994
rect 674576 644065 674604 649966
rect 674562 644056 674618 644065
rect 674562 643991 674618 644000
rect 674392 643810 674512 643838
rect 674484 643770 674512 643810
rect 674484 643742 674604 643770
rect 674576 643686 674604 643742
rect 674564 643680 674616 643686
rect 674564 643622 674616 643628
rect 674564 643340 674616 643346
rect 674616 643288 674696 643294
rect 674564 643282 674696 643288
rect 674576 643266 674696 643282
rect 674472 643136 674524 643142
rect 674472 643078 674524 643084
rect 674116 642621 674328 642649
rect 673840 640306 673960 640334
rect 673932 630674 673960 640306
rect 674116 636857 674144 642621
rect 674484 642546 674512 643078
rect 674300 642518 674512 642546
rect 674102 636848 674158 636857
rect 674102 636783 674158 636792
rect 673472 596146 673684 596174
rect 673748 630646 673960 630674
rect 673472 591297 673500 596146
rect 673748 592034 673776 630646
rect 674010 626376 674066 626385
rect 674010 626311 674066 626320
rect 674024 625870 674052 626311
rect 674012 625864 674064 625870
rect 674012 625806 674064 625812
rect 674012 625592 674064 625598
rect 674010 625560 674012 625569
rect 674064 625560 674066 625569
rect 674010 625495 674066 625504
rect 674010 625152 674066 625161
rect 674010 625087 674012 625096
rect 674064 625087 674066 625096
rect 674012 625058 674064 625064
rect 674010 624744 674066 624753
rect 674010 624679 674012 624688
rect 674064 624679 674066 624688
rect 674012 624650 674064 624656
rect 674012 624368 674064 624374
rect 674010 624336 674012 624345
rect 674064 624336 674066 624345
rect 674010 624271 674066 624280
rect 674010 623928 674066 623937
rect 674010 623863 674012 623872
rect 674064 623863 674066 623872
rect 674012 623834 674064 623840
rect 674012 623552 674064 623558
rect 674010 623520 674012 623529
rect 674064 623520 674066 623529
rect 674010 623455 674066 623464
rect 674010 623112 674066 623121
rect 674010 623047 674012 623056
rect 674064 623047 674066 623056
rect 674012 623018 674064 623024
rect 674012 622736 674064 622742
rect 674010 622704 674012 622713
rect 674064 622704 674066 622713
rect 674010 622639 674066 622648
rect 674010 622296 674066 622305
rect 674010 622231 674012 622240
rect 674064 622231 674066 622240
rect 674012 622202 674064 622208
rect 674012 621240 674064 621246
rect 674010 621208 674012 621217
rect 674064 621208 674066 621217
rect 674010 621143 674066 621152
rect 674300 621014 674328 642518
rect 674470 640248 674526 640257
rect 674470 640183 674526 640192
rect 674484 637574 674512 640183
rect 674668 637574 674696 643266
rect 674392 637546 674512 637574
rect 674576 637546 674696 637574
rect 674392 630674 674420 637546
rect 674576 637022 674604 637546
rect 674564 637016 674616 637022
rect 674564 636958 674616 636964
rect 674392 630646 674512 630674
rect 674024 620986 674328 621014
rect 674024 611354 674052 620986
rect 674484 618225 674512 630646
rect 674760 626657 674788 649966
rect 675404 649777 675432 650012
rect 675390 649768 675446 649777
rect 675390 649703 675446 649712
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675772 648689 675800 648788
rect 675758 648680 675814 648689
rect 675758 648615 675814 648624
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 675114 647320 675170 647329
rect 675114 647255 675170 647264
rect 674932 645244 674984 645250
rect 674932 645186 674984 645192
rect 674944 642649 674972 645186
rect 675128 644489 675156 647255
rect 675312 645646 675418 645674
rect 675312 645250 675340 645646
rect 675300 645244 675352 645250
rect 675300 645186 675352 645192
rect 675312 645102 675418 645130
rect 675312 644745 675340 645102
rect 675298 644736 675354 644745
rect 675298 644671 675354 644680
rect 675128 644461 675418 644489
rect 675128 643810 675418 643838
rect 675128 643278 675156 643810
rect 675390 643648 675446 643657
rect 675390 643583 675446 643592
rect 675404 643280 675432 643583
rect 675116 643272 675168 643278
rect 675116 643214 675168 643220
rect 675114 643104 675170 643113
rect 675114 643039 675170 643048
rect 674852 642621 674972 642649
rect 674852 631938 674880 642621
rect 675128 641458 675156 643039
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 674944 640781 675418 640809
rect 674944 632210 674972 640781
rect 675312 640138 675418 640166
rect 674944 632182 675064 632210
rect 675036 631938 675064 632182
rect 674852 631910 674972 631938
rect 675036 631910 675156 631938
rect 674944 631854 674972 631910
rect 674932 631848 674984 631854
rect 674932 631790 674984 631796
rect 675128 631122 675156 631910
rect 674944 631094 675156 631122
rect 674746 626648 674802 626657
rect 674746 626583 674802 626592
rect 674944 626534 674972 631094
rect 675312 630850 675340 640138
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 675484 637016 675536 637022
rect 675484 636958 675536 636964
rect 675496 636585 675524 636958
rect 675852 636880 675904 636886
rect 675850 636848 675852 636857
rect 683396 636880 683448 636886
rect 675904 636848 675906 636857
rect 683396 636822 683448 636828
rect 675850 636783 675906 636792
rect 675482 636576 675538 636585
rect 675482 636511 675538 636520
rect 683210 636576 683266 636585
rect 683210 636511 683266 636520
rect 681002 636168 681058 636177
rect 681002 636103 681058 636112
rect 675484 631848 675536 631854
rect 675484 631790 675536 631796
rect 675128 630822 675340 630850
rect 674944 626506 675064 626534
rect 674470 618216 674526 618225
rect 674470 618151 674526 618160
rect 674024 611326 674144 611354
rect 673918 602984 673974 602993
rect 673918 602919 673974 602928
rect 673932 601694 673960 602919
rect 673656 592006 673776 592034
rect 673840 601666 673960 601694
rect 673656 591841 673684 592006
rect 673642 591832 673698 591841
rect 673642 591767 673698 591776
rect 673458 591288 673514 591297
rect 673458 591223 673514 591232
rect 673642 580680 673698 580689
rect 673642 580615 673698 580624
rect 673656 579698 673684 580615
rect 673644 579692 673696 579698
rect 673644 579634 673696 579640
rect 673458 579456 673514 579465
rect 673458 579391 673514 579400
rect 673472 578270 673500 579391
rect 673460 578264 673512 578270
rect 673460 578206 673512 578212
rect 673642 578232 673698 578241
rect 673642 578167 673698 578176
rect 673656 577182 673684 578167
rect 673644 577176 673696 577182
rect 673644 577118 673696 577124
rect 673414 577040 673466 577046
rect 673466 576988 673500 576994
rect 673414 576982 673500 576988
rect 673426 576966 673500 576982
rect 673472 576745 673500 576966
rect 673458 576736 673514 576745
rect 673458 576671 673514 576680
rect 673642 574560 673698 574569
rect 673642 574495 673698 574504
rect 673656 574190 673684 574495
rect 673644 574184 673696 574190
rect 673644 574126 673696 574132
rect 673642 572520 673698 572529
rect 673642 572455 673698 572464
rect 673656 571742 673684 572455
rect 673644 571736 673696 571742
rect 673644 571678 673696 571684
rect 673642 558104 673698 558113
rect 673642 558039 673698 558048
rect 673276 557864 673328 557870
rect 673276 557806 673328 557812
rect 673274 557560 673330 557569
rect 673274 557495 673330 557504
rect 673288 557410 673316 557495
rect 673104 557382 673316 557410
rect 673104 549250 673132 557382
rect 673276 555484 673328 555490
rect 673276 555426 673328 555432
rect 673104 549222 673224 549250
rect 673196 548962 673224 549222
rect 673288 549114 673316 555426
rect 673460 550656 673512 550662
rect 673460 550598 673512 550604
rect 673472 549273 673500 550598
rect 673458 549264 673514 549273
rect 673458 549199 673514 549208
rect 673288 549086 673408 549114
rect 673184 548956 673236 548962
rect 673184 548898 673236 548904
rect 673012 548814 673224 548842
rect 673000 548548 673052 548554
rect 673000 548490 673052 548496
rect 673012 539594 673040 548490
rect 672828 539566 672948 539594
rect 673012 539566 673132 539594
rect 672552 538186 672672 538214
rect 672448 531956 672500 531962
rect 672448 531898 672500 531904
rect 672264 528488 672316 528494
rect 672264 528430 672316 528436
rect 672460 488510 672488 531898
rect 672644 531758 672672 538186
rect 672632 531752 672684 531758
rect 672632 531694 672684 531700
rect 672724 530256 672776 530262
rect 672724 530198 672776 530204
rect 672736 526522 672764 530198
rect 672920 527649 672948 539566
rect 672906 527640 672962 527649
rect 672906 527575 672962 527584
rect 672724 526516 672776 526522
rect 672724 526458 672776 526464
rect 672908 493332 672960 493338
rect 672908 493274 672960 493280
rect 672920 491337 672948 493274
rect 672906 491328 672962 491337
rect 672906 491263 672962 491272
rect 672632 489660 672684 489666
rect 672632 489602 672684 489608
rect 672448 488504 672500 488510
rect 672448 488446 672500 488452
rect 671988 482384 672040 482390
rect 671988 482326 672040 482332
rect 671986 474872 672042 474881
rect 671986 474807 672042 474816
rect 670608 456408 670660 456414
rect 670608 456350 670660 456356
rect 669410 455424 669466 455433
rect 669410 455359 669466 455368
rect 672000 454866 672028 474807
rect 672000 454850 672120 454866
rect 672000 454844 672132 454850
rect 672000 454838 672080 454844
rect 672080 454786 672132 454792
rect 672448 453960 672500 453966
rect 672448 453902 672500 453908
rect 672460 453801 672488 453902
rect 672446 453792 672502 453801
rect 672446 453727 672502 453736
rect 60002 430672 60058 430681
rect 60002 430607 60058 430616
rect 45834 427408 45890 427417
rect 45834 427343 45890 427352
rect 45834 426864 45890 426873
rect 45834 426799 45890 426808
rect 45558 384840 45614 384849
rect 45558 384775 45614 384784
rect 45848 384033 45876 426799
rect 46018 424008 46074 424017
rect 46018 423943 46074 423952
rect 46032 400217 46060 423943
rect 53838 407824 53894 407833
rect 53838 407759 53894 407768
rect 53852 404326 53880 407759
rect 53840 404320 53892 404326
rect 53840 404262 53892 404268
rect 51080 400240 51132 400246
rect 46018 400208 46074 400217
rect 51080 400182 51132 400188
rect 46018 400143 46074 400152
rect 51092 395729 51120 400182
rect 60016 400110 60044 430607
rect 61382 429312 61438 429321
rect 61382 429247 61438 429256
rect 60004 400104 60056 400110
rect 60004 400046 60056 400052
rect 61396 398313 61424 429247
rect 63130 427136 63186 427145
rect 63130 427071 63186 427080
rect 62120 404320 62172 404326
rect 62120 404262 62172 404268
rect 62132 404161 62160 404262
rect 62118 404152 62174 404161
rect 62118 404087 62174 404096
rect 62120 402960 62172 402966
rect 62120 402902 62172 402908
rect 62132 402665 62160 402902
rect 62118 402656 62174 402665
rect 62118 402591 62174 402600
rect 62118 400616 62174 400625
rect 62118 400551 62174 400560
rect 62132 400246 62160 400551
rect 62120 400240 62172 400246
rect 63144 400217 63172 427071
rect 657542 403336 657598 403345
rect 657542 403271 657598 403280
rect 652022 400888 652078 400897
rect 652022 400823 652078 400832
rect 62120 400182 62172 400188
rect 63130 400208 63186 400217
rect 63130 400143 63186 400152
rect 62120 400104 62172 400110
rect 62120 400046 62172 400052
rect 62132 399401 62160 400046
rect 62118 399392 62174 399401
rect 62118 399327 62174 399336
rect 61382 398304 61438 398313
rect 61382 398239 61438 398248
rect 51078 395720 51134 395729
rect 51078 395655 51134 395664
rect 61382 386472 61438 386481
rect 61382 386407 61438 386416
rect 46018 384432 46074 384441
rect 46018 384367 46074 384376
rect 45834 384024 45890 384033
rect 45834 383959 45890 383968
rect 45650 383616 45706 383625
rect 45650 383551 45706 383560
rect 45282 381440 45338 381449
rect 45282 381375 45338 381384
rect 45296 369854 45324 381375
rect 44836 364306 44956 364334
rect 45020 369826 45140 369854
rect 45204 369826 45324 369854
rect 44546 361584 44602 361593
rect 44546 361519 44602 361528
rect 44192 359650 44680 359666
rect 44192 359644 44692 359650
rect 44192 359638 44640 359644
rect 44640 359586 44692 359592
rect 44836 359514 44864 364306
rect 44824 359508 44876 359514
rect 44824 359450 44876 359456
rect 44822 355192 44878 355201
rect 44822 355127 44878 355136
rect 44638 354920 44694 354929
rect 44638 354855 44694 354864
rect 44652 354754 44680 354855
rect 44836 354754 44864 355127
rect 44640 354748 44692 354754
rect 44640 354690 44692 354696
rect 44824 354748 44876 354754
rect 44824 354690 44876 354696
rect 43732 354606 43944 354634
rect 44008 354606 44895 354634
rect 43916 354498 43944 354606
rect 43916 354482 44772 354498
rect 44867 354482 44895 354606
rect 43916 354476 44784 354482
rect 43916 354470 44732 354476
rect 44732 354418 44784 354424
rect 44855 354476 44907 354482
rect 44855 354418 44907 354424
rect 43258 353696 43314 353705
rect 43258 353631 43314 353640
rect 42338 353016 42394 353025
rect 42338 352951 42394 352960
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35808 344616 35860 344622
rect 35808 344558 35860 344564
rect 39856 344616 39908 344622
rect 39856 344558 39908 344564
rect 35820 344321 35848 344558
rect 35806 344312 35862 344321
rect 35806 344247 35862 344256
rect 35622 343904 35678 343913
rect 35622 343839 35678 343848
rect 35636 343670 35664 343839
rect 35624 343664 35676 343670
rect 35624 343606 35676 343612
rect 35806 343496 35862 343505
rect 35806 343431 35862 343440
rect 35820 342242 35848 343431
rect 35808 342236 35860 342242
rect 35808 342178 35860 342184
rect 39868 341873 39896 344558
rect 40406 343904 40462 343913
rect 40406 343839 40462 343848
rect 40040 343664 40092 343670
rect 40040 343606 40092 343612
rect 35806 341864 35862 341873
rect 35806 341799 35862 341808
rect 39670 341864 39726 341873
rect 39670 341799 39726 341808
rect 39854 341864 39910 341873
rect 39854 341799 39910 341808
rect 35820 341562 35848 341799
rect 35808 341556 35860 341562
rect 35808 341498 35860 341504
rect 35808 341080 35860 341086
rect 35806 341048 35808 341057
rect 35860 341048 35862 341057
rect 35806 340983 35862 340992
rect 39684 340241 39712 341799
rect 40052 341442 40080 343606
rect 40222 342272 40278 342281
rect 40222 342207 40224 342216
rect 40276 342207 40278 342216
rect 40224 342178 40276 342184
rect 40420 341578 40448 343839
rect 45020 342553 45048 369826
rect 45204 343369 45232 369826
rect 45374 362944 45430 362953
rect 45374 362879 45430 362888
rect 45388 360194 45416 362879
rect 45376 360188 45428 360194
rect 45376 360130 45428 360136
rect 45376 359644 45428 359650
rect 45296 359592 45376 359598
rect 45296 359586 45428 359592
rect 45296 359570 45416 359586
rect 45296 353818 45324 359570
rect 45468 359508 45520 359514
rect 45468 359450 45520 359456
rect 45296 353790 45343 353818
rect 45315 353530 45343 353790
rect 45303 353524 45355 353530
rect 45303 353466 45355 353472
rect 45480 353274 45508 359450
rect 45434 353258 45508 353274
rect 45422 353252 45508 353258
rect 45474 353246 45508 353252
rect 45422 353194 45474 353200
rect 45190 343360 45246 343369
rect 45190 343295 45246 343304
rect 45006 342544 45062 342553
rect 45006 342479 45062 342488
rect 45466 342272 45522 342281
rect 45466 342207 45468 342216
rect 45520 342207 45522 342216
rect 45468 342178 45520 342184
rect 40236 341562 40448 341578
rect 40224 341556 40448 341562
rect 40276 341550 40448 341556
rect 40224 341498 40276 341504
rect 40052 341414 40540 341442
rect 40512 341306 40540 341414
rect 42246 341320 42302 341329
rect 40512 341278 42246 341306
rect 42246 341255 42302 341264
rect 40132 341080 40184 341086
rect 40130 341048 40132 341057
rect 40184 341048 40186 341057
rect 40130 340983 40186 340992
rect 45664 340785 45692 383551
rect 45834 353968 45890 353977
rect 45834 353903 45836 353912
rect 45888 353903 45890 353912
rect 45836 353874 45888 353880
rect 45836 353728 45888 353734
rect 45834 353696 45836 353705
rect 45888 353696 45890 353705
rect 45834 353631 45890 353640
rect 46032 343913 46060 384367
rect 47122 383208 47178 383217
rect 47122 383143 47178 383152
rect 46938 382392 46994 382401
rect 46938 382327 46994 382336
rect 46570 363216 46626 363225
rect 46570 363151 46626 363160
rect 46584 361554 46612 363151
rect 46572 361548 46624 361554
rect 46572 361490 46624 361496
rect 46952 353025 46980 382327
rect 47136 354385 47164 383143
rect 51724 357468 51776 357474
rect 51724 357410 51776 357416
rect 47122 354376 47178 354385
rect 47122 354311 47178 354320
rect 51736 353297 51764 357410
rect 61396 356017 61424 386407
rect 63406 385928 63462 385937
rect 63406 385863 63462 385872
rect 62946 381848 63002 381857
rect 62946 381783 63002 381792
rect 62120 361548 62172 361554
rect 62120 361490 62172 361496
rect 62132 360913 62160 361490
rect 62118 360904 62174 360913
rect 62118 360839 62174 360848
rect 62120 360188 62172 360194
rect 62120 360130 62172 360136
rect 62132 359825 62160 360130
rect 62118 359816 62174 359825
rect 62118 359751 62174 359760
rect 62118 357776 62174 357785
rect 62118 357711 62174 357720
rect 62132 357474 62160 357711
rect 62120 357468 62172 357474
rect 62120 357410 62172 357416
rect 61382 356008 61438 356017
rect 61382 355943 61438 355952
rect 62960 354521 62988 381783
rect 63420 357377 63448 385863
rect 651472 373992 651524 373998
rect 651472 373934 651524 373940
rect 651484 373289 651512 373934
rect 651470 373280 651526 373289
rect 651470 373215 651526 373224
rect 652036 372201 652064 400823
rect 652206 395312 652262 395321
rect 652206 395247 652262 395256
rect 652220 373969 652248 395247
rect 654782 382936 654838 382945
rect 654782 382871 654838 382880
rect 652206 373960 652262 373969
rect 652206 373895 652262 373904
rect 652022 372192 652078 372201
rect 652022 372127 652078 372136
rect 654796 371006 654824 382871
rect 657556 373998 657584 403271
rect 672644 401985 672672 489602
rect 673104 483177 673132 539566
rect 673196 531314 673224 548814
rect 673380 544490 673408 549086
rect 673288 544462 673408 544490
rect 673288 534074 673316 544462
rect 673458 535256 673514 535265
rect 673458 535191 673514 535200
rect 673472 534274 673500 535191
rect 673460 534268 673512 534274
rect 673460 534210 673512 534216
rect 673288 534046 673408 534074
rect 673380 531314 673408 534046
rect 673196 531286 673316 531314
rect 673380 531286 673500 531314
rect 673288 529145 673316 531286
rect 673472 530262 673500 531286
rect 673460 530256 673512 530262
rect 673460 530198 673512 530204
rect 673274 529136 673330 529145
rect 673274 529071 673330 529080
rect 673276 526516 673328 526522
rect 673276 526458 673328 526464
rect 673090 483168 673146 483177
rect 673090 483103 673146 483112
rect 673288 455870 673316 526458
rect 673656 484401 673684 558039
rect 673840 556646 673868 601666
rect 674116 599842 674144 611326
rect 674838 600128 674894 600137
rect 674838 600063 674894 600072
rect 674116 599814 674236 599842
rect 674208 599298 674236 599814
rect 674562 599448 674618 599457
rect 674562 599383 674618 599392
rect 674024 599270 674236 599298
rect 674024 581641 674052 599270
rect 674378 598360 674434 598369
rect 674378 598295 674434 598304
rect 674194 597408 674250 597417
rect 674194 597343 674250 597352
rect 674010 581632 674066 581641
rect 674010 581567 674066 581576
rect 674010 581088 674066 581097
rect 674010 581023 674012 581032
rect 674064 581023 674066 581032
rect 674012 580994 674064 581000
rect 674012 580304 674064 580310
rect 674010 580272 674012 580281
rect 674064 580272 674066 580281
rect 674010 580207 674066 580216
rect 674012 580032 674064 580038
rect 674012 579974 674064 579980
rect 674024 579873 674052 579974
rect 674010 579864 674066 579873
rect 674010 579799 674066 579808
rect 674010 579048 674066 579057
rect 674010 578983 674066 578992
rect 674024 578814 674052 578983
rect 674012 578808 674064 578814
rect 674012 578750 674064 578756
rect 674010 578640 674066 578649
rect 674010 578575 674066 578584
rect 674024 578406 674052 578575
rect 674012 578400 674064 578406
rect 674012 578342 674064 578348
rect 674012 577448 674064 577454
rect 674010 577416 674012 577425
rect 674064 577416 674066 577425
rect 674010 577351 674066 577360
rect 674010 577008 674066 577017
rect 674010 576943 674012 576952
rect 674064 576943 674066 576952
rect 674012 576914 674064 576920
rect 674012 575952 674064 575958
rect 674012 575894 674064 575900
rect 674024 575793 674052 575894
rect 674010 575784 674066 575793
rect 674010 575719 674066 575728
rect 674012 574456 674064 574462
rect 674012 574398 674064 574404
rect 674024 574161 674052 574398
rect 674010 574152 674066 574161
rect 674010 574087 674066 574096
rect 674010 572928 674066 572937
rect 674010 572863 674012 572872
rect 674064 572863 674066 572872
rect 674012 572834 674064 572840
rect 674010 572112 674066 572121
rect 674010 572047 674066 572056
rect 674024 571470 674052 572047
rect 674012 571464 674064 571470
rect 674012 571406 674064 571412
rect 674012 565888 674064 565894
rect 674010 565856 674012 565865
rect 674064 565856 674066 565865
rect 674010 565791 674066 565800
rect 673828 556640 673880 556646
rect 673828 556582 673880 556588
rect 674012 556640 674064 556646
rect 674012 556582 674064 556588
rect 674024 555642 674052 556582
rect 674024 555614 674144 555642
rect 673918 555520 673974 555529
rect 673918 555455 673974 555464
rect 673932 555234 673960 555455
rect 673748 555206 673960 555234
rect 673748 543734 673776 555206
rect 674116 554962 674144 555614
rect 673932 554934 674144 554962
rect 673932 554933 673960 554934
rect 673840 554905 673960 554933
rect 673840 547074 673868 554905
rect 674012 554872 674064 554878
rect 674012 554814 674064 554820
rect 674024 554713 674052 554814
rect 674010 554704 674066 554713
rect 674010 554639 674066 554648
rect 674012 553444 674064 553450
rect 674208 553394 674236 597343
rect 674064 553392 674144 553394
rect 674012 553386 674144 553392
rect 674024 553366 674144 553386
rect 674208 553366 674328 553394
rect 674116 552945 674144 553366
rect 674102 552936 674158 552945
rect 674102 552871 674158 552880
rect 674300 552786 674328 553366
rect 674208 552758 674328 552786
rect 674208 550338 674236 552758
rect 674392 551253 674420 598295
rect 674576 582374 674604 599383
rect 674852 598641 674880 600063
rect 674838 598632 674894 598641
rect 674838 598567 674894 598576
rect 675036 595898 675064 626506
rect 674760 595870 675064 595898
rect 674760 592929 674788 595870
rect 675128 595762 675156 630822
rect 675496 626534 675524 631790
rect 675850 626648 675906 626657
rect 675850 626583 675906 626592
rect 675220 626506 675524 626534
rect 675220 599162 675248 626506
rect 675864 623082 675892 626583
rect 675852 623076 675904 623082
rect 675852 623018 675904 623024
rect 681016 622033 681044 636103
rect 683224 634814 683252 636511
rect 683224 634786 683344 634814
rect 683120 623076 683172 623082
rect 683120 623018 683172 623024
rect 681002 622024 681058 622033
rect 681002 621959 681058 621968
rect 683132 617545 683160 623018
rect 683316 622962 683344 634786
rect 683224 622934 683344 622962
rect 683224 617794 683252 622934
rect 683408 617953 683436 636822
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683394 617944 683450 617953
rect 683394 617879 683450 617888
rect 683224 617766 683344 617794
rect 683118 617536 683174 617545
rect 683118 617471 683174 617480
rect 683316 617137 683344 617766
rect 683302 617128 683358 617137
rect 683302 617063 683358 617072
rect 675850 616856 675906 616865
rect 675850 616791 675906 616800
rect 675864 615534 675892 616791
rect 675852 615528 675904 615534
rect 683120 615528 683172 615534
rect 675852 615470 675904 615476
rect 683118 615496 683120 615505
rect 683172 615496 683174 615505
rect 683118 615431 683174 615440
rect 675390 611416 675446 611425
rect 675390 611351 675446 611360
rect 675404 608668 675432 611351
rect 675390 608288 675446 608297
rect 675390 608223 675446 608232
rect 675404 608124 675432 608223
rect 675390 608016 675446 608025
rect 675390 607951 675446 607960
rect 675404 607479 675432 607951
rect 675404 606529 675432 606832
rect 675390 606520 675446 606529
rect 675390 606455 675446 606464
rect 675496 604625 675524 604996
rect 675482 604616 675538 604625
rect 675482 604551 675538 604560
rect 675404 604353 675432 604452
rect 675390 604344 675446 604353
rect 675390 604279 675446 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 675404 602993 675432 603160
rect 675390 602984 675446 602993
rect 675390 602919 675446 602928
rect 675496 600409 675524 600644
rect 675482 600400 675538 600409
rect 675482 600335 675538 600344
rect 675772 599865 675800 600100
rect 675758 599856 675814 599865
rect 675758 599791 675814 599800
rect 675482 599720 675538 599729
rect 675482 599655 675538 599664
rect 675496 599488 675524 599655
rect 675482 599176 675538 599185
rect 675220 599134 675482 599162
rect 675482 599111 675538 599120
rect 675298 599040 675354 599049
rect 675298 598975 675354 598984
rect 675312 596442 675340 598975
rect 675772 598641 675800 598808
rect 675482 598632 675538 598641
rect 675482 598567 675538 598576
rect 675758 598632 675814 598641
rect 675758 598567 675814 598576
rect 675496 598264 675524 598567
rect 675496 597417 675524 597652
rect 675482 597408 675538 597417
rect 675482 597343 675538 597352
rect 675312 596414 675418 596442
rect 675298 596320 675354 596329
rect 675298 596255 675354 596264
rect 675312 596174 675340 596255
rect 674944 595734 675156 595762
rect 675220 596146 675340 596174
rect 674746 592920 674802 592929
rect 674746 592855 674802 592864
rect 674944 589257 674972 595734
rect 675220 595218 675248 596146
rect 675404 595513 675432 595816
rect 675390 595504 675446 595513
rect 675390 595439 675446 595448
rect 675036 595190 675248 595218
rect 675036 592034 675064 595190
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675404 593609 675432 593980
rect 675390 593600 675446 593609
rect 675390 593535 675446 593544
rect 675850 592920 675906 592929
rect 675850 592855 675852 592864
rect 675904 592855 675906 592864
rect 678244 592884 678296 592890
rect 675852 592826 675904 592832
rect 678244 592826 678296 592832
rect 675482 592104 675538 592113
rect 675482 592039 675538 592048
rect 675036 592006 675156 592034
rect 674930 589248 674986 589257
rect 674930 589183 674986 589192
rect 675128 586265 675156 592006
rect 675496 586265 675524 592039
rect 675850 591832 675906 591841
rect 675850 591767 675906 591776
rect 675864 591462 675892 591767
rect 675852 591456 675904 591462
rect 675852 591398 675904 591404
rect 675852 591320 675904 591326
rect 675850 591288 675852 591297
rect 675904 591288 675906 591297
rect 675850 591223 675906 591232
rect 675852 589280 675904 589286
rect 675850 589248 675852 589257
rect 675904 589248 675906 589257
rect 675850 589183 675906 589192
rect 675114 586256 675170 586265
rect 675114 586191 675170 586200
rect 675482 586256 675538 586265
rect 675482 586191 675538 586200
rect 674116 550310 674236 550338
rect 674300 551225 674420 551253
rect 674484 582346 674604 582374
rect 674116 547346 674144 550310
rect 674300 547466 674328 551225
rect 674288 547460 674340 547466
rect 674288 547402 674340 547408
rect 674116 547318 674328 547346
rect 674300 547194 674328 547318
rect 674288 547188 674340 547194
rect 674288 547130 674340 547136
rect 673840 547058 674328 547074
rect 673840 547052 674340 547058
rect 673840 547046 674288 547052
rect 674288 546994 674340 547000
rect 673748 543706 674052 543734
rect 674024 538214 674052 543706
rect 674024 538186 674328 538214
rect 673826 536072 673882 536081
rect 673826 536007 673882 536016
rect 673840 535498 673868 536007
rect 674012 535696 674064 535702
rect 674010 535664 674012 535673
rect 674064 535664 674066 535673
rect 674010 535599 674066 535608
rect 673828 535492 673880 535498
rect 673828 535434 673880 535440
rect 674010 534848 674066 534857
rect 674010 534783 674066 534792
rect 674024 534546 674052 534783
rect 674012 534540 674064 534546
rect 674012 534482 674064 534488
rect 673826 534440 673882 534449
rect 673826 534375 673882 534384
rect 674012 534404 674064 534410
rect 673840 534138 673868 534375
rect 674012 534346 674064 534352
rect 674024 534177 674052 534346
rect 674010 534168 674066 534177
rect 673828 534132 673880 534138
rect 674010 534103 674066 534112
rect 673828 534074 673880 534080
rect 674010 533624 674066 533633
rect 674010 533559 674012 533568
rect 674064 533559 674066 533568
rect 674012 533530 674064 533536
rect 674012 533384 674064 533390
rect 674010 533352 674012 533361
rect 674064 533352 674066 533361
rect 674010 533287 674066 533296
rect 674010 532808 674066 532817
rect 674010 532743 674012 532752
rect 674064 532743 674066 532752
rect 674012 532714 674064 532720
rect 674012 532568 674064 532574
rect 674010 532536 674012 532545
rect 674064 532536 674066 532545
rect 674010 532471 674066 532480
rect 674010 531992 674066 532001
rect 674010 531927 674012 531936
rect 674064 531927 674066 531936
rect 674012 531898 674064 531904
rect 674012 531752 674064 531758
rect 674010 531720 674012 531729
rect 674064 531720 674066 531729
rect 674010 531655 674066 531664
rect 674010 531176 674066 531185
rect 674010 531111 674066 531120
rect 673828 530120 673880 530126
rect 673826 530088 673828 530097
rect 673880 530088 673882 530097
rect 673826 530023 673882 530032
rect 674024 529990 674052 531111
rect 674012 529984 674064 529990
rect 674012 529926 674064 529932
rect 674012 529712 674064 529718
rect 674010 529680 674012 529689
rect 674064 529680 674066 529689
rect 674010 529615 674066 529624
rect 674300 529258 674328 538186
rect 674484 537169 674512 582346
rect 674654 581632 674710 581641
rect 674654 581567 674710 581576
rect 674668 571441 674696 581567
rect 675850 577824 675906 577833
rect 675850 577759 675906 577768
rect 675864 576745 675892 577759
rect 675850 576736 675906 576745
rect 675850 576671 675906 576680
rect 678256 576473 678284 592826
rect 684038 592648 684094 592657
rect 684038 592583 684094 592592
rect 683396 591456 683448 591462
rect 683396 591398 683448 591404
rect 681004 589280 681056 589286
rect 681004 589222 681056 589228
rect 678242 576464 678298 576473
rect 678242 576399 678298 576408
rect 674654 571432 674710 571441
rect 674654 571367 674710 571376
rect 681016 571334 681044 589222
rect 683408 571985 683436 591398
rect 684052 575657 684080 592583
rect 684224 591320 684276 591326
rect 684224 591262 684276 591268
rect 684038 575648 684094 575657
rect 684038 575583 684094 575592
rect 684236 574025 684264 591262
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 684222 574016 684278 574025
rect 684222 573951 684278 573960
rect 683394 571976 683450 571985
rect 683394 571911 683450 571920
rect 681004 571328 681056 571334
rect 681004 571270 681056 571276
rect 683120 571328 683172 571334
rect 683120 571270 683172 571276
rect 683132 570761 683160 571270
rect 683118 570752 683174 570761
rect 683118 570687 683174 570696
rect 676218 569528 676274 569537
rect 676218 569463 676274 569472
rect 675390 565856 675446 565865
rect 675390 565791 675446 565800
rect 675404 563448 675432 565791
rect 676232 565593 676260 569463
rect 676218 565584 676274 565593
rect 676218 565519 676274 565528
rect 675772 562737 675800 562904
rect 675758 562728 675814 562737
rect 675758 562663 675814 562672
rect 675114 562320 675170 562329
rect 675170 562278 675418 562306
rect 675114 562255 675170 562264
rect 675390 561912 675446 561921
rect 675390 561847 675446 561856
rect 675404 561612 675432 561847
rect 675312 559830 675432 559858
rect 675312 559790 675340 559830
rect 674852 559762 675340 559790
rect 675404 559776 675432 559830
rect 674656 554940 674708 554946
rect 674656 554882 674708 554888
rect 674470 537160 674526 537169
rect 674470 537095 674526 537104
rect 674300 529230 674420 529258
rect 674010 529136 674066 529145
rect 674010 529071 674066 529080
rect 674024 528630 674052 529071
rect 674012 528624 674064 528630
rect 674012 528566 674064 528572
rect 674012 528488 674064 528494
rect 674010 528456 674012 528465
rect 674064 528456 674066 528465
rect 674010 528391 674066 528400
rect 674012 524680 674064 524686
rect 674010 524648 674012 524657
rect 674064 524648 674066 524657
rect 674010 524583 674066 524592
rect 674392 524414 674420 529230
rect 674392 524386 674512 524414
rect 674484 505094 674512 524386
rect 674392 505066 674512 505094
rect 674392 492425 674420 505066
rect 674378 492416 674434 492425
rect 674378 492351 674434 492360
rect 673826 492144 673882 492153
rect 673826 492079 673882 492088
rect 673840 491366 673868 492079
rect 674010 491736 674066 491745
rect 674010 491671 674066 491680
rect 674024 491502 674052 491671
rect 674012 491496 674064 491502
rect 674012 491438 674064 491444
rect 673828 491360 673880 491366
rect 673828 491302 673880 491308
rect 674012 490952 674064 490958
rect 674010 490920 674012 490929
rect 674064 490920 674066 490929
rect 674010 490855 674066 490864
rect 674012 490136 674064 490142
rect 674010 490104 674012 490113
rect 674064 490104 674066 490113
rect 674010 490039 674066 490048
rect 674010 489696 674066 489705
rect 674010 489631 674012 489640
rect 674064 489631 674066 489640
rect 674012 489602 674064 489608
rect 674012 489320 674064 489326
rect 674010 489288 674012 489297
rect 674064 489288 674066 489297
rect 674010 489223 674066 489232
rect 674012 488504 674064 488510
rect 674010 488472 674012 488481
rect 674064 488472 674066 488481
rect 674010 488407 674066 488416
rect 674010 486024 674066 486033
rect 674010 485959 674066 485968
rect 674024 485858 674052 485959
rect 674012 485852 674064 485858
rect 674012 485794 674064 485800
rect 673826 485616 673882 485625
rect 673826 485551 673882 485560
rect 673840 484430 673868 485551
rect 674010 485208 674066 485217
rect 674010 485143 674066 485152
rect 674024 484566 674052 485143
rect 674012 484560 674064 484566
rect 674012 484502 674064 484508
rect 673828 484424 673880 484430
rect 673642 484392 673698 484401
rect 673828 484366 673880 484372
rect 673642 484327 673698 484336
rect 674668 482769 674696 554882
rect 674852 553466 674880 559762
rect 675128 559218 675418 559246
rect 675128 555529 675156 559218
rect 675404 558113 675432 558620
rect 675390 558104 675446 558113
rect 675390 558039 675446 558048
rect 675404 557569 675432 557940
rect 675390 557560 675446 557569
rect 675390 557495 675446 557504
rect 675114 555520 675170 555529
rect 675114 555455 675170 555464
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675116 554940 675168 554946
rect 675168 554905 675418 554933
rect 675116 554882 675168 554888
rect 675114 554704 675170 554713
rect 675114 554639 675170 554648
rect 674760 553438 674880 553466
rect 674760 553330 674788 553438
rect 674760 553302 675064 553330
rect 674838 549808 674894 549817
rect 674838 549743 674894 549752
rect 674654 482760 674710 482769
rect 674654 482695 674710 482704
rect 674012 482384 674064 482390
rect 674010 482352 674012 482361
rect 674064 482352 674066 482361
rect 674010 482287 674066 482296
rect 674852 480049 674880 549743
rect 675036 501945 675064 553302
rect 675128 553093 675156 554639
rect 675772 553897 675800 554268
rect 675758 553888 675814 553897
rect 675758 553823 675814 553832
rect 675404 553489 675432 553656
rect 675390 553480 675446 553489
rect 675390 553415 675446 553424
rect 675128 553065 675418 553093
rect 675206 552936 675262 552945
rect 675206 552871 675262 552880
rect 675220 551253 675248 552871
rect 675772 552129 675800 552432
rect 675758 552120 675814 552129
rect 675758 552055 675814 552064
rect 675220 551225 675418 551253
rect 675128 550582 675418 550610
rect 675128 511994 675156 550582
rect 675404 549817 675432 549951
rect 675390 549808 675446 549817
rect 675390 549743 675446 549752
rect 675390 549264 675446 549273
rect 675390 549199 675446 549208
rect 675404 548760 675432 549199
rect 675482 547632 675538 547641
rect 676034 547632 676090 547641
rect 675482 547567 675484 547576
rect 675536 547567 675538 547576
rect 675852 547596 675904 547602
rect 675484 547538 675536 547544
rect 676034 547567 676090 547576
rect 677414 547632 677470 547641
rect 677414 547567 677470 547576
rect 684224 547596 684276 547602
rect 675852 547538 675904 547544
rect 675864 547448 675892 547538
rect 676048 547466 676076 547567
rect 675496 547420 675892 547448
rect 676036 547460 676088 547466
rect 675496 547330 675524 547420
rect 676036 547402 676088 547408
rect 675484 547324 675536 547330
rect 675484 547266 675536 547272
rect 675852 547324 675904 547330
rect 675852 547266 675904 547272
rect 675864 547210 675892 547266
rect 675496 547182 675892 547210
rect 675496 547058 675524 547182
rect 675484 547052 675536 547058
rect 675484 546994 675536 547000
rect 675298 544504 675354 544513
rect 675298 544439 675354 544448
rect 675312 511994 675340 544439
rect 675850 537160 675906 537169
rect 675850 537095 675906 537104
rect 675864 533390 675892 537095
rect 675852 533384 675904 533390
rect 675852 533326 675904 533332
rect 675850 524648 675906 524657
rect 675850 524583 675852 524592
rect 675904 524583 675906 524592
rect 675852 524554 675904 524560
rect 675852 518900 675904 518906
rect 675852 518842 675904 518848
rect 675574 513768 675630 513777
rect 675574 513703 675630 513712
rect 675128 511966 675248 511994
rect 675312 511966 675432 511994
rect 675220 508881 675248 511966
rect 675206 508872 675262 508881
rect 675206 508807 675262 508816
rect 675404 507226 675432 511966
rect 675312 507198 675432 507226
rect 675312 503946 675340 507198
rect 675588 505594 675616 513703
rect 675496 505566 675616 505594
rect 675496 503946 675524 505566
rect 675300 503940 675352 503946
rect 675300 503882 675352 503888
rect 675484 503940 675536 503946
rect 675484 503882 675536 503888
rect 675300 503668 675352 503674
rect 675300 503610 675352 503616
rect 675484 503668 675536 503674
rect 675484 503610 675536 503616
rect 675022 501936 675078 501945
rect 675022 501871 675078 501880
rect 675312 487665 675340 503610
rect 675298 487656 675354 487665
rect 675298 487591 675354 487600
rect 675114 481944 675170 481953
rect 675114 481879 675170 481888
rect 674838 480040 674894 480049
rect 674838 479975 674894 479984
rect 673458 464808 673514 464817
rect 673458 464743 673514 464752
rect 673276 455864 673328 455870
rect 673276 455806 673328 455812
rect 673274 455424 673330 455433
rect 673274 455359 673276 455368
rect 673328 455359 673330 455368
rect 673276 455330 673328 455336
rect 673472 455274 673500 464743
rect 673828 455864 673880 455870
rect 673826 455832 673828 455841
rect 673880 455832 673882 455841
rect 673826 455767 673882 455776
rect 673400 455258 673500 455274
rect 673388 455252 673500 455258
rect 673440 455246 673500 455252
rect 673388 455194 673440 455200
rect 673276 455048 673328 455054
rect 673274 455016 673276 455025
rect 673328 455016 673330 455025
rect 673274 454951 673330 454960
rect 673046 454640 673098 454646
rect 673044 454608 673046 454617
rect 673098 454608 673100 454617
rect 673044 454543 673100 454552
rect 672954 454368 673006 454374
rect 672952 454336 672954 454345
rect 674288 454368 674340 454374
rect 673006 454336 673008 454345
rect 672952 454271 673008 454280
rect 674286 454336 674288 454345
rect 674340 454336 674342 454345
rect 674286 454271 674342 454280
rect 672816 454096 672868 454102
rect 672814 454064 672816 454073
rect 672868 454064 672870 454073
rect 672814 453999 672870 454008
rect 675128 453801 675156 481879
rect 675298 480720 675354 480729
rect 675298 480655 675354 480664
rect 675312 454073 675340 480655
rect 675496 454374 675524 503610
rect 675864 502334 675892 518842
rect 676036 518696 676088 518702
rect 676036 518638 676088 518644
rect 676048 513777 676076 518638
rect 676034 513768 676090 513777
rect 676034 513703 676090 513712
rect 676126 508872 676182 508881
rect 676126 508807 676182 508816
rect 676140 503810 676168 508807
rect 676128 503804 676180 503810
rect 676128 503746 676180 503752
rect 677428 503674 677456 547567
rect 684224 547538 684276 547544
rect 683396 547460 683448 547466
rect 683396 547402 683448 547408
rect 678242 547360 678298 547369
rect 678242 547295 678298 547304
rect 683212 547324 683264 547330
rect 678256 530641 678284 547295
rect 683212 547266 683264 547272
rect 681002 547088 681058 547097
rect 681002 547023 681058 547032
rect 681016 531049 681044 547023
rect 681002 531040 681058 531049
rect 681002 530975 681058 530984
rect 678242 530632 678298 530641
rect 678242 530567 678298 530576
rect 683224 527377 683252 547266
rect 683210 527368 683266 527377
rect 683210 527303 683266 527312
rect 683408 526561 683436 547402
rect 683580 533384 683632 533390
rect 683580 533326 683632 533332
rect 683592 526969 683620 533326
rect 684236 528193 684264 547538
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 684222 528184 684278 528193
rect 684222 528119 684278 528128
rect 683578 526960 683634 526969
rect 683578 526895 683634 526904
rect 683394 526552 683450 526561
rect 683394 526487 683450 526496
rect 677874 525736 677930 525745
rect 677874 525671 677930 525680
rect 677690 524512 677746 524521
rect 677690 524447 677746 524456
rect 677704 518906 677732 524447
rect 677692 518900 677744 518906
rect 677692 518842 677744 518848
rect 677888 518838 677916 525671
rect 683118 524920 683174 524929
rect 683118 524855 683174 524864
rect 683132 524618 683160 524855
rect 683120 524612 683172 524618
rect 683120 524554 683172 524560
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 678244 503804 678296 503810
rect 678244 503746 678296 503752
rect 677416 503668 677468 503674
rect 677416 503610 677468 503616
rect 675680 502306 675892 502334
rect 675680 454617 675708 502306
rect 675850 501936 675906 501945
rect 675850 501871 675906 501880
rect 675864 500818 675892 501871
rect 675852 500812 675904 500818
rect 675852 500754 675904 500760
rect 676034 492416 676090 492425
rect 676034 492351 676090 492360
rect 675850 490512 675906 490521
rect 675850 490447 675906 490456
rect 675864 485774 675892 490447
rect 676048 490074 676076 492351
rect 676036 490068 676088 490074
rect 676036 490010 676088 490016
rect 676588 490068 676640 490074
rect 676588 490010 676640 490016
rect 676034 488064 676090 488073
rect 676090 488022 676260 488050
rect 676034 487999 676090 488008
rect 676232 487218 676260 488022
rect 676220 487212 676272 487218
rect 676220 487154 676272 487160
rect 675864 485746 675984 485774
rect 675666 454608 675722 454617
rect 675666 454543 675722 454552
rect 675484 454368 675536 454374
rect 675484 454310 675536 454316
rect 675298 454064 675354 454073
rect 675298 453999 675354 454008
rect 675114 453792 675170 453801
rect 675114 453727 675170 453736
rect 675956 447817 675984 485746
rect 676600 484571 676628 490010
rect 678256 487257 678284 503746
rect 683396 503668 683448 503674
rect 683396 503610 683448 503616
rect 681004 500812 681056 500818
rect 681004 500754 681056 500760
rect 678242 487248 678298 487257
rect 677508 487212 677560 487218
rect 678242 487183 678298 487192
rect 677508 487154 677560 487160
rect 676586 484562 676642 484571
rect 676586 484497 676642 484506
rect 676128 480412 676180 480418
rect 676128 480354 676180 480360
rect 676140 480049 676168 480354
rect 676126 480040 676182 480049
rect 676126 479975 676182 479984
rect 676218 477456 676274 477465
rect 676218 477391 676274 477400
rect 676232 456210 676260 477391
rect 676220 456204 676272 456210
rect 676220 456146 676272 456152
rect 676174 456000 676226 456006
rect 676140 455948 676174 455954
rect 676140 455942 676226 455948
rect 676140 455926 676214 455942
rect 676140 455841 676168 455926
rect 676126 455832 676182 455841
rect 676126 455767 676182 455776
rect 675942 447808 675998 447817
rect 675942 447743 675998 447752
rect 677520 440337 677548 487154
rect 681016 486441 681044 500754
rect 683408 486849 683436 503610
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683394 486840 683450 486849
rect 683394 486775 683450 486784
rect 681002 486432 681058 486441
rect 681002 486367 681058 486376
rect 683118 481128 683174 481137
rect 683118 481063 683174 481072
rect 683132 480418 683160 481063
rect 683120 480412 683172 480418
rect 683120 480354 683172 480360
rect 677506 440328 677562 440337
rect 677506 440263 677562 440272
rect 676034 410544 676090 410553
rect 676034 410479 676090 410488
rect 674562 403472 674618 403481
rect 674562 403407 674618 403416
rect 672630 401976 672686 401985
rect 672630 401911 672686 401920
rect 672814 401704 672870 401713
rect 672814 401639 672870 401648
rect 671986 397216 672042 397225
rect 671986 397151 672042 397160
rect 669226 393544 669282 393553
rect 669226 393479 669282 393488
rect 668858 386064 668914 386073
rect 668858 385999 668914 386008
rect 668872 382945 668900 385999
rect 668858 382936 668914 382945
rect 668858 382871 668914 382880
rect 657544 373992 657596 373998
rect 657544 373934 657596 373940
rect 651472 371000 651524 371006
rect 651472 370942 651524 370948
rect 654784 371000 654836 371006
rect 654784 370942 654836 370948
rect 651484 370705 651512 370942
rect 651470 370696 651526 370705
rect 651470 370631 651526 370640
rect 654782 358592 654838 358601
rect 654782 358527 654838 358536
rect 63406 357368 63462 357377
rect 63406 357303 63462 357312
rect 652022 356688 652078 356697
rect 652022 356623 652078 356632
rect 62946 354512 63002 354521
rect 62946 354447 63002 354456
rect 51722 353288 51778 353297
rect 51722 353223 51778 353232
rect 46938 353016 46994 353025
rect 46938 352951 46994 352960
rect 46018 343904 46074 343913
rect 46018 343839 46074 343848
rect 63132 342236 63184 342242
rect 63132 342178 63184 342184
rect 62946 341728 63002 341737
rect 62946 341663 63002 341672
rect 62762 341456 62818 341465
rect 62762 341391 62818 341400
rect 45650 340776 45706 340785
rect 45650 340711 45706 340720
rect 39670 340232 39726 340241
rect 39670 340167 39726 340176
rect 35530 339824 35586 339833
rect 35530 339759 35586 339768
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35544 339658 35572 339759
rect 35532 339652 35584 339658
rect 35532 339594 35584 339600
rect 35820 339522 35848 339759
rect 37096 339652 37148 339658
rect 37096 339594 37148 339600
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 37108 336569 37136 339594
rect 38844 339516 38896 339522
rect 38844 339458 38896 339464
rect 37094 336560 37150 336569
rect 37094 336495 37150 336504
rect 38856 335753 38884 339458
rect 46938 339280 46994 339289
rect 46938 339215 46994 339224
rect 45558 338872 45614 338881
rect 45558 338807 45614 338816
rect 45374 337920 45430 337929
rect 45374 337855 45430 337864
rect 45388 337770 45416 337855
rect 45388 337742 45508 337770
rect 35806 335744 35862 335753
rect 35806 335679 35862 335688
rect 38842 335744 38898 335753
rect 38842 335679 38898 335688
rect 35820 335374 35848 335679
rect 35808 335368 35860 335374
rect 35808 335310 35860 335316
rect 39856 335368 39908 335374
rect 39856 335310 39908 335316
rect 35806 334520 35862 334529
rect 35806 334455 35862 334464
rect 35820 334150 35848 334455
rect 35808 334144 35860 334150
rect 35808 334086 35860 334092
rect 39868 332489 39896 335310
rect 44178 334656 44234 334665
rect 44178 334591 44234 334600
rect 44362 334656 44418 334665
rect 44362 334591 44418 334600
rect 40316 334144 40368 334150
rect 40316 334086 40368 334092
rect 40328 332897 40356 334086
rect 40314 332888 40370 332897
rect 40314 332823 40370 332832
rect 42890 332888 42946 332897
rect 42890 332823 42946 332832
rect 39854 332480 39910 332489
rect 39854 332415 39910 332424
rect 42430 327040 42486 327049
rect 42430 326975 42486 326984
rect 42444 326278 42472 326975
rect 42168 326210 42196 326264
rect 42260 326250 42472 326278
rect 42260 326210 42288 326250
rect 42168 326182 42288 326210
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42182 323734 42656 323762
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42182 321898 42472 321926
rect 42076 321201 42104 321368
rect 42062 321192 42118 321201
rect 42062 321127 42118 321136
rect 42168 320521 42196 320725
rect 42154 320512 42210 320521
rect 42154 320447 42210 320456
rect 42076 319977 42104 320076
rect 41878 319968 41934 319977
rect 41878 319903 41934 319912
rect 42062 319968 42118 319977
rect 42062 319903 42118 319912
rect 41892 319532 41920 319903
rect 42444 319705 42472 321898
rect 42628 320793 42656 323734
rect 42904 321201 42932 332823
rect 43074 332480 43130 332489
rect 43074 332415 43130 332424
rect 42890 321192 42946 321201
rect 42890 321127 42946 321136
rect 42614 320784 42670 320793
rect 42614 320719 42670 320728
rect 43088 320521 43116 332415
rect 43074 320512 43130 320521
rect 43074 320447 43130 320456
rect 44192 319977 44220 334591
rect 44376 322833 44404 334591
rect 45282 327040 45338 327049
rect 45480 327026 45508 337742
rect 45338 326998 45508 327026
rect 45282 326975 45338 326984
rect 44362 322824 44418 322833
rect 44362 322759 44418 322768
rect 44178 319968 44234 319977
rect 44178 319903 44234 319912
rect 42430 319696 42486 319705
rect 42430 319631 42486 319640
rect 42246 319016 42302 319025
rect 42246 318951 42302 318960
rect 41786 317384 41842 317393
rect 41786 317319 41842 317328
rect 41800 317045 41828 317319
rect 42260 316418 42288 318951
rect 42182 316390 42288 316418
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 42168 315757 42196 315959
rect 45572 315489 45600 338807
rect 42154 315480 42210 315489
rect 42154 315415 42210 315424
rect 45558 315480 45614 315489
rect 45558 315415 45614 315424
rect 42168 315180 42196 315415
rect 42062 313712 42118 313721
rect 42062 313647 42118 313656
rect 42076 313344 42104 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 42168 312174 42288 312202
rect 42168 312052 42196 312174
rect 42260 312066 42288 312174
rect 42260 312038 42472 312066
rect 42076 309097 42104 311508
rect 42444 310457 42472 312038
rect 46952 310457 46980 339215
rect 51722 334112 51778 334121
rect 51722 334047 51778 334056
rect 50342 333160 50398 333169
rect 50342 333095 50398 333104
rect 42430 310448 42486 310457
rect 42430 310383 42486 310392
rect 46938 310448 46994 310457
rect 46938 310383 46994 310392
rect 42062 309088 42118 309097
rect 42062 309023 42118 309032
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 35622 300928 35678 300937
rect 35622 300863 35678 300872
rect 35636 298790 35664 300863
rect 46202 300520 46258 300529
rect 46202 300455 46258 300464
rect 44178 299704 44234 299713
rect 44178 299639 44234 299648
rect 35806 298888 35862 298897
rect 35806 298823 35862 298832
rect 35624 298784 35676 298790
rect 35624 298726 35676 298732
rect 35820 298314 35848 298823
rect 41604 298784 41656 298790
rect 41786 298752 41842 298761
rect 41656 298732 41786 298738
rect 41604 298726 41786 298732
rect 41616 298710 41786 298726
rect 41786 298687 41842 298696
rect 35808 298308 35860 298314
rect 35808 298250 35860 298256
rect 41604 298308 41656 298314
rect 41604 298250 41656 298256
rect 41616 296562 41644 298250
rect 41786 296576 41842 296585
rect 41616 296534 41786 296562
rect 41786 296511 41842 296520
rect 42798 296576 42854 296585
rect 42798 296511 42854 296520
rect 35438 296440 35494 296449
rect 35438 296375 35494 296384
rect 35452 295526 35480 296375
rect 35622 296032 35678 296041
rect 35622 295967 35678 295976
rect 35440 295520 35492 295526
rect 35440 295462 35492 295468
rect 35636 295390 35664 295967
rect 35808 295656 35860 295662
rect 35806 295624 35808 295633
rect 40684 295656 40736 295662
rect 35860 295624 35862 295633
rect 40684 295598 40736 295604
rect 35806 295559 35862 295568
rect 35624 295384 35676 295390
rect 35624 295326 35676 295332
rect 35806 295216 35862 295225
rect 35806 295151 35862 295160
rect 33782 294808 33838 294817
rect 33782 294743 33838 294752
rect 32402 294400 32458 294409
rect 32402 294335 32458 294344
rect 32416 284889 32444 294335
rect 33796 286346 33824 294743
rect 35820 294166 35848 295151
rect 35808 294160 35860 294166
rect 35808 294102 35860 294108
rect 35806 293176 35862 293185
rect 35806 293111 35862 293120
rect 35820 292942 35848 293111
rect 35808 292936 35860 292942
rect 35808 292878 35860 292884
rect 35806 292768 35862 292777
rect 35806 292703 35862 292712
rect 35820 292602 35848 292703
rect 35808 292596 35860 292602
rect 35808 292538 35860 292544
rect 35806 291136 35862 291145
rect 35806 291071 35862 291080
rect 35622 290320 35678 290329
rect 35622 290255 35678 290264
rect 35636 289134 35664 290255
rect 35820 289950 35848 291071
rect 35808 289944 35860 289950
rect 35808 289886 35860 289892
rect 35624 289128 35676 289134
rect 35624 289070 35676 289076
rect 33784 286340 33836 286346
rect 33784 286282 33836 286288
rect 32402 284880 32458 284889
rect 32402 284815 32458 284824
rect 40696 284345 40724 295598
rect 41328 295520 41380 295526
rect 41328 295462 41380 295468
rect 41340 292482 41368 295462
rect 41604 295384 41656 295390
rect 41786 295352 41842 295361
rect 41656 295332 41786 295338
rect 41604 295326 41786 295332
rect 41616 295310 41786 295326
rect 41786 295287 41842 295296
rect 41696 294160 41748 294166
rect 41696 294102 41748 294108
rect 41512 292868 41564 292874
rect 41512 292810 41564 292816
rect 41340 292454 41460 292482
rect 41432 292346 41460 292454
rect 41524 292448 41552 292810
rect 41708 292574 41736 294102
rect 41708 292546 42564 292574
rect 42064 292460 42116 292466
rect 41524 292420 42064 292448
rect 42064 292402 42116 292408
rect 41432 292318 42472 292346
rect 41604 292256 41656 292262
rect 41786 292224 41842 292233
rect 41656 292204 41786 292210
rect 41604 292198 41786 292204
rect 41616 292182 41786 292198
rect 41786 292159 41842 292168
rect 41786 291952 41842 291961
rect 41524 291910 41786 291938
rect 41524 289814 41552 291910
rect 41786 291887 41842 291896
rect 41786 290320 41842 290329
rect 41786 290255 41842 290264
rect 41800 290170 41828 290255
rect 41708 290154 41828 290170
rect 41696 290148 41828 290154
rect 41748 290142 41828 290148
rect 41696 290090 41748 290096
rect 41524 289786 41828 289814
rect 41800 289241 41828 289786
rect 41786 289232 41842 289241
rect 41786 289167 41842 289176
rect 41696 289060 41748 289066
rect 41696 289002 41748 289008
rect 41708 288946 41736 289002
rect 41708 288918 42380 288946
rect 41696 286340 41748 286346
rect 41696 286282 41748 286288
rect 41708 286226 41736 286282
rect 41708 286198 42288 286226
rect 40682 284336 40738 284345
rect 40682 284271 40738 284280
rect 42260 283059 42288 286198
rect 42182 283031 42288 283059
rect 42352 281874 42380 288918
rect 42182 281846 42380 281874
rect 42168 281302 42288 281330
rect 42168 281180 42196 281302
rect 42260 281194 42288 281302
rect 42444 281194 42472 292318
rect 42536 282914 42564 292546
rect 42536 282886 42656 282914
rect 42260 281166 42472 281194
rect 42182 280554 42472 280582
rect 42248 280152 42300 280158
rect 42248 280094 42300 280100
rect 42260 279426 42288 280094
rect 42168 279398 42288 279426
rect 42168 279344 42196 279398
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42182 278718 42288 278746
rect 41786 278488 41842 278497
rect 41786 278423 41842 278432
rect 41800 278188 41828 278423
rect 42062 277808 42118 277817
rect 42062 277743 42118 277752
rect 42076 277508 42104 277743
rect 41786 277128 41842 277137
rect 41786 277063 41842 277072
rect 41800 276896 41828 277063
rect 42062 276720 42118 276729
rect 42062 276655 42118 276664
rect 42076 276352 42104 276655
rect 42260 275913 42288 278718
rect 42430 278695 42486 278704
rect 42628 276729 42656 282886
rect 42614 276720 42670 276729
rect 42614 276655 42670 276664
rect 42246 275904 42302 275913
rect 42246 275839 42302 275848
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42168 273170 42196 273224
rect 42338 273184 42394 273193
rect 42168 273142 42338 273170
rect 42338 273119 42394 273128
rect 42430 272912 42486 272921
rect 42430 272847 42486 272856
rect 42444 272558 42472 272847
rect 42182 272530 42472 272558
rect 41970 272368 42026 272377
rect 41970 272303 42026 272312
rect 41984 272000 42012 272303
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 41878 270056 41934 270065
rect 41878 269991 41934 270000
rect 41892 269521 41920 269991
rect 42156 269068 42208 269074
rect 42156 269010 42208 269016
rect 42168 268872 42196 269010
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 42168 266257 42196 268328
rect 42154 266248 42210 266257
rect 42154 266183 42210 266192
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 42812 255921 42840 296511
rect 43166 295352 43222 295361
rect 43166 295287 43222 295296
rect 42984 292460 43036 292466
rect 42984 292402 43036 292408
rect 42996 280158 43024 292402
rect 42984 280152 43036 280158
rect 42984 280094 43036 280100
rect 43180 269074 43208 295287
rect 43626 292224 43682 292233
rect 43626 292159 43682 292168
rect 43350 290320 43406 290329
rect 43350 290255 43406 290264
rect 43364 282914 43392 290255
rect 43364 282886 43484 282914
rect 43168 269068 43220 269074
rect 43168 269010 43220 269016
rect 35806 255912 35862 255921
rect 35806 255847 35862 255856
rect 39762 255912 39818 255921
rect 39762 255847 39818 255856
rect 42798 255912 42854 255921
rect 42798 255847 42854 255856
rect 35820 255474 35848 255847
rect 39776 255474 39804 255847
rect 35808 255468 35860 255474
rect 35808 255410 35860 255416
rect 39764 255468 39816 255474
rect 39764 255410 39816 255416
rect 35808 254108 35860 254114
rect 35808 254050 35860 254056
rect 39580 254108 39632 254114
rect 39580 254050 39632 254056
rect 35820 253881 35848 254050
rect 39592 253881 39620 254050
rect 35806 253872 35862 253881
rect 35806 253807 35862 253816
rect 39578 253872 39634 253881
rect 39578 253807 39634 253816
rect 42798 253872 42854 253881
rect 42798 253807 42854 253816
rect 35622 253464 35678 253473
rect 35622 253399 35678 253408
rect 35636 252618 35664 253399
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 40958 253056 41014 253065
rect 40958 252991 41014 253000
rect 35820 252754 35848 252991
rect 35808 252748 35860 252754
rect 35808 252690 35860 252696
rect 40972 252618 41000 252991
rect 41696 252748 41748 252754
rect 41696 252690 41748 252696
rect 35624 252612 35676 252618
rect 35624 252554 35676 252560
rect 40960 252612 41012 252618
rect 40960 252554 41012 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 40498 252240 40554 252249
rect 40498 252175 40554 252184
rect 35820 251394 35848 252175
rect 40512 251394 40540 252175
rect 35808 251388 35860 251394
rect 35808 251330 35860 251336
rect 40500 251388 40552 251394
rect 40500 251330 40552 251336
rect 35806 250608 35862 250617
rect 35806 250543 35862 250552
rect 35820 249966 35848 250543
rect 35808 249960 35860 249966
rect 35808 249902 35860 249908
rect 39396 249960 39448 249966
rect 39396 249902 39448 249908
rect 39408 249393 39436 249902
rect 35806 249384 35862 249393
rect 35806 249319 35862 249328
rect 39394 249384 39450 249393
rect 39394 249319 39450 249328
rect 35820 248538 35848 249319
rect 41708 248554 41736 252690
rect 42430 252240 42486 252249
rect 42430 252175 42486 252184
rect 35808 248532 35860 248538
rect 35808 248474 35860 248480
rect 39212 248532 39264 248538
rect 41708 248526 42380 248554
rect 39212 248474 39264 248480
rect 35622 247752 35678 247761
rect 35622 247687 35678 247696
rect 35636 247110 35664 247687
rect 35808 247240 35860 247246
rect 35808 247182 35860 247188
rect 35624 247104 35676 247110
rect 35624 247046 35676 247052
rect 35820 246945 35848 247182
rect 35806 246936 35862 246945
rect 35806 246871 35862 246880
rect 39224 245041 39252 248474
rect 41696 247240 41748 247246
rect 41696 247182 41748 247188
rect 41512 247104 41564 247110
rect 41512 247046 41564 247052
rect 41524 246945 41552 247046
rect 41510 246936 41566 246945
rect 41510 246871 41566 246880
rect 39210 245032 39266 245041
rect 39210 244967 39266 244976
rect 41708 244274 41736 247182
rect 41708 244246 42288 244274
rect 42062 240136 42118 240145
rect 42062 240071 42118 240080
rect 42076 239836 42104 240071
rect 42260 238754 42288 244246
rect 42168 238726 42288 238754
rect 42168 238649 42196 238726
rect 42352 238014 42380 248526
rect 42182 237986 42380 238014
rect 42444 237425 42472 252175
rect 42812 251174 42840 253807
rect 43258 253056 43314 253065
rect 43258 252991 43314 253000
rect 42720 251146 42840 251174
rect 43272 251174 43300 252991
rect 43272 251146 43392 251174
rect 42720 241514 42748 251146
rect 43166 249384 43222 249393
rect 43166 249319 43222 249328
rect 42982 245032 43038 245041
rect 42982 244967 43038 244976
rect 42720 241486 42840 241514
rect 42430 237416 42486 237425
rect 42430 237351 42486 237360
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42430 235920 42486 235929
rect 42430 235855 42486 235864
rect 42444 234983 42472 235855
rect 42182 234955 42472 234983
rect 42432 234592 42484 234598
rect 42432 234534 42484 234540
rect 42444 234342 42472 234534
rect 42182 234314 42472 234342
rect 42182 233667 42472 233695
rect 42444 233481 42472 233667
rect 42430 233472 42486 233481
rect 42430 233407 42486 233416
rect 42430 233200 42486 233209
rect 42168 233158 42430 233186
rect 42168 233104 42196 233158
rect 42430 233135 42486 233144
rect 42246 233064 42302 233073
rect 42246 232999 42302 233008
rect 42062 231024 42118 231033
rect 42062 230959 42118 230968
rect 42076 230656 42104 230959
rect 42260 230466 42288 232999
rect 42168 230438 42288 230466
rect 42432 230444 42484 230450
rect 42168 229976 42196 230438
rect 42432 230386 42484 230392
rect 42444 229378 42472 230386
rect 42182 229350 42472 229378
rect 41970 228984 42026 228993
rect 41970 228919 42026 228928
rect 41984 228820 42012 228919
rect 42432 227724 42484 227730
rect 42432 227666 42484 227672
rect 42444 226998 42472 227666
rect 42168 226930 42196 226984
rect 42260 226970 42472 226998
rect 42260 226930 42288 226970
rect 42168 226902 42288 226930
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42260 226290 42472 226318
rect 42246 226128 42302 226137
rect 42246 226063 42302 226072
rect 42260 225706 42288 226063
rect 42182 225678 42288 225706
rect 42168 223281 42196 225148
rect 42444 224913 42472 226290
rect 42614 225584 42670 225593
rect 42614 225519 42670 225528
rect 42430 224904 42486 224913
rect 42430 224839 42486 224848
rect 42154 223272 42210 223281
rect 42154 223207 42210 223216
rect 42628 219434 42656 225519
rect 41708 219406 42656 219434
rect 35806 217968 35862 217977
rect 35806 217903 35862 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35820 214713 35848 217903
rect 35806 214704 35862 214713
rect 35806 214639 35862 214648
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 41708 213994 41736 219406
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 41696 213988 41748 213994
rect 41696 213930 41748 213936
rect 35438 212256 35494 212265
rect 35438 212191 35494 212200
rect 35452 211206 35480 212191
rect 42812 211857 42840 241486
rect 42996 234598 43024 244967
rect 42984 234592 43036 234598
rect 42984 234534 43036 234540
rect 43180 230466 43208 249319
rect 43364 244274 43392 251146
rect 43088 230450 43208 230466
rect 43076 230444 43208 230450
rect 43128 230438 43208 230444
rect 43272 244246 43392 244274
rect 43076 230386 43128 230392
rect 43272 227730 43300 244246
rect 43260 227724 43312 227730
rect 43260 227666 43312 227672
rect 43456 215294 43484 282886
rect 43640 277817 43668 292159
rect 43626 277808 43682 277817
rect 43626 277743 43682 277752
rect 44192 256873 44220 299639
rect 45006 298072 45062 298081
rect 45006 298007 45062 298016
rect 44362 297256 44418 297265
rect 44362 297191 44418 297200
rect 44178 256864 44234 256873
rect 44178 256799 44234 256808
rect 44376 254425 44404 297191
rect 44730 293992 44786 294001
rect 44730 293927 44786 293936
rect 44546 293584 44602 293593
rect 44546 293519 44602 293528
rect 44560 273193 44588 293519
rect 44546 273184 44602 273193
rect 44546 273119 44602 273128
rect 44744 272921 44772 293927
rect 44730 272912 44786 272921
rect 44730 272847 44786 272856
rect 44822 256456 44878 256465
rect 44822 256391 44878 256400
rect 44638 254824 44694 254833
rect 44638 254759 44694 254768
rect 44362 254416 44418 254425
rect 44362 254351 44418 254360
rect 44362 252784 44418 252793
rect 44362 252719 44418 252728
rect 44178 251560 44234 251569
rect 44178 251495 44234 251504
rect 43626 246936 43682 246945
rect 43626 246871 43682 246880
rect 43456 215266 43576 215294
rect 35622 211848 35678 211857
rect 35622 211783 35678 211792
rect 39578 211848 39634 211857
rect 39578 211783 39634 211792
rect 42798 211848 42854 211857
rect 42798 211783 42854 211792
rect 35636 211342 35664 211783
rect 39592 211614 39620 211783
rect 35808 211608 35860 211614
rect 35808 211550 35860 211556
rect 39580 211608 39632 211614
rect 39580 211550 39632 211556
rect 35820 211449 35848 211550
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35624 211336 35676 211342
rect 35624 211278 35676 211284
rect 41696 211336 41748 211342
rect 41696 211278 41748 211284
rect 35440 211200 35492 211206
rect 35440 211142 35492 211148
rect 41328 211200 41380 211206
rect 41328 211142 41380 211148
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35820 209846 35848 210151
rect 35808 209840 35860 209846
rect 35808 209782 35860 209788
rect 40224 209840 40276 209846
rect 40224 209782 40276 209788
rect 35622 208992 35678 209001
rect 35622 208927 35678 208936
rect 35636 208418 35664 208927
rect 35806 208584 35862 208593
rect 35806 208519 35808 208528
rect 35860 208519 35862 208528
rect 35808 208490 35860 208496
rect 35624 208412 35676 208418
rect 35624 208354 35676 208360
rect 40040 208412 40092 208418
rect 40040 208354 40092 208360
rect 40052 208185 40080 208354
rect 40038 208176 40094 208185
rect 40038 208111 40094 208120
rect 35806 207768 35862 207777
rect 35806 207703 35862 207712
rect 35820 207194 35848 207703
rect 35808 207188 35860 207194
rect 35808 207130 35860 207136
rect 35806 206136 35862 206145
rect 35806 206071 35862 206080
rect 35820 205834 35848 206071
rect 35808 205828 35860 205834
rect 35808 205770 35860 205776
rect 40236 205737 40264 209782
rect 40500 208548 40552 208554
rect 40500 208490 40552 208496
rect 40512 207777 40540 208490
rect 40498 207768 40554 207777
rect 40498 207703 40554 207712
rect 40776 207188 40828 207194
rect 40776 207130 40828 207136
rect 40222 205728 40278 205737
rect 40222 205663 40278 205672
rect 35622 204912 35678 204921
rect 35622 204847 35678 204856
rect 35636 204338 35664 204847
rect 35808 204604 35860 204610
rect 35808 204546 35860 204552
rect 40408 204604 40460 204610
rect 40408 204546 40460 204552
rect 35624 204332 35676 204338
rect 35624 204274 35676 204280
rect 35820 204105 35848 204546
rect 40420 204105 40448 204546
rect 35806 204096 35862 204105
rect 35806 204031 35862 204040
rect 40406 204096 40462 204105
rect 40406 204031 40462 204040
rect 28538 203688 28594 203697
rect 28538 203623 28594 203632
rect 28552 199345 28580 203623
rect 40788 203289 40816 207130
rect 41340 206553 41368 211142
rect 41708 208185 41736 211278
rect 41694 208176 41750 208185
rect 41694 208111 41750 208120
rect 42982 207768 43038 207777
rect 42982 207703 43038 207712
rect 41326 206544 41382 206553
rect 41326 206479 41382 206488
rect 40960 205828 41012 205834
rect 40960 205770 41012 205776
rect 40972 204513 41000 205770
rect 40958 204504 41014 204513
rect 40958 204439 41014 204448
rect 41696 204400 41748 204406
rect 42064 204400 42116 204406
rect 41748 204348 42064 204354
rect 41696 204342 42116 204348
rect 41708 204326 42104 204342
rect 40774 203280 40830 203289
rect 40774 203215 40830 203224
rect 42798 203280 42854 203289
rect 42798 203215 42854 203224
rect 28538 199336 28594 199345
rect 28538 199271 28594 199280
rect 42246 199336 42302 199345
rect 42246 199271 42302 199280
rect 42062 197024 42118 197033
rect 42062 196959 42118 196968
rect 42076 196656 42104 196959
rect 42260 195786 42288 199271
rect 42168 195758 42288 195786
rect 42168 195432 42196 195758
rect 41878 195256 41934 195265
rect 41878 195191 41934 195200
rect 41892 194820 41920 195191
rect 42246 194984 42302 194993
rect 42246 194919 42302 194928
rect 41786 193216 41842 193225
rect 41786 193151 41842 193160
rect 41800 192984 41828 193151
rect 42076 191593 42104 191760
rect 42062 191584 42118 191593
rect 42062 191519 42118 191528
rect 42168 191026 42196 191148
rect 42260 191026 42288 194919
rect 42168 190998 42288 191026
rect 42246 190904 42302 190913
rect 42246 190839 42302 190848
rect 42260 190482 42288 190839
rect 42182 190454 42288 190482
rect 42432 190188 42484 190194
rect 42432 190130 42484 190136
rect 42444 189938 42472 190130
rect 42182 189910 42472 189938
rect 42432 187672 42484 187678
rect 42432 187614 42484 187620
rect 42444 187459 42472 187614
rect 42182 187431 42472 187459
rect 42430 186824 42486 186833
rect 42182 186782 42430 186810
rect 42430 186759 42486 186768
rect 41786 186416 41842 186425
rect 41786 186351 41842 186360
rect 41800 186184 41828 186351
rect 41786 186008 41842 186017
rect 41786 185943 41842 185952
rect 41800 185605 41828 185943
rect 41786 184104 41842 184113
rect 41786 184039 41842 184048
rect 41800 183765 41828 184039
rect 42812 183274 42840 203215
rect 42996 190194 43024 207703
rect 43166 204504 43222 204513
rect 43166 204439 43222 204448
rect 42984 190188 43036 190194
rect 42984 190130 43036 190136
rect 43180 187678 43208 204439
rect 43352 204400 43404 204406
rect 43350 204368 43352 204377
rect 43404 204368 43406 204377
rect 43350 204303 43406 204312
rect 43548 195974 43576 215266
rect 43456 195946 43576 195974
rect 43168 187672 43220 187678
rect 43168 187614 43220 187620
rect 42536 183246 42840 183274
rect 42536 183138 42564 183246
rect 42182 183110 42564 183138
rect 42182 182463 42472 182491
rect 42076 179353 42104 181900
rect 42444 180713 42472 182463
rect 42430 180704 42486 180713
rect 42430 180639 42486 180648
rect 42062 179344 42118 179353
rect 42062 179279 42118 179288
rect 43456 44198 43484 195946
rect 43640 44334 43668 246871
rect 44192 240145 44220 251495
rect 44178 240136 44234 240145
rect 44178 240071 44234 240080
rect 44376 226137 44404 252719
rect 44362 226128 44418 226137
rect 44362 226063 44418 226072
rect 44652 212129 44680 254759
rect 44836 213761 44864 256391
rect 45020 255241 45048 298007
rect 46216 292466 46244 300455
rect 46204 292460 46256 292466
rect 46204 292402 46256 292408
rect 48962 289912 49018 289921
rect 48962 289847 49018 289856
rect 46204 285728 46256 285734
rect 46204 285670 46256 285676
rect 46216 258097 46244 285670
rect 47768 280356 47820 280362
rect 47768 280298 47820 280304
rect 46202 258088 46258 258097
rect 46202 258023 46258 258032
rect 45558 255640 45614 255649
rect 45558 255575 45614 255584
rect 45006 255232 45062 255241
rect 45006 255167 45062 255176
rect 45006 251968 45062 251977
rect 45006 251903 45062 251912
rect 45020 233209 45048 251903
rect 45190 249112 45246 249121
rect 45190 249047 45246 249056
rect 45006 233200 45062 233209
rect 45006 233135 45062 233144
rect 45204 231033 45232 249047
rect 45190 231024 45246 231033
rect 45190 230959 45246 230968
rect 44822 213752 44878 213761
rect 44822 213687 44878 213696
rect 45572 212945 45600 255575
rect 45926 251152 45982 251161
rect 45926 251087 45982 251096
rect 45742 248704 45798 248713
rect 45742 248639 45798 248648
rect 45756 233481 45784 248639
rect 45742 233472 45798 233481
rect 45742 233407 45798 233416
rect 45940 224913 45968 251087
rect 46110 248296 46166 248305
rect 46110 248231 46166 248240
rect 46124 235929 46152 248231
rect 47582 246664 47638 246673
rect 47582 246599 47638 246608
rect 46110 235920 46166 235929
rect 46110 235855 46166 235864
rect 45926 224904 45982 224913
rect 45926 224839 45982 224848
rect 45558 212936 45614 212945
rect 45558 212871 45614 212880
rect 44638 212120 44694 212129
rect 44638 212055 44694 212064
rect 46938 209672 46994 209681
rect 46938 209607 46994 209616
rect 44362 208448 44418 208457
rect 44362 208383 44418 208392
rect 44178 207224 44234 207233
rect 44178 207159 44234 207168
rect 43994 204368 44050 204377
rect 43994 204303 44050 204312
rect 43810 204096 43866 204105
rect 43810 204031 43866 204040
rect 43824 45218 43852 204031
rect 44008 191593 44036 204303
rect 43994 191584 44050 191593
rect 43994 191519 44050 191528
rect 44192 186833 44220 207159
rect 44376 197033 44404 208383
rect 44638 205320 44694 205329
rect 44638 205255 44694 205264
rect 44362 197024 44418 197033
rect 44362 196959 44418 196968
rect 44652 190913 44680 205255
rect 44822 204912 44878 204921
rect 44822 204847 44878 204856
rect 44638 190904 44694 190913
rect 44638 190839 44694 190848
rect 44178 186824 44234 186833
rect 44178 186759 44234 186768
rect 44836 74534 44864 204847
rect 46202 203552 46258 203561
rect 46202 203487 46258 203496
rect 44836 74506 45508 74534
rect 45480 49026 45508 74506
rect 46216 51746 46244 203487
rect 46952 180713 46980 209607
rect 46938 180704 46994 180713
rect 46938 180639 46994 180648
rect 47596 53106 47624 246599
rect 47780 214985 47808 280298
rect 47766 214976 47822 214985
rect 47766 214911 47822 214920
rect 47766 213344 47822 213353
rect 47766 213279 47822 213288
rect 47780 190505 47808 213279
rect 47950 210896 48006 210905
rect 47950 210831 48006 210840
rect 47964 195922 47992 210831
rect 48778 206544 48834 206553
rect 48778 206479 48834 206488
rect 47964 195894 48360 195922
rect 48332 194449 48360 195894
rect 48318 194440 48374 194449
rect 48318 194375 48374 194384
rect 48792 192409 48820 206479
rect 48778 192400 48834 192409
rect 48778 192335 48834 192344
rect 47766 190496 47822 190505
rect 47766 190431 47822 190440
rect 48976 53242 49004 289847
rect 49146 247480 49202 247489
rect 49146 247415 49202 247424
rect 48964 53236 49016 53242
rect 48964 53178 49016 53184
rect 47584 53100 47636 53106
rect 47584 53042 47636 53048
rect 46204 51740 46256 51746
rect 46204 51682 46256 51688
rect 49160 50386 49188 247415
rect 49514 208176 49570 208185
rect 49514 208111 49570 208120
rect 49528 196489 49556 208111
rect 49514 196480 49570 196489
rect 49514 196415 49570 196424
rect 50356 51882 50384 333095
rect 50526 290728 50582 290737
rect 50526 290663 50582 290672
rect 50540 53378 50568 290663
rect 50712 218884 50764 218890
rect 50712 218826 50764 218832
rect 50724 179353 50752 218826
rect 50710 179344 50766 179353
rect 50710 179279 50766 179288
rect 50528 53372 50580 53378
rect 50528 53314 50580 53320
rect 50344 51876 50396 51882
rect 50344 51818 50396 51824
rect 49148 50380 49200 50386
rect 49148 50322 49200 50328
rect 51736 49162 51764 334047
rect 53838 320784 53894 320793
rect 53838 320719 53894 320728
rect 53102 319696 53158 319705
rect 53102 319631 53158 319640
rect 53116 315994 53144 319631
rect 53852 317422 53880 320719
rect 53840 317416 53892 317422
rect 62120 317416 62172 317422
rect 53840 317358 53892 317364
rect 62118 317384 62120 317393
rect 62172 317384 62174 317393
rect 62118 317319 62174 317328
rect 62118 316024 62174 316033
rect 53104 315988 53156 315994
rect 62118 315959 62120 315968
rect 53104 315930 53156 315936
rect 62172 315959 62174 315968
rect 62120 315930 62172 315936
rect 62118 314800 62174 314809
rect 59912 314764 59964 314770
rect 62118 314735 62120 314744
rect 59912 314706 59964 314712
rect 62172 314735 62174 314744
rect 62120 314706 62172 314712
rect 59924 309097 59952 314706
rect 62776 311817 62804 341391
rect 62960 313041 62988 341663
rect 63144 314129 63172 342178
rect 651380 328296 651432 328302
rect 651380 328238 651432 328244
rect 651392 328137 651420 328238
rect 651378 328128 651434 328137
rect 651378 328063 651434 328072
rect 652036 326913 652064 356623
rect 652390 352608 652446 352617
rect 652390 352543 652446 352552
rect 652404 329769 652432 352543
rect 653402 338736 653458 338745
rect 653402 338671 653458 338680
rect 652390 329760 652446 329769
rect 652390 329695 652446 329704
rect 652022 326904 652078 326913
rect 652022 326839 652078 326848
rect 651378 325680 651434 325689
rect 653416 325650 653444 338671
rect 654796 328302 654824 358527
rect 658922 346488 658978 346497
rect 658922 346423 658978 346432
rect 654784 328296 654836 328302
rect 654784 328238 654836 328244
rect 651378 325615 651380 325624
rect 651432 325615 651434 325624
rect 653404 325644 653456 325650
rect 651380 325586 651432 325592
rect 653404 325586 653456 325592
rect 63130 314120 63186 314129
rect 63130 314055 63186 314064
rect 653402 313304 653458 313313
rect 653402 313239 653458 313248
rect 62946 313032 63002 313041
rect 62946 312967 63002 312976
rect 62762 311808 62818 311817
rect 62762 311743 62818 311752
rect 652298 309904 652354 309913
rect 652298 309839 652354 309848
rect 59910 309088 59966 309097
rect 59910 309023 59966 309032
rect 651380 303544 651432 303550
rect 651380 303486 651432 303492
rect 651392 303385 651420 303486
rect 651378 303376 651434 303385
rect 651378 303311 651434 303320
rect 652312 302161 652340 309839
rect 653416 303550 653444 313239
rect 653404 303544 653456 303550
rect 653404 303486 653456 303492
rect 652298 302152 652354 302161
rect 652298 302087 652354 302096
rect 53102 301336 53158 301345
rect 53102 301271 53158 301280
rect 53116 291174 53144 301271
rect 654782 300928 654838 300937
rect 654782 300863 654838 300872
rect 651472 300824 651524 300830
rect 651472 300766 651524 300772
rect 651484 300665 651512 300766
rect 651470 300656 651526 300665
rect 651470 300591 651526 300600
rect 62762 298752 62818 298761
rect 62762 298687 62818 298696
rect 651470 298752 651526 298761
rect 651470 298687 651526 298696
rect 62118 295488 62174 295497
rect 58624 295452 58676 295458
rect 62118 295423 62120 295432
rect 58624 295394 58676 295400
rect 62172 295423 62174 295432
rect 62120 295394 62172 295400
rect 57244 294092 57296 294098
rect 57244 294034 57296 294040
rect 54484 292596 54536 292602
rect 54484 292538 54536 292544
rect 53104 291168 53156 291174
rect 53104 291110 53156 291116
rect 54496 266257 54524 292538
rect 55864 288516 55916 288522
rect 55864 288458 55916 288464
rect 54482 266248 54538 266257
rect 54482 266183 54538 266192
rect 55876 223281 55904 288458
rect 57256 275913 57284 294034
rect 58636 278769 58664 295394
rect 62118 294128 62174 294137
rect 62118 294063 62120 294072
rect 62172 294063 62174 294072
rect 62120 294034 62172 294040
rect 62302 292768 62358 292777
rect 62302 292703 62358 292712
rect 62316 292602 62344 292703
rect 62304 292596 62356 292602
rect 62304 292538 62356 292544
rect 62118 292496 62174 292505
rect 62118 292431 62120 292440
rect 62172 292431 62174 292440
rect 62120 292402 62172 292408
rect 62120 291168 62172 291174
rect 62120 291110 62172 291116
rect 62132 291009 62160 291110
rect 62118 291000 62174 291009
rect 62118 290935 62174 290944
rect 62776 289785 62804 298687
rect 651484 298178 651512 298687
rect 651472 298172 651524 298178
rect 651472 298114 651524 298120
rect 651470 297528 651526 297537
rect 651470 297463 651526 297472
rect 651484 297090 651512 297463
rect 651472 297084 651524 297090
rect 651472 297026 651524 297032
rect 652666 296848 652722 296857
rect 652666 296783 652722 296792
rect 652680 296002 652708 296783
rect 652668 295996 652720 296002
rect 652668 295938 652720 295944
rect 652114 295352 652170 295361
rect 652114 295287 652170 295296
rect 651470 294264 651526 294273
rect 651470 294199 651526 294208
rect 651484 294030 651512 294199
rect 651472 294024 651524 294030
rect 651472 293966 651524 293972
rect 651470 293040 651526 293049
rect 651470 292975 651526 292984
rect 651484 292602 651512 292975
rect 651472 292596 651524 292602
rect 651472 292538 651524 292544
rect 651470 290456 651526 290465
rect 651470 290391 651526 290400
rect 651484 289882 651512 290391
rect 651472 289876 651524 289882
rect 651472 289818 651524 289824
rect 62762 289776 62818 289785
rect 62762 289711 62818 289720
rect 651470 289232 651526 289241
rect 651470 289167 651526 289176
rect 62118 288552 62174 288561
rect 62118 288487 62120 288496
rect 62172 288487 62174 288496
rect 62120 288458 62172 288464
rect 651484 288454 651512 289167
rect 651746 288552 651802 288561
rect 651746 288487 651802 288496
rect 651472 288448 651524 288454
rect 651472 288390 651524 288396
rect 651470 287464 651526 287473
rect 651470 287399 651526 287408
rect 63130 287192 63186 287201
rect 63130 287127 63186 287136
rect 62118 285968 62174 285977
rect 62118 285903 62174 285912
rect 62132 285734 62160 285903
rect 62120 285728 62172 285734
rect 62120 285670 62172 285676
rect 62118 284472 62174 284481
rect 60004 284436 60056 284442
rect 62118 284407 62120 284416
rect 60004 284378 60056 284384
rect 62172 284407 62174 284416
rect 62120 284378 62172 284384
rect 58622 278760 58678 278769
rect 58622 278695 58678 278704
rect 57242 275904 57298 275913
rect 57242 275839 57298 275848
rect 60016 256737 60044 284378
rect 62762 283248 62818 283257
rect 62762 283183 62818 283192
rect 62118 280936 62174 280945
rect 62118 280871 62174 280880
rect 61382 280392 61438 280401
rect 62132 280362 62160 280871
rect 61382 280327 61438 280336
rect 62120 280356 62172 280362
rect 60002 256728 60058 256737
rect 60002 256663 60058 256672
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 55862 223272 55918 223281
rect 55862 223207 55918 223216
rect 56520 218210 56548 226986
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 55692 217138 55720 218146
rect 57256 218074 57284 228346
rect 60648 227452 60700 227458
rect 60648 227394 60700 227400
rect 58992 225616 59044 225622
rect 58992 225558 59044 225564
rect 57428 218204 57480 218210
rect 57428 218146 57480 218152
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56520 217138 56548 218010
rect 57440 217274 57468 218146
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217246 57468 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217246
rect 58176 217138 58204 218010
rect 59004 217274 59032 225558
rect 59360 221468 59412 221474
rect 59360 221410 59412 221416
rect 59372 218074 59400 221410
rect 59820 218748 59872 218754
rect 59820 218690 59872 218696
rect 59360 218068 59412 218074
rect 59360 218010 59412 218016
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218690
rect 60660 217274 60688 227394
rect 61396 219434 61424 280327
rect 62120 280298 62172 280304
rect 61660 228540 61712 228546
rect 61660 228482 61712 228488
rect 61304 219406 61424 219434
rect 61304 217977 61332 219406
rect 61672 218210 61700 228482
rect 62028 225208 62080 225214
rect 62028 225150 62080 225156
rect 61660 218204 61712 218210
rect 61660 218146 61712 218152
rect 62040 218074 62068 225150
rect 62304 219020 62356 219026
rect 62304 218962 62356 218968
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 62028 218068 62080 218074
rect 62028 218010 62080 218016
rect 61290 217968 61346 217977
rect 61290 217903 61346 217912
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217138 62344 218962
rect 62776 218890 62804 283183
rect 62946 282160 63002 282169
rect 62946 282095 63002 282104
rect 62960 225593 62988 282095
rect 63144 267073 63172 287127
rect 651484 287094 651512 287399
rect 651472 287088 651524 287094
rect 651472 287030 651524 287036
rect 651470 285968 651526 285977
rect 651470 285903 651526 285912
rect 651484 285734 651512 285903
rect 651472 285728 651524 285734
rect 651472 285670 651524 285676
rect 651470 284744 651526 284753
rect 651470 284679 651526 284688
rect 651484 284374 651512 284679
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 651760 282282 651788 288487
rect 652128 283529 652156 295287
rect 652390 291544 652446 291553
rect 652390 291479 652446 291488
rect 652114 283520 652170 283529
rect 652114 283455 652170 283464
rect 651760 282254 652156 282282
rect 651930 282160 651986 282169
rect 651930 282095 651986 282104
rect 651654 280936 651710 280945
rect 651654 280871 651710 280880
rect 651470 280392 651526 280401
rect 651470 280327 651472 280336
rect 651524 280327 651526 280336
rect 651472 280298 651524 280304
rect 651668 280226 651696 280871
rect 651656 280220 651708 280226
rect 651656 280162 651708 280168
rect 65904 273970 65932 278052
rect 67100 274378 67128 278052
rect 67088 274372 67140 274378
rect 67088 274314 67140 274320
rect 65892 273964 65944 273970
rect 65892 273906 65944 273912
rect 68204 271182 68232 278052
rect 69400 272678 69428 278052
rect 69388 272672 69440 272678
rect 69388 272614 69440 272620
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 70596 269958 70624 278052
rect 71792 275330 71820 278052
rect 71780 275324 71832 275330
rect 71780 275266 71832 275272
rect 72988 272542 73016 278052
rect 74184 274718 74212 278052
rect 74172 274712 74224 274718
rect 74172 274654 74224 274660
rect 72976 272536 73028 272542
rect 72976 272478 73028 272484
rect 75380 271318 75408 278052
rect 76484 275602 76512 278052
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 76748 274712 76800 274718
rect 76748 274654 76800 274660
rect 75368 271312 75420 271318
rect 75368 271254 75420 271260
rect 70584 269952 70636 269958
rect 70584 269894 70636 269900
rect 76760 269822 76788 274654
rect 77680 274106 77708 278052
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 76748 269816 76800 269822
rect 76748 269758 76800 269764
rect 78876 269550 78904 278052
rect 80072 277394 80100 278052
rect 80072 277366 80192 277394
rect 80164 269958 80192 277366
rect 81268 275466 81296 278052
rect 81256 275460 81308 275466
rect 81256 275402 81308 275408
rect 82464 272814 82492 278052
rect 83674 278038 84148 278066
rect 84778 278038 85528 278066
rect 82452 272808 82504 272814
rect 82452 272750 82504 272756
rect 79968 269952 80020 269958
rect 79968 269894 80020 269900
rect 80152 269952 80204 269958
rect 80152 269894 80204 269900
rect 78864 269544 78916 269550
rect 78864 269486 78916 269492
rect 79980 267170 80008 269894
rect 84120 269074 84148 278038
rect 85500 270094 85528 278038
rect 85960 274718 85988 278052
rect 86224 275596 86276 275602
rect 86224 275538 86276 275544
rect 85948 274712 86000 274718
rect 85948 274654 86000 274660
rect 85488 270088 85540 270094
rect 85488 270030 85540 270036
rect 84108 269068 84160 269074
rect 84108 269010 84160 269016
rect 86236 267442 86264 275538
rect 87156 271454 87184 278052
rect 87144 271448 87196 271454
rect 87144 271390 87196 271396
rect 88352 270366 88380 278052
rect 89456 278038 89562 278066
rect 89456 274242 89484 278038
rect 90744 275602 90772 278052
rect 91862 278038 92428 278066
rect 90732 275596 90784 275602
rect 90732 275538 90784 275544
rect 90364 274712 90416 274718
rect 90364 274654 90416 274660
rect 89444 274236 89496 274242
rect 89444 274178 89496 274184
rect 88340 270360 88392 270366
rect 88340 270302 88392 270308
rect 86224 267436 86276 267442
rect 86224 267378 86276 267384
rect 79968 267164 80020 267170
rect 79968 267106 80020 267112
rect 63130 267064 63186 267073
rect 90376 267034 90404 274654
rect 92400 268394 92428 278038
rect 93044 275738 93072 278052
rect 93032 275732 93084 275738
rect 93032 275674 93084 275680
rect 94240 271590 94268 278052
rect 95436 274378 95464 278052
rect 95884 274508 95936 274514
rect 95884 274450 95936 274456
rect 95424 274372 95476 274378
rect 95424 274314 95476 274320
rect 94228 271584 94280 271590
rect 94228 271526 94280 271532
rect 92388 268388 92440 268394
rect 92388 268330 92440 268336
rect 95896 267578 95924 274450
rect 96632 273834 96660 278052
rect 97842 278038 97948 278066
rect 96620 273828 96672 273834
rect 96620 273770 96672 273776
rect 97920 270230 97948 278038
rect 99024 272950 99052 278052
rect 100128 275874 100156 278052
rect 100116 275868 100168 275874
rect 100116 275810 100168 275816
rect 101324 273086 101352 278052
rect 101312 273080 101364 273086
rect 101312 273022 101364 273028
rect 99012 272944 99064 272950
rect 99012 272886 99064 272892
rect 97908 270224 97960 270230
rect 97908 270166 97960 270172
rect 102520 268530 102548 278052
rect 103716 274718 103744 278052
rect 104926 278038 105216 278066
rect 103704 274712 103756 274718
rect 103704 274654 103756 274660
rect 104808 274712 104860 274718
rect 104808 274654 104860 274660
rect 102508 268524 102560 268530
rect 102508 268466 102560 268472
rect 95884 267572 95936 267578
rect 95884 267514 95936 267520
rect 104820 267306 104848 274654
rect 105188 274514 105216 278038
rect 105176 274508 105228 274514
rect 105176 274450 105228 274456
rect 106108 271726 106136 278052
rect 107212 276010 107240 278052
rect 107200 276004 107252 276010
rect 107200 275946 107252 275952
rect 108408 271862 108436 278052
rect 109618 278038 110276 278066
rect 108396 271856 108448 271862
rect 108396 271798 108448 271804
rect 106096 271720 106148 271726
rect 106096 271662 106148 271668
rect 110248 268666 110276 278038
rect 110800 275058 110828 278052
rect 110788 275052 110840 275058
rect 110788 274994 110840 275000
rect 111996 268938 112024 278052
rect 113206 278038 113496 278066
rect 113468 274650 113496 278038
rect 113456 274644 113508 274650
rect 113456 274586 113508 274592
rect 114388 273222 114416 278052
rect 115506 278038 115888 278066
rect 114376 273216 114428 273222
rect 114376 273158 114428 273164
rect 111984 268932 112036 268938
rect 111984 268874 112036 268880
rect 115860 268802 115888 278038
rect 116688 271046 116716 278052
rect 117898 278038 118280 278066
rect 118252 273834 118280 278038
rect 117964 273828 118016 273834
rect 117964 273770 118016 273776
rect 118240 273828 118292 273834
rect 118240 273770 118292 273776
rect 116676 271040 116728 271046
rect 116676 270982 116728 270988
rect 115848 268796 115900 268802
rect 115848 268738 115900 268744
rect 110236 268660 110288 268666
rect 110236 268602 110288 268608
rect 117976 267714 118004 273770
rect 119080 272270 119108 278052
rect 120276 272406 120304 278052
rect 121486 278038 121684 278066
rect 120264 272400 120316 272406
rect 120264 272342 120316 272348
rect 119068 272264 119120 272270
rect 119068 272206 119120 272212
rect 121460 270360 121512 270366
rect 121460 270302 121512 270308
rect 117964 267708 118016 267714
rect 117964 267650 118016 267656
rect 104808 267300 104860 267306
rect 104808 267242 104860 267248
rect 63130 266999 63186 267008
rect 90364 267028 90416 267034
rect 90364 266970 90416 266976
rect 121472 266898 121500 270302
rect 121656 269278 121684 278038
rect 122576 270366 122604 278052
rect 123772 273698 123800 278052
rect 123760 273692 123812 273698
rect 123760 273634 123812 273640
rect 124968 270910 124996 278052
rect 126178 278038 126928 278066
rect 124956 270904 125008 270910
rect 124956 270846 125008 270852
rect 122564 270360 122616 270366
rect 122564 270302 122616 270308
rect 126900 269686 126928 278038
rect 127360 270774 127388 278052
rect 127348 270768 127400 270774
rect 127348 270710 127400 270716
rect 126888 269680 126940 269686
rect 126888 269622 126940 269628
rect 121644 269272 121696 269278
rect 121644 269214 121696 269220
rect 128556 268258 128584 278052
rect 129476 278038 129674 278066
rect 129476 270502 129504 278038
rect 130856 272134 130884 278052
rect 132052 274922 132080 278052
rect 133262 278038 133828 278066
rect 132040 274916 132092 274922
rect 132040 274858 132092 274864
rect 130844 272128 130896 272134
rect 130844 272070 130896 272076
rect 129464 270496 129516 270502
rect 129464 270438 129516 270444
rect 133800 269550 133828 278038
rect 134444 273562 134472 278052
rect 134432 273556 134484 273562
rect 134432 273498 134484 273504
rect 135640 273426 135668 278052
rect 136836 274786 136864 278052
rect 136824 274780 136876 274786
rect 136824 274722 136876 274728
rect 137652 274780 137704 274786
rect 137652 274722 137704 274728
rect 136824 273964 136876 273970
rect 136824 273906 136876 273912
rect 135628 273420 135680 273426
rect 135628 273362 135680 273368
rect 130384 269544 130436 269550
rect 130384 269486 130436 269492
rect 133788 269544 133840 269550
rect 133788 269486 133840 269492
rect 128544 268252 128596 268258
rect 128544 268194 128596 268200
rect 121460 266892 121512 266898
rect 121460 266834 121512 266840
rect 130396 266762 130424 269486
rect 130384 266756 130436 266762
rect 130384 266698 130436 266704
rect 136836 264330 136864 273906
rect 137664 269074 137692 274722
rect 137940 270638 137968 278052
rect 139136 275194 139164 278052
rect 140346 278038 140728 278066
rect 139124 275188 139176 275194
rect 139124 275130 139176 275136
rect 139400 272672 139452 272678
rect 139400 272614 139452 272620
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137928 270632 137980 270638
rect 137928 270574 137980 270580
rect 137468 269068 137520 269074
rect 137468 269010 137520 269016
rect 137652 269068 137704 269074
rect 137652 269010 137704 269016
rect 137480 266626 137508 269010
rect 138112 267572 138164 267578
rect 138112 267514 138164 267520
rect 137468 266620 137520 266626
rect 137468 266562 137520 266568
rect 136836 264302 137310 264330
rect 138124 264316 138152 267514
rect 138492 264330 138520 271118
rect 139412 264330 139440 272614
rect 140700 269414 140728 278038
rect 141056 275324 141108 275330
rect 141056 275266 141108 275272
rect 140688 269408 140740 269414
rect 140688 269350 140740 269356
rect 140596 267164 140648 267170
rect 140596 267106 140648 267112
rect 138492 264302 138966 264330
rect 139412 264302 139794 264330
rect 140608 264316 140636 267106
rect 141068 264330 141096 275266
rect 141528 272678 141556 278052
rect 141516 272672 141568 272678
rect 141516 272614 141568 272620
rect 142160 272536 142212 272542
rect 142160 272478 142212 272484
rect 142172 264330 142200 272478
rect 142724 271318 142752 278052
rect 143920 274786 143948 278052
rect 143908 274780 143960 274786
rect 143908 274722 143960 274728
rect 144368 274780 144420 274786
rect 144368 274722 144420 274728
rect 142712 271312 142764 271318
rect 142712 271254 142764 271260
rect 144184 271312 144236 271318
rect 144184 271254 144236 271260
rect 142712 271176 142764 271182
rect 142712 271118 142764 271124
rect 142724 264330 142752 271118
rect 143908 269816 143960 269822
rect 143908 269758 143960 269764
rect 141068 264302 141450 264330
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143920 264316 143948 269758
rect 144196 267170 144224 271254
rect 144380 269822 144408 274722
rect 144920 274100 144972 274106
rect 144920 274042 144972 274048
rect 144368 269816 144420 269822
rect 144368 269758 144420 269764
rect 144932 267734 144960 274042
rect 145116 273970 145144 278052
rect 145564 275460 145616 275466
rect 145564 275402 145616 275408
rect 145104 273964 145156 273970
rect 145104 273906 145156 273912
rect 144932 267706 145144 267734
rect 144736 267436 144788 267442
rect 144736 267378 144788 267384
rect 144184 267164 144236 267170
rect 144184 267106 144236 267112
rect 144748 264316 144776 267378
rect 144920 266892 144972 266898
rect 144920 266834 144972 266840
rect 144932 266490 144960 266834
rect 144920 266484 144972 266490
rect 144920 266426 144972 266432
rect 145116 264330 145144 267706
rect 145380 266892 145432 266898
rect 145380 266834 145432 266840
rect 145392 266626 145420 266834
rect 145576 266626 145604 275402
rect 146220 275330 146248 278052
rect 146208 275324 146260 275330
rect 146208 275266 146260 275272
rect 146944 275188 146996 275194
rect 146944 275130 146996 275136
rect 146956 274786 146984 275130
rect 146944 274780 146996 274786
rect 146944 274722 146996 274728
rect 147416 274106 147444 278052
rect 147404 274100 147456 274106
rect 147404 274042 147456 274048
rect 146944 273420 146996 273426
rect 146944 273362 146996 273368
rect 146392 269952 146444 269958
rect 146392 269894 146444 269900
rect 145380 266620 145432 266626
rect 145380 266562 145432 266568
rect 145564 266620 145616 266626
rect 145564 266562 145616 266568
rect 145116 264302 145590 264330
rect 146404 264316 146432 269894
rect 146956 267442 146984 273362
rect 148416 272808 148468 272814
rect 148416 272750 148468 272756
rect 146944 267436 146996 267442
rect 146944 267378 146996 267384
rect 147220 266756 147272 266762
rect 147220 266698 147272 266704
rect 147232 264316 147260 266698
rect 148048 266620 148100 266626
rect 148048 266562 148100 266568
rect 148060 264316 148088 266562
rect 148428 264330 148456 272750
rect 148612 271182 148640 278052
rect 149808 275194 149836 278052
rect 151018 278038 151768 278066
rect 149796 275188 149848 275194
rect 149796 275130 149848 275136
rect 149704 275052 149756 275058
rect 149704 274994 149756 275000
rect 148600 271176 148652 271182
rect 148600 271118 148652 271124
rect 149428 270088 149480 270094
rect 149428 270030 149480 270036
rect 149440 264330 149468 270030
rect 149716 266762 149744 274994
rect 151740 268258 151768 278038
rect 152004 274236 152056 274242
rect 152004 274178 152056 274184
rect 150440 268252 150492 268258
rect 150440 268194 150492 268200
rect 151728 268252 151780 268258
rect 151728 268194 151780 268200
rect 150452 267578 150480 268194
rect 150440 267572 150492 267578
rect 150440 267514 150492 267520
rect 151360 267028 151412 267034
rect 151360 266970 151412 266976
rect 150532 266892 150584 266898
rect 150532 266834 150584 266840
rect 149704 266756 149756 266762
rect 149704 266698 149756 266704
rect 148428 264302 148902 264330
rect 149440 264302 149730 264330
rect 150544 264316 150572 266834
rect 151372 264316 151400 266970
rect 152016 265674 152044 274178
rect 152200 272542 152228 278052
rect 153396 275058 153424 278052
rect 154316 278038 154514 278066
rect 153384 275052 153436 275058
rect 153384 274994 153436 275000
rect 152188 272536 152240 272542
rect 152188 272478 152240 272484
rect 152188 271448 152240 271454
rect 152188 271390 152240 271396
rect 152004 265668 152056 265674
rect 152004 265610 152056 265616
rect 152200 264316 152228 271390
rect 154316 271318 154344 278038
rect 154764 275596 154816 275602
rect 154764 275538 154816 275544
rect 154488 275052 154540 275058
rect 154488 274994 154540 275000
rect 154304 271312 154356 271318
rect 154304 271254 154356 271260
rect 154500 267034 154528 274994
rect 154776 267734 154804 275538
rect 155696 274242 155724 278052
rect 155960 275732 156012 275738
rect 155960 275674 156012 275680
rect 155684 274236 155736 274242
rect 155684 274178 155736 274184
rect 155500 268388 155552 268394
rect 155500 268330 155552 268336
rect 154684 267706 154804 267734
rect 154488 267028 154540 267034
rect 154488 266970 154540 266976
rect 153844 266484 153896 266490
rect 153844 266426 153896 266432
rect 152740 265668 152792 265674
rect 152740 265610 152792 265616
rect 152752 264330 152780 265610
rect 152752 264302 153042 264330
rect 153856 264316 153884 266426
rect 154684 264316 154712 267706
rect 155512 264316 155540 268330
rect 155972 265674 156000 275674
rect 156892 275602 156920 278052
rect 156880 275596 156932 275602
rect 156880 275538 156932 275544
rect 157616 274372 157668 274378
rect 157616 274314 157668 274320
rect 156144 271584 156196 271590
rect 156144 271526 156196 271532
rect 155960 265668 156012 265674
rect 155960 265610 156012 265616
rect 156156 264330 156184 271526
rect 156788 265668 156840 265674
rect 156788 265610 156840 265616
rect 156800 264330 156828 265610
rect 157628 264330 157656 274314
rect 158088 272814 158116 278052
rect 158076 272808 158128 272814
rect 158076 272750 158128 272756
rect 159284 271454 159312 278052
rect 160480 275466 160508 278052
rect 161584 275874 161612 278052
rect 162124 276004 162176 276010
rect 162124 275946 162176 275952
rect 161388 275868 161440 275874
rect 161388 275810 161440 275816
rect 161572 275868 161624 275874
rect 161572 275810 161624 275816
rect 161756 275868 161808 275874
rect 161756 275810 161808 275816
rect 160468 275460 160520 275466
rect 160468 275402 160520 275408
rect 161400 273170 161428 275810
rect 161768 275754 161796 275810
rect 161676 275726 161796 275754
rect 161676 275058 161704 275726
rect 161848 275460 161900 275466
rect 161848 275402 161900 275408
rect 161860 275058 161888 275402
rect 161664 275052 161716 275058
rect 161664 274994 161716 275000
rect 161848 275052 161900 275058
rect 161848 274994 161900 275000
rect 161400 273142 161612 273170
rect 160928 273080 160980 273086
rect 160928 273022 160980 273028
rect 160100 272944 160152 272950
rect 160100 272886 160152 272892
rect 159272 271448 159324 271454
rect 159272 271390 159324 271396
rect 158812 270224 158864 270230
rect 158812 270166 158864 270172
rect 156156 264302 156354 264330
rect 156800 264302 157182 264330
rect 157628 264302 158010 264330
rect 158824 264316 158852 270166
rect 159640 267708 159692 267714
rect 159640 267650 159692 267656
rect 159652 264316 159680 267650
rect 160112 264330 160140 272886
rect 160940 264330 160968 273022
rect 161584 267734 161612 273142
rect 161584 267706 161704 267734
rect 161676 264330 161704 267706
rect 162136 266422 162164 275946
rect 162780 272950 162808 278052
rect 163976 277394 164004 278052
rect 165186 278038 165476 278066
rect 163976 277366 164096 277394
rect 164068 275738 164096 277366
rect 163136 275732 163188 275738
rect 163136 275674 163188 275680
rect 164056 275732 164108 275738
rect 164056 275674 164108 275680
rect 162768 272944 162820 272950
rect 162768 272886 162820 272892
rect 162952 268524 163004 268530
rect 162952 268466 163004 268472
rect 162124 266416 162176 266422
rect 162124 266358 162176 266364
rect 160112 264302 160494 264330
rect 160940 264302 161322 264330
rect 161676 264302 162150 264330
rect 162964 264316 162992 268466
rect 163148 268122 163176 275674
rect 163320 274508 163372 274514
rect 163320 274450 163372 274456
rect 163136 268116 163188 268122
rect 163136 268058 163188 268064
rect 163332 264330 163360 274450
rect 164976 271720 165028 271726
rect 164976 271662 165028 271668
rect 164608 267300 164660 267306
rect 164608 267242 164660 267248
rect 163332 264302 163806 264330
rect 164620 264316 164648 267242
rect 164988 264330 165016 271662
rect 165448 269958 165476 278038
rect 166368 274378 166396 278052
rect 167000 275868 167052 275874
rect 167000 275810 167052 275816
rect 166356 274372 166408 274378
rect 166356 274314 166408 274320
rect 165896 271856 165948 271862
rect 165896 271798 165948 271804
rect 165436 269952 165488 269958
rect 165436 269894 165488 269900
rect 165908 264330 165936 271798
rect 167012 268666 167040 275810
rect 167564 274922 167592 278052
rect 167552 274916 167604 274922
rect 167552 274858 167604 274864
rect 168760 274514 168788 278052
rect 169878 278038 170168 278066
rect 169024 274916 169076 274922
rect 169024 274858 169076 274864
rect 168748 274508 168800 274514
rect 168748 274450 168800 274456
rect 167828 269272 167880 269278
rect 167828 269214 167880 269220
rect 167000 268660 167052 268666
rect 167000 268602 167052 268608
rect 167644 268388 167696 268394
rect 167644 268330 167696 268336
rect 167092 266416 167144 266422
rect 167092 266358 167144 266364
rect 164988 264302 165462 264330
rect 165908 264302 166290 264330
rect 167104 264316 167132 266358
rect 167656 264330 167684 268330
rect 167840 267714 167868 269214
rect 168748 268932 168800 268938
rect 168748 268874 168800 268880
rect 168012 268388 168064 268394
rect 168012 268330 168064 268336
rect 168024 268122 168052 268330
rect 168012 268116 168064 268122
rect 168012 268058 168064 268064
rect 167828 267708 167880 267714
rect 167828 267650 167880 267656
rect 167656 264302 167946 264330
rect 168760 264316 168788 268874
rect 169036 267306 169064 274858
rect 169944 274644 169996 274650
rect 169944 274586 169996 274592
rect 169024 267300 169076 267306
rect 169024 267242 169076 267248
rect 169576 266756 169628 266762
rect 169576 266698 169628 266704
rect 169588 264316 169616 266698
rect 169956 264330 169984 274586
rect 170140 271590 170168 278038
rect 171060 275738 171088 278052
rect 171048 275732 171100 275738
rect 171048 275674 171100 275680
rect 171600 273216 171652 273222
rect 171600 273158 171652 273164
rect 170128 271584 170180 271590
rect 170128 271526 170180 271532
rect 171232 268524 171284 268530
rect 171232 268466 171284 268472
rect 169956 264302 170430 264330
rect 171244 264316 171272 268466
rect 171612 264330 171640 273158
rect 172256 273086 172284 278052
rect 173466 278038 173756 278066
rect 172244 273080 172296 273086
rect 172244 273022 172296 273028
rect 172520 272264 172572 272270
rect 172520 272206 172572 272212
rect 172532 265674 172560 272206
rect 172704 271040 172756 271046
rect 172704 270982 172756 270988
rect 172520 265668 172572 265674
rect 172520 265610 172572 265616
rect 172716 264330 172744 270982
rect 173728 270094 173756 278038
rect 174648 274854 174676 278052
rect 174636 274848 174688 274854
rect 174636 274790 174688 274796
rect 174452 274780 174504 274786
rect 174452 274722 174504 274728
rect 174176 273828 174228 273834
rect 174176 273770 174228 273776
rect 173716 270088 173768 270094
rect 173716 270030 173768 270036
rect 173348 265668 173400 265674
rect 173348 265610 173400 265616
rect 173360 264330 173388 265610
rect 174188 264330 174216 273770
rect 174464 272270 174492 274722
rect 175280 272400 175332 272406
rect 175280 272342 175332 272348
rect 174452 272264 174504 272270
rect 174452 272206 174504 272212
rect 175292 264330 175320 272342
rect 175752 271726 175780 278052
rect 175924 275052 175976 275058
rect 175924 274994 175976 275000
rect 175936 273834 175964 274994
rect 175924 273828 175976 273834
rect 175924 273770 175976 273776
rect 175740 271720 175792 271726
rect 175740 271662 175792 271668
rect 176200 270360 176252 270366
rect 176200 270302 176252 270308
rect 171612 264302 172086 264330
rect 172716 264302 172914 264330
rect 173360 264302 173742 264330
rect 174188 264302 174570 264330
rect 175292 264302 175398 264330
rect 176212 264316 176240 270302
rect 176948 268530 176976 278052
rect 178144 275874 178172 278052
rect 178132 275868 178184 275874
rect 178132 275810 178184 275816
rect 177488 273692 177540 273698
rect 177488 273634 177540 273640
rect 176936 268524 176988 268530
rect 176936 268466 176988 268472
rect 177028 267708 177080 267714
rect 177028 267650 177080 267656
rect 177040 264316 177068 267650
rect 177500 264330 177528 273634
rect 178684 270904 178736 270910
rect 178684 270846 178736 270852
rect 178316 269680 178368 269686
rect 178316 269622 178368 269628
rect 178328 264330 178356 269622
rect 178696 266422 178724 270846
rect 179340 270230 179368 278052
rect 180550 278038 180748 278066
rect 181746 278038 182036 278066
rect 179880 270768 179932 270774
rect 179880 270710 179932 270716
rect 179328 270224 179380 270230
rect 179328 270166 179380 270172
rect 178684 266416 178736 266422
rect 178684 266358 178736 266364
rect 179512 266416 179564 266422
rect 179512 266358 179564 266364
rect 177500 264302 177882 264330
rect 178328 264302 178710 264330
rect 179524 264316 179552 266358
rect 179892 264330 179920 270710
rect 180720 270366 180748 278038
rect 181168 270496 181220 270502
rect 181168 270438 181220 270444
rect 180708 270360 180760 270366
rect 180708 270302 180760 270308
rect 179892 264302 180366 264330
rect 181180 264316 181208 270438
rect 182008 267714 182036 278038
rect 182732 274848 182784 274854
rect 182732 274790 182784 274796
rect 182456 272128 182508 272134
rect 182456 272070 182508 272076
rect 181996 267708 182048 267714
rect 181996 267650 182048 267656
rect 181996 267572 182048 267578
rect 181996 267514 182048 267520
rect 182008 264316 182036 267514
rect 182468 264330 182496 272070
rect 182744 267714 182772 274790
rect 182928 274650 182956 278052
rect 182916 274644 182968 274650
rect 182916 274586 182968 274592
rect 184124 273222 184152 278052
rect 185228 276010 185256 278052
rect 185216 276004 185268 276010
rect 185216 275946 185268 275952
rect 185124 273556 185176 273562
rect 185124 273498 185176 273504
rect 184112 273216 184164 273222
rect 184112 273158 184164 273164
rect 184940 272672 184992 272678
rect 184940 272614 184992 272620
rect 184952 272406 184980 272614
rect 184940 272400 184992 272406
rect 184940 272342 184992 272348
rect 183652 269544 183704 269550
rect 183652 269486 183704 269492
rect 182732 267708 182784 267714
rect 182732 267650 182784 267656
rect 182468 264302 182850 264330
rect 183664 264316 183692 269486
rect 184480 268660 184532 268666
rect 184480 268602 184532 268608
rect 184492 264316 184520 268602
rect 185136 264330 185164 273498
rect 186424 269550 186452 278052
rect 187344 278038 187634 278066
rect 186412 269544 186464 269550
rect 186412 269486 186464 269492
rect 186136 269068 186188 269074
rect 186136 269010 186188 269016
rect 185136 264302 185334 264330
rect 186148 264316 186176 269010
rect 187344 268666 187372 278038
rect 188816 271862 188844 278052
rect 189080 275324 189132 275330
rect 189080 275266 189132 275272
rect 189092 272678 189120 275266
rect 190012 275058 190040 278052
rect 191222 278038 191512 278066
rect 192418 278038 192800 278066
rect 193522 278038 193628 278066
rect 190000 275052 190052 275058
rect 190000 274994 190052 275000
rect 189080 272672 189132 272678
rect 189080 272614 189132 272620
rect 189172 272400 189224 272406
rect 189172 272342 189224 272348
rect 188804 271856 188856 271862
rect 188804 271798 188856 271804
rect 187700 270632 187752 270638
rect 187700 270574 187752 270580
rect 187332 268660 187384 268666
rect 187332 268602 187384 268608
rect 186964 267436 187016 267442
rect 186964 267378 187016 267384
rect 186976 264316 187004 267378
rect 187712 264330 187740 270574
rect 188620 269408 188672 269414
rect 188620 269350 188672 269356
rect 187712 264302 187818 264330
rect 188632 264316 188660 269350
rect 189184 265674 189212 272342
rect 189356 272264 189408 272270
rect 189356 272206 189408 272212
rect 189172 265668 189224 265674
rect 189172 265610 189224 265616
rect 189368 264330 189396 272206
rect 191484 271998 191512 278038
rect 191748 275188 191800 275194
rect 191748 275130 191800 275136
rect 191472 271992 191524 271998
rect 191472 271934 191524 271940
rect 191760 270502 191788 275130
rect 192392 273964 192444 273970
rect 192392 273906 192444 273912
rect 191748 270496 191800 270502
rect 191748 270438 191800 270444
rect 190828 269816 190880 269822
rect 190828 269758 190880 269764
rect 189908 265668 189960 265674
rect 189908 265610 189960 265616
rect 189920 264330 189948 265610
rect 190840 264330 190868 269758
rect 191932 267164 191984 267170
rect 191932 267106 191984 267112
rect 189368 264302 189474 264330
rect 189920 264302 190302 264330
rect 190840 264302 191130 264330
rect 191944 264316 191972 267106
rect 192404 264330 192432 273906
rect 192576 271856 192628 271862
rect 192576 271798 192628 271804
rect 192588 267170 192616 271798
rect 192772 271046 192800 278038
rect 193404 274100 193456 274106
rect 193404 274042 193456 274048
rect 192760 271040 192812 271046
rect 192760 270982 192812 270988
rect 192576 267164 192628 267170
rect 192576 267106 192628 267112
rect 193416 264330 193444 274042
rect 193600 272406 193628 278038
rect 194704 272678 194732 278052
rect 195900 273970 195928 278052
rect 195888 273964 195940 273970
rect 195888 273906 195940 273912
rect 194048 272672 194100 272678
rect 194048 272614 194100 272620
rect 194692 272672 194744 272678
rect 194692 272614 194744 272620
rect 193588 272400 193640 272406
rect 193588 272342 193640 272348
rect 194060 264330 194088 272614
rect 197096 271182 197124 278052
rect 198292 274106 198320 278052
rect 198740 275460 198792 275466
rect 198740 275402 198792 275408
rect 198280 274100 198332 274106
rect 198280 274042 198332 274048
rect 197544 272536 197596 272542
rect 197544 272478 197596 272484
rect 194784 271176 194836 271182
rect 194784 271118 194836 271124
rect 197084 271176 197136 271182
rect 197084 271118 197136 271124
rect 194796 264330 194824 271118
rect 196900 270496 196952 270502
rect 196900 270438 196952 270444
rect 196072 268252 196124 268258
rect 196072 268194 196124 268200
rect 192404 264302 192786 264330
rect 193416 264302 193614 264330
rect 194060 264302 194442 264330
rect 194796 264302 195270 264330
rect 196084 264316 196112 268194
rect 196912 264316 196940 270438
rect 197556 264330 197584 272478
rect 198096 271312 198148 271318
rect 198096 271254 198148 271260
rect 198108 264330 198136 271254
rect 198752 267850 198780 275402
rect 199488 272542 199516 278052
rect 200592 277394 200620 278052
rect 200500 277366 200620 277394
rect 200120 274236 200172 274242
rect 200120 274178 200172 274184
rect 199476 272536 199528 272542
rect 199476 272478 199528 272484
rect 198740 267844 198792 267850
rect 198740 267786 198792 267792
rect 199384 267028 199436 267034
rect 199384 266970 199436 266976
rect 197556 264302 197754 264330
rect 198108 264302 198582 264330
rect 199396 264316 199424 266970
rect 200132 264330 200160 274178
rect 200500 269686 200528 277366
rect 200672 272808 200724 272814
rect 200672 272750 200724 272756
rect 200488 269680 200540 269686
rect 200488 269622 200540 269628
rect 200684 264330 200712 272750
rect 201788 270502 201816 278052
rect 202328 271448 202380 271454
rect 202328 271390 202380 271396
rect 201776 270496 201828 270502
rect 201776 270438 201828 270444
rect 201868 267844 201920 267850
rect 201868 267786 201920 267792
rect 200132 264302 200238 264330
rect 200684 264302 201066 264330
rect 201880 264316 201908 267786
rect 202340 264330 202368 271390
rect 202984 269822 203012 278052
rect 203904 278038 204194 278066
rect 202972 269816 203024 269822
rect 202972 269758 203024 269764
rect 203904 268394 203932 278038
rect 205376 274242 205404 278052
rect 206376 275596 206428 275602
rect 206376 275538 206428 275544
rect 205364 274236 205416 274242
rect 205364 274178 205416 274184
rect 204260 273828 204312 273834
rect 204260 273770 204312 273776
rect 204076 269544 204128 269550
rect 204076 269486 204128 269492
rect 203524 268388 203576 268394
rect 203524 268330 203576 268336
rect 203892 268388 203944 268394
rect 203892 268330 203944 268336
rect 202340 264302 202722 264330
rect 203536 264316 203564 268330
rect 204088 266898 204116 269486
rect 204076 266892 204128 266898
rect 204076 266834 204128 266840
rect 204272 264330 204300 273770
rect 204720 272944 204772 272950
rect 204720 272886 204772 272892
rect 204732 264330 204760 272886
rect 206008 269952 206060 269958
rect 206008 269894 206060 269900
rect 204272 264302 204378 264330
rect 204732 264302 205206 264330
rect 206020 264316 206048 269894
rect 206388 264330 206416 275538
rect 206572 273834 206600 278052
rect 207768 274378 207796 278052
rect 208492 274508 208544 274514
rect 208492 274450 208544 274456
rect 207296 274372 207348 274378
rect 207296 274314 207348 274320
rect 207756 274372 207808 274378
rect 207756 274314 207808 274320
rect 206560 273828 206612 273834
rect 206560 273770 206612 273776
rect 207308 264330 207336 274314
rect 206388 264302 206862 264330
rect 207308 264302 207690 264330
rect 208504 264316 208532 274450
rect 208872 272814 208900 278052
rect 208860 272808 208912 272814
rect 208860 272750 208912 272756
rect 209780 271584 209832 271590
rect 209780 271526 209832 271532
rect 209320 267300 209372 267306
rect 209320 267242 209372 267248
rect 209332 264316 209360 267242
rect 209792 264330 209820 271526
rect 210068 269958 210096 278052
rect 211264 277394 211292 278052
rect 212276 278038 212474 278066
rect 211264 277366 211384 277394
rect 211068 275732 211120 275738
rect 211068 275674 211120 275680
rect 210608 273080 210660 273086
rect 210608 273022 210660 273028
rect 210056 269952 210108 269958
rect 210056 269894 210108 269900
rect 210620 264330 210648 273022
rect 211080 271810 211108 275674
rect 211080 271782 211200 271810
rect 211172 267734 211200 271782
rect 211356 268802 211384 277366
rect 212276 271318 212304 278038
rect 213000 271720 213052 271726
rect 213000 271662 213052 271668
rect 212264 271312 212316 271318
rect 212264 271254 212316 271260
rect 212632 270088 212684 270094
rect 212632 270030 212684 270036
rect 211344 268796 211396 268802
rect 211344 268738 211396 268744
rect 211172 267706 211384 267734
rect 211356 264330 211384 267706
rect 209792 264302 210174 264330
rect 210620 264302 211002 264330
rect 211356 264302 211830 264330
rect 212644 264316 212672 270030
rect 213012 264330 213040 271662
rect 213656 271454 213684 278052
rect 214852 275466 214880 278052
rect 215970 278038 216536 278066
rect 214840 275460 214892 275466
rect 214840 275402 214892 275408
rect 214564 274644 214616 274650
rect 214564 274586 214616 274592
rect 213644 271448 213696 271454
rect 213644 271390 213696 271396
rect 214104 270224 214156 270230
rect 214104 270166 214156 270172
rect 214116 266558 214144 270166
rect 214288 267708 214340 267714
rect 214288 267650 214340 267656
rect 214104 266552 214156 266558
rect 214104 266494 214156 266500
rect 213012 264302 213486 264330
rect 214300 264316 214328 267650
rect 214576 266694 214604 274586
rect 215300 270360 215352 270366
rect 215300 270302 215352 270308
rect 215116 268524 215168 268530
rect 215116 268466 215168 268472
rect 214564 266688 214616 266694
rect 214564 266630 214616 266636
rect 215128 264316 215156 268466
rect 215312 266422 215340 270302
rect 216508 270094 216536 278038
rect 217152 275874 217180 278052
rect 216680 275868 216732 275874
rect 216680 275810 216732 275816
rect 217140 275868 217192 275874
rect 217140 275810 217192 275816
rect 216496 270088 216548 270094
rect 216496 270030 216548 270036
rect 215944 266552 215996 266558
rect 215944 266494 215996 266500
rect 215300 266416 215352 266422
rect 215300 266358 215352 266364
rect 215956 264316 215984 266494
rect 216692 264330 216720 275810
rect 218348 275330 218376 278052
rect 218336 275324 218388 275330
rect 218336 275266 218388 275272
rect 218704 275052 218756 275058
rect 218704 274994 218756 275000
rect 218716 267306 218744 274994
rect 218888 273216 218940 273222
rect 218888 273158 218940 273164
rect 218704 267300 218756 267306
rect 218704 267242 218756 267248
rect 218900 267034 218928 273158
rect 219544 272950 219572 278052
rect 220464 278038 220754 278066
rect 219532 272944 219584 272950
rect 219532 272886 219584 272892
rect 219440 268660 219492 268666
rect 219440 268602 219492 268608
rect 219256 267572 219308 267578
rect 219256 267514 219308 267520
rect 218888 267028 218940 267034
rect 218888 266970 218940 266976
rect 218428 266688 218480 266694
rect 218428 266630 218480 266636
rect 217600 266416 217652 266422
rect 217600 266358 217652 266364
rect 216692 264302 216798 264330
rect 217612 264316 217640 266358
rect 218440 264316 218468 266630
rect 219268 264316 219296 267514
rect 219452 266422 219480 268602
rect 220464 268530 220492 278038
rect 221280 276004 221332 276010
rect 221280 275946 221332 275952
rect 220452 268524 220504 268530
rect 220452 268466 220504 268472
rect 220084 267028 220136 267034
rect 220084 266970 220136 266976
rect 219440 266416 219492 266422
rect 219440 266358 219492 266364
rect 220096 264316 220124 266970
rect 220912 266892 220964 266898
rect 220912 266834 220964 266840
rect 220924 264316 220952 266834
rect 221292 264330 221320 275946
rect 221936 275602 221964 278052
rect 221924 275596 221976 275602
rect 221924 275538 221976 275544
rect 223132 271590 223160 278052
rect 224040 275868 224092 275874
rect 224040 275810 224092 275816
rect 224052 273086 224080 275810
rect 224236 275738 224264 278052
rect 224224 275732 224276 275738
rect 224224 275674 224276 275680
rect 224040 273080 224092 273086
rect 224040 273022 224092 273028
rect 224224 272400 224276 272406
rect 224224 272342 224276 272348
rect 223120 271584 223172 271590
rect 223120 271526 223172 271532
rect 223488 268796 223540 268802
rect 223488 268738 223540 268744
rect 223500 267306 223528 268738
rect 223028 267300 223080 267306
rect 223028 267242 223080 267248
rect 223488 267300 223540 267306
rect 223488 267242 223540 267248
rect 222568 266416 222620 266422
rect 222568 266358 222620 266364
rect 221292 264302 221766 264330
rect 222580 264316 222608 266358
rect 223040 264330 223068 267242
rect 223948 267164 224000 267170
rect 223948 267106 224000 267112
rect 223960 264330 223988 267106
rect 224236 266422 224264 272342
rect 225432 271862 225460 278052
rect 225052 271856 225104 271862
rect 225052 271798 225104 271804
rect 225420 271856 225472 271862
rect 225420 271798 225472 271804
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 223040 264302 223422 264330
rect 223960 264302 224250 264330
rect 225064 264316 225092 271798
rect 225512 271040 225564 271046
rect 225512 270982 225564 270988
rect 225524 264330 225552 270982
rect 226628 270230 226656 278052
rect 227824 274514 227852 278052
rect 227812 274508 227864 274514
rect 227812 274450 227864 274456
rect 229020 273970 229048 278052
rect 229192 274100 229244 274106
rect 229192 274042 229244 274048
rect 227904 273964 227956 273970
rect 227904 273906 227956 273912
rect 229008 273964 229060 273970
rect 229008 273906 229060 273912
rect 227168 272672 227220 272678
rect 227168 272614 227220 272620
rect 226616 270224 226668 270230
rect 226616 270166 226668 270172
rect 226892 269680 226944 269686
rect 226892 269622 226944 269628
rect 226904 266626 226932 269622
rect 226892 266620 226944 266626
rect 226892 266562 226944 266568
rect 226708 266416 226760 266422
rect 226708 266358 226760 266364
rect 225524 264302 225906 264330
rect 226720 264316 226748 266358
rect 227180 264330 227208 272614
rect 227916 264330 227944 273906
rect 229204 273850 229232 274042
rect 229112 273822 229232 273850
rect 228364 271856 228416 271862
rect 228364 271798 228416 271804
rect 228376 267034 228404 271798
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 229112 265674 229140 273822
rect 230216 271182 230244 278052
rect 231334 278038 231716 278066
rect 230572 272536 230624 272542
rect 230572 272478 230624 272484
rect 229284 271176 229336 271182
rect 229284 271118 229336 271124
rect 230204 271176 230256 271182
rect 230204 271118 230256 271124
rect 229100 265668 229152 265674
rect 229100 265610 229152 265616
rect 229296 265554 229324 271118
rect 229652 265668 229704 265674
rect 229652 265610 229704 265616
rect 229204 265526 229324 265554
rect 227180 264302 227562 264330
rect 227916 264302 228390 264330
rect 229204 264316 229232 265526
rect 229664 264330 229692 265610
rect 230584 264330 230612 272478
rect 231688 268394 231716 278038
rect 232516 275874 232544 278052
rect 232504 275868 232556 275874
rect 232504 275810 232556 275816
rect 232780 275732 232832 275738
rect 232780 275674 232832 275680
rect 232228 270496 232280 270502
rect 232228 270438 232280 270444
rect 230756 268388 230808 268394
rect 230756 268330 230808 268336
rect 231676 268388 231728 268394
rect 231676 268330 231728 268336
rect 230768 266762 230796 268330
rect 230756 266756 230808 266762
rect 230756 266698 230808 266704
rect 231676 266620 231728 266626
rect 231676 266562 231728 266568
rect 229664 264302 230046 264330
rect 230584 264302 230874 264330
rect 231688 264316 231716 266562
rect 232240 264330 232268 270438
rect 232792 270366 232820 275674
rect 233712 272542 233740 278052
rect 233884 274372 233936 274378
rect 233884 274314 233936 274320
rect 233700 272536 233752 272542
rect 233700 272478 233752 272484
rect 232780 270360 232832 270366
rect 232780 270302 232832 270308
rect 233332 269816 233384 269822
rect 233332 269758 233384 269764
rect 232240 264302 232530 264330
rect 233344 264316 233372 269758
rect 233896 266422 233924 274314
rect 234908 274242 234936 278052
rect 236104 275738 236132 278052
rect 236092 275732 236144 275738
rect 236092 275674 236144 275680
rect 236644 275460 236696 275466
rect 236644 275402 236696 275408
rect 234712 274236 234764 274242
rect 234712 274178 234764 274184
rect 234896 274236 234948 274242
rect 234896 274178 234948 274184
rect 234160 266756 234212 266762
rect 234160 266698 234212 266704
rect 233884 266416 233936 266422
rect 233884 266358 233936 266364
rect 234172 264316 234200 266698
rect 234724 264330 234752 274178
rect 235448 273828 235500 273834
rect 235448 273770 235500 273776
rect 235460 264330 235488 273770
rect 236656 267442 236684 275402
rect 237300 274106 237328 278052
rect 237288 274100 237340 274106
rect 237288 274042 237340 274048
rect 237380 272808 237432 272814
rect 237380 272750 237432 272756
rect 236644 267436 236696 267442
rect 236644 267378 236696 267384
rect 236644 266416 236696 266422
rect 236644 266358 236696 266364
rect 234724 264302 235014 264330
rect 235460 264302 235842 264330
rect 236656 264316 236684 266358
rect 237392 264330 237420 272750
rect 238496 272678 238524 278052
rect 239404 275596 239456 275602
rect 239404 275538 239456 275544
rect 239416 275346 239444 275538
rect 239600 275466 239628 278052
rect 240810 278038 241468 278066
rect 239864 275868 239916 275874
rect 239864 275810 239916 275816
rect 239588 275460 239640 275466
rect 239588 275402 239640 275408
rect 239416 275318 239536 275346
rect 238484 272672 238536 272678
rect 238484 272614 238536 272620
rect 239312 271312 239364 271318
rect 239312 271254 239364 271260
rect 238300 269952 238352 269958
rect 238300 269894 238352 269900
rect 237392 264302 237498 264330
rect 238312 264316 238340 269894
rect 239324 267734 239352 271254
rect 239508 267734 239536 275318
rect 239876 271726 239904 275810
rect 239864 271720 239916 271726
rect 239864 271662 239916 271668
rect 240416 271448 240468 271454
rect 240416 271390 240468 271396
rect 239324 267706 239444 267734
rect 239508 267706 239628 267734
rect 239128 267300 239180 267306
rect 239128 267242 239180 267248
rect 239140 264316 239168 267242
rect 239416 264466 239444 267706
rect 239600 266422 239628 267706
rect 239588 266416 239640 266422
rect 239588 266358 239640 266364
rect 239416 264438 239536 264466
rect 239508 264330 239536 264438
rect 240428 264330 240456 271390
rect 241440 269822 241468 278038
rect 241992 269958 242020 278052
rect 243188 275602 243216 278052
rect 244398 278038 244688 278066
rect 243176 275596 243228 275602
rect 243176 275538 243228 275544
rect 243084 275324 243136 275330
rect 243084 275266 243136 275272
rect 242440 270088 242492 270094
rect 242440 270030 242492 270036
rect 241980 269952 242032 269958
rect 241980 269894 242032 269900
rect 241428 269816 241480 269822
rect 241428 269758 241480 269764
rect 241612 267436 241664 267442
rect 241612 267378 241664 267384
rect 239508 264302 239982 264330
rect 240428 264302 240810 264330
rect 241624 264316 241652 267378
rect 242452 264316 242480 270030
rect 243096 265674 243124 275266
rect 243268 273080 243320 273086
rect 243268 273022 243320 273028
rect 243084 265668 243136 265674
rect 243084 265610 243136 265616
rect 243280 264316 243308 273022
rect 244464 272944 244516 272950
rect 244464 272886 244516 272892
rect 243820 265668 243872 265674
rect 243820 265610 243872 265616
rect 243832 264330 243860 265610
rect 244476 264330 244504 272886
rect 244660 271318 244688 278038
rect 244648 271312 244700 271318
rect 244648 271254 244700 271260
rect 245580 268666 245608 278052
rect 246790 278038 246988 278066
rect 247894 278038 248368 278066
rect 245568 268660 245620 268666
rect 245568 268602 245620 268608
rect 245752 268524 245804 268530
rect 245752 268466 245804 268472
rect 243832 264302 244122 264330
rect 244476 264302 244950 264330
rect 245764 264316 245792 268466
rect 246960 267170 246988 278038
rect 247224 271584 247276 271590
rect 247224 271526 247276 271532
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 246580 266416 246632 266422
rect 246580 266358 246632 266364
rect 246592 264316 246620 266358
rect 247236 264330 247264 271526
rect 247868 270360 247920 270366
rect 247868 270302 247920 270308
rect 247880 264330 247908 270302
rect 248340 270094 248368 278038
rect 248880 274508 248932 274514
rect 248880 274450 248932 274456
rect 248328 270088 248380 270094
rect 248328 270030 248380 270036
rect 248892 266558 248920 274450
rect 249076 274378 249104 278052
rect 249064 274372 249116 274378
rect 249064 274314 249116 274320
rect 250272 271454 250300 278052
rect 250444 273964 250496 273970
rect 250444 273906 250496 273912
rect 250260 271448 250312 271454
rect 250260 271390 250312 271396
rect 249892 270224 249944 270230
rect 249892 270166 249944 270172
rect 249064 266892 249116 266898
rect 249064 266834 249116 266840
rect 248880 266552 248932 266558
rect 248880 266494 248932 266500
rect 247236 264302 247434 264330
rect 247880 264302 248262 264330
rect 249076 264316 249104 266834
rect 249904 264316 249932 270166
rect 250456 266422 250484 273906
rect 251468 272814 251496 278052
rect 251916 275460 251968 275466
rect 251916 275402 251968 275408
rect 251456 272808 251508 272814
rect 251456 272750 251508 272756
rect 251732 271176 251784 271182
rect 251732 271118 251784 271124
rect 251744 267734 251772 271118
rect 251928 267734 251956 275402
rect 252664 272950 252692 278052
rect 253388 275732 253440 275738
rect 253388 275674 253440 275680
rect 252652 272944 252704 272950
rect 252652 272886 252704 272892
rect 253204 268388 253256 268394
rect 253204 268330 253256 268336
rect 251744 267706 251864 267734
rect 251928 267706 252048 267734
rect 250720 266552 250772 266558
rect 250720 266494 250772 266500
rect 250444 266416 250496 266422
rect 250444 266358 250496 266364
rect 250732 264316 250760 266494
rect 251548 266416 251600 266422
rect 251548 266358 251600 266364
rect 251560 264316 251588 266358
rect 251836 264330 251864 267706
rect 252020 266762 252048 267706
rect 252008 266756 252060 266762
rect 252008 266698 252060 266704
rect 251836 264302 252402 264330
rect 253216 264316 253244 268330
rect 253400 266422 253428 275674
rect 253860 274718 253888 278052
rect 253848 274712 253900 274718
rect 253848 274654 253900 274660
rect 253940 272536 253992 272542
rect 253940 272478 253992 272484
rect 253388 266416 253440 266422
rect 253388 266358 253440 266364
rect 253952 265674 253980 272478
rect 254124 271720 254176 271726
rect 254124 271662 254176 271668
rect 253940 265668 253992 265674
rect 253940 265610 253992 265616
rect 254136 265554 254164 271662
rect 254964 271182 254992 278052
rect 255320 275596 255372 275602
rect 255320 275538 255372 275544
rect 255332 274242 255360 275538
rect 256160 275330 256188 278052
rect 257356 275602 257384 278052
rect 257344 275596 257396 275602
rect 257344 275538 257396 275544
rect 256148 275324 256200 275330
rect 256148 275266 256200 275272
rect 258356 274712 258408 274718
rect 258356 274654 258408 274660
rect 255320 274236 255372 274242
rect 255320 274178 255372 274184
rect 255412 274100 255464 274106
rect 255412 274042 255464 274048
rect 254952 271176 255004 271182
rect 254952 271118 255004 271124
rect 254492 265668 254544 265674
rect 254492 265610 254544 265616
rect 254044 265526 254164 265554
rect 254044 264316 254072 265526
rect 254504 264330 254532 265610
rect 255424 264330 255452 274042
rect 256976 273964 257028 273970
rect 256976 273906 257028 273912
rect 256516 266416 256568 266422
rect 256516 266358 256568 266364
rect 254504 264302 254886 264330
rect 255424 264302 255714 264330
rect 256528 264316 256556 266358
rect 256988 264330 257016 273906
rect 258080 272672 258132 272678
rect 258080 272614 258132 272620
rect 258092 264330 258120 272614
rect 258368 268394 258396 274654
rect 258552 273970 258580 278052
rect 258540 273964 258592 273970
rect 258540 273906 258592 273912
rect 259748 270230 259776 278052
rect 260958 278038 261248 278066
rect 261024 274236 261076 274242
rect 261024 274178 261076 274184
rect 259736 270224 259788 270230
rect 259736 270166 259788 270172
rect 260380 269952 260432 269958
rect 260380 269894 260432 269900
rect 259828 269816 259880 269822
rect 259828 269758 259880 269764
rect 258356 268388 258408 268394
rect 258356 268330 258408 268336
rect 259000 266756 259052 266762
rect 259000 266698 259052 266704
rect 256988 264302 257370 264330
rect 258092 264302 258198 264330
rect 259012 264316 259040 266698
rect 259840 264316 259868 269758
rect 260392 264330 260420 269894
rect 261036 264330 261064 274178
rect 261220 274106 261248 278038
rect 261956 278038 262062 278066
rect 261208 274100 261260 274106
rect 261208 274042 261260 274048
rect 261956 269822 261984 278038
rect 262864 275596 262916 275602
rect 262864 275538 262916 275544
rect 262220 271312 262272 271318
rect 262220 271254 262272 271260
rect 261944 269816 261996 269822
rect 261944 269758 261996 269764
rect 262232 264330 262260 271254
rect 262876 270366 262904 275538
rect 263244 275466 263272 278052
rect 263232 275460 263284 275466
rect 263232 275402 263284 275408
rect 264440 272542 264468 278052
rect 265256 274372 265308 274378
rect 265256 274314 265308 274320
rect 264428 272536 264480 272542
rect 264428 272478 264480 272484
rect 262864 270360 262916 270366
rect 262864 270302 262916 270308
rect 264796 270088 264848 270094
rect 264796 270030 264848 270036
rect 263140 268660 263192 268666
rect 263140 268602 263192 268608
rect 260392 264302 260682 264330
rect 261036 264302 261510 264330
rect 262232 264302 262338 264330
rect 263152 264316 263180 268602
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 263980 264316 264008 267106
rect 264808 264316 264836 270030
rect 265268 264330 265296 274314
rect 265636 271454 265664 278052
rect 266832 272678 266860 278052
rect 268028 274718 268056 278052
rect 268844 275324 268896 275330
rect 268844 275266 268896 275272
rect 268016 274712 268068 274718
rect 268016 274654 268068 274660
rect 267924 272944 267976 272950
rect 267924 272886 267976 272892
rect 267004 272808 267056 272814
rect 267004 272750 267056 272756
rect 266820 272672 266872 272678
rect 266820 272614 266872 272620
rect 265624 271448 265676 271454
rect 265624 271390 265676 271396
rect 266452 271312 266504 271318
rect 266452 271254 266504 271260
rect 265268 264302 265650 264330
rect 266464 264316 266492 271254
rect 267016 264330 267044 272750
rect 267936 264330 267964 272886
rect 268856 271930 268884 275266
rect 269224 275126 269252 278052
rect 269212 275120 269264 275126
rect 269212 275062 269264 275068
rect 268844 271924 268896 271930
rect 268844 271866 268896 271872
rect 270328 271182 270356 278052
rect 271524 272814 271552 278052
rect 272432 274712 272484 274718
rect 272432 274654 272484 274660
rect 272064 273964 272116 273970
rect 272064 273906 272116 273912
rect 271512 272808 271564 272814
rect 271512 272750 271564 272756
rect 270500 271924 270552 271930
rect 270500 271866 270552 271872
rect 269304 271176 269356 271182
rect 269304 271118 269356 271124
rect 270316 271176 270368 271182
rect 270316 271118 270368 271124
rect 268936 268388 268988 268394
rect 268936 268330 268988 268336
rect 267016 264302 267306 264330
rect 267936 264302 268134 264330
rect 268948 264316 268976 268330
rect 269316 264330 269344 271118
rect 270512 264330 270540 271866
rect 271420 270224 271472 270230
rect 271420 270166 271472 270172
rect 269316 264302 269790 264330
rect 270512 264302 270618 264330
rect 271432 264316 271460 270166
rect 272076 264330 272104 273906
rect 272444 269278 272472 274654
rect 272720 273970 272748 278052
rect 273260 275460 273312 275466
rect 273260 275402 273312 275408
rect 272708 273964 272760 273970
rect 272708 273906 272760 273912
rect 273076 269952 273128 269958
rect 273076 269894 273128 269900
rect 272432 269272 272484 269278
rect 272432 269214 272484 269220
rect 272076 264302 272274 264330
rect 273088 264316 273116 269894
rect 273272 269006 273300 275402
rect 273916 275330 273944 278052
rect 273904 275324 273956 275330
rect 273904 275266 273956 275272
rect 274916 275120 274968 275126
rect 274916 275062 274968 275068
rect 273536 274100 273588 274106
rect 273536 274042 273588 274048
rect 273260 269000 273312 269006
rect 273260 268942 273312 268948
rect 273548 264330 273576 274042
rect 274732 269816 274784 269822
rect 274732 269758 274784 269764
rect 273548 264302 273930 264330
rect 274744 264316 274772 269758
rect 274928 269142 274956 275062
rect 275112 274106 275140 278052
rect 276322 278038 276704 278066
rect 275100 274100 275152 274106
rect 275100 274042 275152 274048
rect 276020 272536 276072 272542
rect 276020 272478 276072 272484
rect 274916 269136 274968 269142
rect 274916 269078 274968 269084
rect 275560 269000 275612 269006
rect 275560 268942 275612 268948
rect 275572 264316 275600 268942
rect 276032 264330 276060 272478
rect 276676 271318 276704 278038
rect 277504 275670 277532 278052
rect 277492 275664 277544 275670
rect 277492 275606 277544 275612
rect 278608 273154 278636 278052
rect 279818 278038 280108 278066
rect 278596 273148 278648 273154
rect 278596 273090 278648 273096
rect 277584 272672 277636 272678
rect 277584 272614 277636 272620
rect 276848 271448 276900 271454
rect 276848 271390 276900 271396
rect 276664 271312 276716 271318
rect 276664 271254 276716 271260
rect 276860 264330 276888 271390
rect 277596 264330 277624 272614
rect 280080 269822 280108 278038
rect 280344 272808 280396 272814
rect 280344 272750 280396 272756
rect 280068 269816 280120 269822
rect 280068 269758 280120 269764
rect 278872 269272 278924 269278
rect 278872 269214 278924 269220
rect 276032 264302 276414 264330
rect 276860 264302 277242 264330
rect 277596 264302 278070 264330
rect 278884 264316 278912 269214
rect 279700 269136 279752 269142
rect 279700 269078 279752 269084
rect 279712 264316 279740 269078
rect 280356 265674 280384 272750
rect 281000 272678 281028 278052
rect 282196 274310 282224 278052
rect 282920 275324 282972 275330
rect 282920 275266 282972 275272
rect 282184 274304 282236 274310
rect 282184 274246 282236 274252
rect 281816 273964 281868 273970
rect 281816 273906 281868 273912
rect 280988 272672 281040 272678
rect 280988 272614 281040 272620
rect 280528 271176 280580 271182
rect 280528 271118 280580 271124
rect 280344 265668 280396 265674
rect 280344 265610 280396 265616
rect 280540 264316 280568 271118
rect 280988 265668 281040 265674
rect 280988 265610 281040 265616
rect 281000 264330 281028 265610
rect 281828 264330 281856 273906
rect 282932 264330 282960 275266
rect 283392 274718 283420 278052
rect 284588 275874 284616 278052
rect 284576 275868 284628 275874
rect 284576 275810 284628 275816
rect 284300 275664 284352 275670
rect 284300 275606 284352 275612
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283472 274100 283524 274106
rect 283472 274042 283524 274048
rect 283484 264330 283512 274042
rect 284312 265674 284340 275606
rect 285692 275466 285720 278052
rect 286888 275602 286916 278052
rect 286876 275596 286928 275602
rect 286876 275538 286928 275544
rect 285680 275460 285732 275466
rect 285680 275402 285732 275408
rect 288084 275058 288112 278052
rect 288072 275052 288124 275058
rect 288072 274994 288124 275000
rect 289280 274854 289308 278052
rect 290096 275868 290148 275874
rect 290096 275810 290148 275816
rect 289268 274848 289320 274854
rect 289268 274790 289320 274796
rect 289176 274712 289228 274718
rect 289176 274654 289228 274660
rect 287704 274304 287756 274310
rect 287704 274246 287756 274252
rect 285864 273148 285916 273154
rect 285864 273090 285916 273096
rect 284484 271312 284536 271318
rect 284484 271254 284536 271260
rect 284300 265668 284352 265674
rect 284300 265610 284352 265616
rect 284496 264330 284524 271254
rect 285220 265668 285272 265674
rect 285220 265610 285272 265616
rect 285232 264330 285260 265610
rect 285876 264330 285904 273090
rect 286324 272672 286376 272678
rect 286324 272614 286376 272620
rect 286336 266898 286364 272614
rect 287152 269816 287204 269822
rect 287152 269758 287204 269764
rect 286324 266892 286376 266898
rect 286324 266834 286376 266840
rect 281000 264302 281382 264330
rect 281828 264302 282210 264330
rect 282932 264302 283038 264330
rect 283484 264302 283866 264330
rect 284496 264302 284694 264330
rect 285232 264302 285522 264330
rect 285876 264302 286350 264330
rect 287164 264316 287192 269758
rect 287716 266422 287744 274246
rect 287980 266892 288032 266898
rect 287980 266834 288032 266840
rect 287704 266416 287756 266422
rect 287704 266358 287756 266364
rect 287992 264316 288020 266834
rect 288808 266416 288860 266422
rect 288808 266358 288860 266364
rect 288820 264316 288848 266358
rect 289188 264330 289216 274654
rect 290108 264330 290136 275810
rect 290476 275330 290504 278052
rect 291672 275670 291700 278052
rect 291660 275664 291712 275670
rect 291660 275606 291712 275612
rect 291752 275528 291804 275534
rect 291752 275470 291804 275476
rect 291200 275460 291252 275466
rect 291200 275402 291252 275408
rect 290464 275324 290516 275330
rect 290464 275266 290516 275272
rect 291212 264330 291240 275402
rect 291764 264330 291792 275470
rect 292868 275194 292896 278052
rect 292856 275188 292908 275194
rect 292856 275130 292908 275136
rect 292672 275052 292724 275058
rect 292672 274994 292724 275000
rect 292684 264330 292712 274994
rect 293972 274990 294000 278052
rect 294144 275324 294196 275330
rect 294144 275266 294196 275272
rect 293960 274984 294012 274990
rect 293960 274926 294012 274932
rect 293408 274848 293460 274854
rect 293408 274790 293460 274796
rect 293420 264330 293448 274790
rect 294156 264330 294184 275266
rect 295168 274718 295196 278052
rect 295340 275664 295392 275670
rect 295340 275606 295392 275612
rect 295156 274712 295208 274718
rect 295156 274654 295208 274660
rect 295352 264330 295380 275606
rect 295800 275188 295852 275194
rect 295800 275130 295852 275136
rect 295812 264330 295840 275130
rect 296364 274854 296392 278052
rect 297180 274984 297232 274990
rect 297180 274926 297232 274932
rect 296352 274848 296404 274854
rect 296352 274790 296404 274796
rect 296812 274712 296864 274718
rect 296812 274654 296864 274660
rect 296824 265674 296852 274654
rect 297192 267734 297220 274926
rect 297560 274718 297588 278052
rect 298756 275262 298784 278052
rect 299952 275398 299980 278052
rect 299940 275392 299992 275398
rect 299940 275334 299992 275340
rect 298744 275256 298796 275262
rect 298744 275198 298796 275204
rect 300032 275256 300084 275262
rect 300032 275198 300084 275204
rect 298376 274848 298428 274854
rect 298376 274790 298428 274796
rect 297548 274712 297600 274718
rect 297548 274654 297600 274660
rect 297100 267706 297220 267734
rect 296812 265668 296864 265674
rect 296812 265610 296864 265616
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291212 264302 291318 264330
rect 291764 264302 292146 264330
rect 292684 264302 292974 264330
rect 293420 264302 293802 264330
rect 294156 264302 294630 264330
rect 295352 264302 295458 264330
rect 295812 264302 296286 264330
rect 297100 264316 297128 267706
rect 297548 265668 297600 265674
rect 297548 265610 297600 265616
rect 297560 264330 297588 265610
rect 298388 264330 298416 274790
rect 299572 274712 299624 274718
rect 299572 274654 299624 274660
rect 297560 264302 297942 264330
rect 298388 264302 298770 264330
rect 299584 264316 299612 274654
rect 300044 264330 300072 275198
rect 301056 266422 301084 278052
rect 302266 278038 302464 278066
rect 301228 275392 301280 275398
rect 301228 275334 301280 275340
rect 301044 266416 301096 266422
rect 301044 266358 301096 266364
rect 300044 264302 300426 264330
rect 301240 264316 301268 275334
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 302068 264316 302096 266358
rect 302436 264330 302464 278038
rect 303448 274718 303476 278052
rect 303724 278038 304658 278066
rect 305012 278038 305854 278066
rect 306392 278038 307050 278066
rect 307772 278038 308154 278066
rect 309152 278038 309350 278066
rect 303436 274712 303488 274718
rect 303436 274654 303488 274660
rect 303724 266422 303752 278038
rect 303988 274712 304040 274718
rect 303988 274654 304040 274660
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 304000 264330 304028 274654
rect 304540 266416 304592 266422
rect 304540 266358 304592 266364
rect 302436 264302 302910 264330
rect 303738 264302 304028 264330
rect 304552 264316 304580 266358
rect 305012 264330 305040 278038
rect 306392 266370 306420 278038
rect 307772 267734 307800 278038
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266688 308732 266694
rect 308680 266630 308732 266636
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266630
rect 309152 266422 309180 278038
rect 310532 266694 310560 278052
rect 310992 278038 311742 278066
rect 311912 278038 312938 278066
rect 313292 278038 314134 278066
rect 314672 278038 315238 278066
rect 316052 278038 316434 278066
rect 317432 278038 317630 278066
rect 310520 266688 310572 266694
rect 310520 266630 310572 266636
rect 310336 266552 310388 266558
rect 310336 266494 310388 266500
rect 309140 266416 309192 266422
rect 309140 266358 309192 266364
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309520 264316 309548 266358
rect 310348 264316 310376 266494
rect 310992 266422 311020 278038
rect 311912 266558 311940 278038
rect 312820 267164 312872 267170
rect 312820 267106 312872 267112
rect 311900 266552 311952 266558
rect 311900 266494 311952 266500
rect 312268 266552 312320 266558
rect 312268 266494 312320 266500
rect 310980 266416 311032 266422
rect 310980 266358 311032 266364
rect 311164 266416 311216 266422
rect 311164 266358 311216 266364
rect 311176 264316 311204 266358
rect 312280 264330 312308 266494
rect 312018 264302 312308 264330
rect 312832 264316 312860 267106
rect 313292 266422 313320 278038
rect 314476 267300 314528 267306
rect 314476 267242 314528 267248
rect 313648 266756 313700 266762
rect 313648 266698 313700 266704
rect 313280 266416 313332 266422
rect 313280 266358 313332 266364
rect 313660 264316 313688 266698
rect 314488 264316 314516 267242
rect 314672 266558 314700 278038
rect 315304 267436 315356 267442
rect 315304 267378 315356 267384
rect 314660 266552 314712 266558
rect 314660 266494 314712 266500
rect 315316 264316 315344 267378
rect 316052 267170 316080 278038
rect 316040 267164 316092 267170
rect 316040 267106 316092 267112
rect 316960 267028 317012 267034
rect 316960 266970 317012 266976
rect 316132 266552 316184 266558
rect 316132 266494 316184 266500
rect 316144 264316 316172 266494
rect 316972 264316 317000 266970
rect 317432 266762 317460 278038
rect 318616 273284 318668 273290
rect 318616 273226 318668 273232
rect 317420 266756 317472 266762
rect 317420 266698 317472 266704
rect 317788 266688 317840 266694
rect 317788 266630 317840 266636
rect 317800 264316 317828 266630
rect 318628 264316 318656 273226
rect 318812 267306 318840 278052
rect 318996 278038 320022 278066
rect 320192 278038 321218 278066
rect 321940 278038 322414 278066
rect 322952 278038 323518 278066
rect 318996 267442 319024 278038
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 318984 267436 319036 267442
rect 318984 267378 319036 267384
rect 318800 267300 318852 267306
rect 318800 267242 318852 267248
rect 319456 264316 319484 269078
rect 320192 266558 320220 278038
rect 321192 274712 321244 274718
rect 321192 274654 321244 274660
rect 321204 267734 321232 274654
rect 321376 270768 321428 270774
rect 321376 270710 321428 270716
rect 321112 267706 321232 267734
rect 320180 266552 320232 266558
rect 320180 266494 320232 266500
rect 320272 266416 320324 266422
rect 320272 266358 320324 266364
rect 320284 264316 320312 266358
rect 321112 264316 321140 267706
rect 321388 266422 321416 270710
rect 321940 267034 321968 278038
rect 322756 272672 322808 272678
rect 322756 272614 322808 272620
rect 321928 267028 321980 267034
rect 321928 266970 321980 266976
rect 321928 266892 321980 266898
rect 321928 266834 321980 266840
rect 321376 266416 321428 266422
rect 321376 266358 321428 266364
rect 321940 264316 321968 266834
rect 322768 264316 322796 272614
rect 322952 266694 322980 278038
rect 324044 273964 324096 273970
rect 324044 273906 324096 273912
rect 322940 266688 322992 266694
rect 322940 266630 322992 266636
rect 324056 264330 324084 273906
rect 324700 273290 324728 278052
rect 325712 278038 325910 278066
rect 325332 274236 325384 274242
rect 325332 274178 325384 274184
rect 324688 273284 324740 273290
rect 324688 273226 324740 273232
rect 325344 266422 325372 274178
rect 325516 272536 325568 272542
rect 325516 272478 325568 272484
rect 324412 266416 324464 266422
rect 324412 266358 324464 266364
rect 325332 266416 325384 266422
rect 325332 266358 325384 266364
rect 323610 264302 324084 264330
rect 324424 264316 324452 266358
rect 325528 264330 325556 272478
rect 325712 269142 325740 278038
rect 326436 271040 326488 271046
rect 326436 270982 326488 270988
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 270982
rect 327092 270774 327120 278052
rect 328288 274718 328316 278052
rect 328276 274712 328328 274718
rect 328276 274654 328328 274660
rect 329484 273290 329512 278052
rect 327540 273284 327592 273290
rect 327540 273226 327592 273232
rect 329472 273284 329524 273290
rect 329472 273226 329524 273232
rect 327080 270768 327132 270774
rect 327080 270710 327132 270716
rect 326896 269952 326948 269958
rect 326896 269894 326948 269900
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269894
rect 327552 266898 327580 273226
rect 329472 273080 329524 273086
rect 329472 273022 329524 273028
rect 327724 270088 327776 270094
rect 327724 270030 327776 270036
rect 327540 266892 327592 266898
rect 327540 266834 327592 266840
rect 327736 264316 327764 270030
rect 329484 266422 329512 273022
rect 330588 272678 330616 278052
rect 331784 273970 331812 278052
rect 332980 274242 333008 278052
rect 333796 274372 333848 274378
rect 333796 274314 333848 274320
rect 332968 274236 333020 274242
rect 332968 274178 333020 274184
rect 332324 274100 332376 274106
rect 332324 274042 332376 274048
rect 331772 273964 331824 273970
rect 331772 273906 331824 273912
rect 331956 273964 332008 273970
rect 331956 273906 332008 273912
rect 330576 272672 330628 272678
rect 330576 272614 330628 272620
rect 329656 271312 329708 271318
rect 329656 271254 329708 271260
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 329472 266416 329524 266422
rect 329472 266358 329524 266364
rect 328564 264316 328592 266358
rect 329668 264330 329696 271254
rect 331128 271176 331180 271182
rect 331128 271118 331180 271124
rect 331140 267734 331168 271118
rect 331048 267706 331168 267734
rect 330208 266416 330260 266422
rect 330208 266358 330260 266364
rect 329406 264302 329696 264330
rect 330220 264316 330248 266358
rect 331048 264316 331076 267706
rect 331968 266422 331996 273906
rect 331956 266416 332008 266422
rect 331956 266358 332008 266364
rect 332336 264330 332364 274042
rect 332692 266892 332744 266898
rect 332692 266834 332744 266840
rect 331890 264302 332364 264330
rect 332704 264316 332732 266834
rect 333808 264330 333836 274314
rect 334176 272542 334204 278052
rect 335372 274666 335400 278052
rect 335096 274638 335400 274666
rect 335556 278038 336582 278066
rect 336752 278038 337778 278066
rect 334164 272536 334216 272542
rect 334164 272478 334216 272484
rect 335096 271046 335124 274638
rect 335268 272944 335320 272950
rect 335268 272886 335320 272892
rect 335084 271040 335136 271046
rect 335084 270982 335136 270988
rect 335084 269816 335136 269822
rect 335084 269758 335136 269764
rect 334348 266416 334400 266422
rect 334348 266358 334400 266364
rect 333546 264302 333836 264330
rect 334360 264316 334388 266358
rect 335096 264330 335124 269758
rect 335280 266422 335308 272886
rect 335556 269958 335584 278038
rect 336372 272808 336424 272814
rect 336372 272750 336424 272756
rect 335544 269952 335596 269958
rect 335544 269894 335596 269900
rect 335268 266416 335320 266422
rect 335268 266358 335320 266364
rect 336384 264330 336412 272750
rect 336752 270094 336780 278038
rect 338868 273086 338896 278052
rect 338856 273080 338908 273086
rect 338856 273022 338908 273028
rect 338028 272672 338080 272678
rect 338028 272614 338080 272620
rect 336740 270088 336792 270094
rect 336740 270030 336792 270036
rect 336832 269952 336884 269958
rect 336832 269894 336884 269900
rect 335096 264302 335202 264330
rect 336030 264302 336412 264330
rect 336844 264316 336872 269894
rect 338040 264330 338068 272614
rect 339224 271448 339276 271454
rect 339224 271390 339276 271396
rect 338488 268524 338540 268530
rect 338488 268466 338540 268472
rect 337686 264302 338068 264330
rect 338500 264316 338528 268466
rect 339236 264330 339264 271390
rect 340064 271318 340092 278052
rect 341260 273970 341288 278052
rect 341248 273964 341300 273970
rect 341248 273906 341300 273912
rect 342076 273964 342128 273970
rect 342076 273906 342128 273912
rect 340052 271312 340104 271318
rect 340052 271254 340104 271260
rect 340604 271312 340656 271318
rect 340604 271254 340656 271260
rect 340616 264330 340644 271254
rect 340972 267572 341024 267578
rect 340972 267514 341024 267520
rect 339236 264302 339342 264330
rect 340170 264302 340644 264330
rect 340984 264316 341012 267514
rect 342088 264330 342116 273906
rect 342456 271182 342484 278052
rect 343456 274236 343508 274242
rect 343456 274178 343508 274184
rect 342444 271176 342496 271182
rect 342444 271118 342496 271124
rect 342628 266688 342680 266694
rect 342628 266630 342680 266636
rect 341826 264302 342116 264330
rect 342640 264316 342668 266630
rect 343468 264316 343496 274178
rect 343652 274106 343680 278052
rect 343836 278038 344862 278066
rect 343640 274100 343692 274106
rect 343640 274042 343692 274048
rect 343836 266898 343864 278038
rect 345952 274378 345980 278052
rect 346872 278038 347162 278066
rect 347792 278038 348358 278066
rect 345940 274372 345992 274378
rect 345940 274314 345992 274320
rect 346872 272950 346900 278038
rect 347044 274372 347096 274378
rect 347044 274314 347096 274320
rect 346860 272944 346912 272950
rect 346860 272886 346912 272892
rect 344652 272536 344704 272542
rect 344652 272478 344704 272484
rect 343824 266892 343876 266898
rect 343824 266834 343876 266840
rect 344664 264330 344692 272478
rect 345112 270224 345164 270230
rect 345112 270166 345164 270172
rect 344310 264302 344692 264330
rect 345124 264316 345152 270166
rect 345940 270088 345992 270094
rect 345940 270030 345992 270036
rect 345952 264316 345980 270030
rect 347056 266694 347084 274314
rect 347596 271176 347648 271182
rect 347596 271118 347648 271124
rect 347044 266688 347096 266694
rect 347044 266630 347096 266636
rect 347412 266552 347464 266558
rect 347412 266494 347464 266500
rect 346768 266416 346820 266422
rect 346768 266358 346820 266364
rect 346780 264316 346808 266358
rect 347424 264330 347452 266494
rect 347608 266422 347636 271118
rect 347792 269822 347820 278038
rect 349540 272814 349568 278052
rect 350552 278038 350750 278066
rect 350356 274100 350408 274106
rect 350356 274042 350408 274048
rect 349804 273080 349856 273086
rect 349804 273022 349856 273028
rect 349528 272808 349580 272814
rect 349528 272750 349580 272756
rect 347780 269816 347832 269822
rect 347780 269758 347832 269764
rect 348424 268388 348476 268394
rect 348424 268330 348476 268336
rect 347596 266416 347648 266422
rect 347596 266358 347648 266364
rect 347424 264302 347622 264330
rect 348436 264316 348464 268330
rect 349816 266558 349844 273022
rect 350080 267436 350132 267442
rect 350080 267378 350132 267384
rect 349804 266552 349856 266558
rect 349804 266494 349856 266500
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 349264 264316 349292 266358
rect 350092 264316 350120 267378
rect 350368 266422 350396 274042
rect 350552 269958 350580 278038
rect 350724 274712 350776 274718
rect 350724 274654 350776 274660
rect 350540 269952 350592 269958
rect 350540 269894 350592 269900
rect 350736 268530 350764 274654
rect 351932 272678 351960 278052
rect 353128 274718 353156 278052
rect 353116 274712 353168 274718
rect 353116 274654 353168 274660
rect 352564 272808 352616 272814
rect 352564 272750 352616 272756
rect 351920 272672 351972 272678
rect 351920 272614 351972 272620
rect 351736 269952 351788 269958
rect 351736 269894 351788 269900
rect 350724 268524 350776 268530
rect 350724 268466 350776 268472
rect 350908 266552 350960 266558
rect 350908 266494 350960 266500
rect 350356 266416 350408 266422
rect 350356 266358 350408 266364
rect 350920 264316 350948 266494
rect 351748 264316 351776 269894
rect 352576 266558 352604 272750
rect 353944 271720 353996 271726
rect 353944 271662 353996 271668
rect 353392 267300 353444 267306
rect 353392 267242 353444 267248
rect 352564 266552 352616 266558
rect 352564 266494 352616 266500
rect 352564 266416 352616 266422
rect 352564 266358 352616 266364
rect 352576 264316 352604 266358
rect 353404 264316 353432 267242
rect 353956 266422 353984 271662
rect 354232 271454 354260 278052
rect 355152 278038 355442 278066
rect 354496 272672 354548 272678
rect 354496 272614 354548 272620
rect 354220 271448 354272 271454
rect 354220 271390 354272 271396
rect 353944 266416 353996 266422
rect 353944 266358 353996 266364
rect 354508 264330 354536 272614
rect 355152 271318 355180 278038
rect 356624 271862 356652 278052
rect 357820 273970 357848 278052
rect 358084 274508 358136 274514
rect 358084 274450 358136 274456
rect 357808 273964 357860 273970
rect 357808 273906 357860 273912
rect 355324 271856 355376 271862
rect 355324 271798 355376 271804
rect 356612 271856 356664 271862
rect 356612 271798 356664 271804
rect 355140 271312 355192 271318
rect 355140 271254 355192 271260
rect 355048 269816 355100 269822
rect 355048 269758 355100 269764
rect 354246 264302 354536 264330
rect 355060 264316 355088 269758
rect 355336 267578 355364 271798
rect 357164 271584 357216 271590
rect 357164 271526 357216 271532
rect 355324 267572 355376 267578
rect 355324 267514 355376 267520
rect 355876 266824 355928 266830
rect 355876 266766 355928 266772
rect 355888 264316 355916 266766
rect 357176 264330 357204 271526
rect 358096 267442 358124 274450
rect 359016 274378 359044 278052
rect 359004 274372 359056 274378
rect 359004 274314 359056 274320
rect 360212 274242 360240 278052
rect 361212 275324 361264 275330
rect 361212 275266 361264 275272
rect 360200 274236 360252 274242
rect 360200 274178 360252 274184
rect 360108 273964 360160 273970
rect 360108 273906 360160 273912
rect 358728 271448 358780 271454
rect 358728 271390 358780 271396
rect 358084 267436 358136 267442
rect 358084 267378 358136 267384
rect 357532 266552 357584 266558
rect 357532 266494 357584 266500
rect 356730 264302 357204 264330
rect 357544 264316 357572 266494
rect 358740 264330 358768 271390
rect 359832 268524 359884 268530
rect 359832 268466 359884 268472
rect 359844 266558 359872 268466
rect 359832 266552 359884 266558
rect 359832 266494 359884 266500
rect 360120 266422 360148 273906
rect 359188 266416 359240 266422
rect 359188 266358 359240 266364
rect 360108 266416 360160 266422
rect 360108 266358 360160 266364
rect 358386 264302 358768 264330
rect 359200 264316 359228 266358
rect 360016 266280 360068 266286
rect 360016 266222 360068 266228
rect 360028 264316 360056 266222
rect 361224 264330 361252 275266
rect 361408 272542 361436 278052
rect 361592 278038 362526 278066
rect 362972 278038 363722 278066
rect 364536 278038 364918 278066
rect 361396 272536 361448 272542
rect 361396 272478 361448 272484
rect 361592 270230 361620 278038
rect 362776 272944 362828 272950
rect 362776 272886 362828 272892
rect 361580 270224 361632 270230
rect 361580 270166 361632 270172
rect 362500 267436 362552 267442
rect 362500 267378 362552 267384
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 360870 264302 361252 264330
rect 361684 264316 361712 266358
rect 362512 264316 362540 267378
rect 362788 266422 362816 272886
rect 362972 270094 363000 278038
rect 363788 272536 363840 272542
rect 363788 272478 363840 272484
rect 362960 270088 363012 270094
rect 362960 270030 363012 270036
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 363800 264330 363828 272478
rect 364536 271182 364564 278038
rect 364984 274236 365036 274242
rect 364984 274178 365036 274184
rect 364524 271176 364576 271182
rect 364524 271118 364576 271124
rect 364156 270224 364208 270230
rect 364156 270166 364208 270172
rect 363354 264302 363828 264330
rect 364168 264316 364196 270166
rect 364996 267306 365024 274178
rect 366100 273086 366128 278052
rect 367112 278038 367310 278066
rect 366364 273216 366416 273222
rect 366364 273158 366416 273164
rect 366088 273080 366140 273086
rect 366088 273022 366140 273028
rect 365444 271312 365496 271318
rect 365444 271254 365496 271260
rect 364984 267300 365036 267306
rect 364984 267242 365036 267248
rect 365456 264330 365484 271254
rect 365812 267164 365864 267170
rect 365812 267106 365864 267112
rect 365010 264302 365484 264330
rect 365824 264316 365852 267106
rect 366376 266558 366404 273158
rect 366916 271176 366968 271182
rect 366916 271118 366968 271124
rect 366364 266552 366416 266558
rect 366364 266494 366416 266500
rect 366928 264330 366956 271118
rect 367112 268394 367140 278038
rect 368492 274106 368520 278052
rect 369596 274514 369624 278052
rect 369584 274508 369636 274514
rect 369584 274450 369636 274456
rect 369124 274372 369176 274378
rect 369124 274314 369176 274320
rect 368480 274100 368532 274106
rect 368480 274042 368532 274048
rect 367468 270360 367520 270366
rect 367468 270302 367520 270308
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 366666 264302 366956 264330
rect 367480 264316 367508 270302
rect 369136 266422 369164 274314
rect 369308 274100 369360 274106
rect 369308 274042 369360 274048
rect 369320 267442 369348 274042
rect 370792 272814 370820 278052
rect 371252 278038 372002 278066
rect 372816 278038 373198 278066
rect 370780 272808 370832 272814
rect 370780 272750 370832 272756
rect 369860 270088 369912 270094
rect 369860 270030 369912 270036
rect 369308 267436 369360 267442
rect 369308 267378 369360 267384
rect 369872 266422 369900 270030
rect 371252 269958 371280 278038
rect 372816 271726 372844 278038
rect 373264 274372 373316 274378
rect 373264 274314 373316 274320
rect 372804 271720 372856 271726
rect 372804 271662 372856 271668
rect 371240 269952 371292 269958
rect 371240 269894 371292 269900
rect 372436 269952 372488 269958
rect 372436 269894 372488 269900
rect 372160 268388 372212 268394
rect 372160 268330 372212 268336
rect 370780 267572 370832 267578
rect 370780 267514 370832 267520
rect 368296 266416 368348 266422
rect 368296 266358 368348 266364
rect 369124 266416 369176 266422
rect 369124 266358 369176 266364
rect 369400 266416 369452 266422
rect 369400 266358 369452 266364
rect 369860 266416 369912 266422
rect 369860 266358 369912 266364
rect 370320 266416 370372 266422
rect 370320 266358 370372 266364
rect 368308 264316 368336 266358
rect 369412 264330 369440 266358
rect 370332 264330 370360 266358
rect 369150 264302 369440 264330
rect 369978 264302 370360 264330
rect 370792 264316 370820 267514
rect 371608 267436 371660 267442
rect 371608 267378 371660 267384
rect 371620 264316 371648 267378
rect 372172 266422 372200 268330
rect 372160 266416 372212 266422
rect 372160 266358 372212 266364
rect 372448 264316 372476 269894
rect 373276 267442 373304 274314
rect 374380 274242 374408 278052
rect 374368 274236 374420 274242
rect 374368 274178 374420 274184
rect 374644 273352 374696 273358
rect 374644 273294 374696 273300
rect 373264 267436 373316 267442
rect 373264 267378 373316 267384
rect 373264 267300 373316 267306
rect 373264 267242 373316 267248
rect 373276 264316 373304 267242
rect 374656 266830 374684 273294
rect 375196 272808 375248 272814
rect 375196 272750 375248 272756
rect 374644 266824 374696 266830
rect 374644 266766 374696 266772
rect 374920 266552 374972 266558
rect 374920 266494 374972 266500
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 266494
rect 375208 266422 375236 272750
rect 375576 272678 375604 278052
rect 376786 278038 376984 278066
rect 375564 272672 375616 272678
rect 375564 272614 375616 272620
rect 376576 271856 376628 271862
rect 376576 271798 376628 271804
rect 375748 267028 375800 267034
rect 375748 266970 375800 266976
rect 375196 266416 375248 266422
rect 375196 266358 375248 266364
rect 375760 264316 375788 266970
rect 376588 264316 376616 271798
rect 376956 269822 376984 278038
rect 377876 273358 377904 278052
rect 377864 273352 377916 273358
rect 377864 273294 377916 273300
rect 377404 273080 377456 273086
rect 377404 273022 377456 273028
rect 376944 269816 376996 269822
rect 376944 269758 376996 269764
rect 377416 267578 377444 273022
rect 379072 271590 379100 278052
rect 379532 278038 380282 278066
rect 379336 274236 379388 274242
rect 379336 274178 379388 274184
rect 379060 271584 379112 271590
rect 379060 271526 379112 271532
rect 377680 269816 377732 269822
rect 377680 269758 377732 269764
rect 377404 267572 377456 267578
rect 377404 267514 377456 267520
rect 377692 264330 377720 269758
rect 378232 267708 378284 267714
rect 378232 267650 378284 267656
rect 377430 264302 377720 264330
rect 378244 264316 378272 267650
rect 379348 264330 379376 274178
rect 379532 268530 379560 278038
rect 381464 271454 381492 278052
rect 382660 273970 382688 278052
rect 382924 274644 382976 274650
rect 382924 274586 382976 274592
rect 382648 273964 382700 273970
rect 382648 273906 382700 273912
rect 382004 272672 382056 272678
rect 382004 272614 382056 272620
rect 381452 271448 381504 271454
rect 381452 271390 381504 271396
rect 381544 271040 381596 271046
rect 381544 270982 381596 270988
rect 379704 269068 379756 269074
rect 379704 269010 379756 269016
rect 379520 268524 379572 268530
rect 379520 268466 379572 268472
rect 379716 266558 379744 269010
rect 380716 267572 380768 267578
rect 380716 267514 380768 267520
rect 379704 266552 379756 266558
rect 379704 266494 379756 266500
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379376 264330
rect 379900 264316 379928 266358
rect 380728 264316 380756 267514
rect 381556 266422 381584 270982
rect 381544 266416 381596 266422
rect 381544 266358 381596 266364
rect 382016 264330 382044 272614
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 382936 267170 382964 274586
rect 383856 273222 383884 278052
rect 385052 275330 385080 278052
rect 385880 278038 386170 278066
rect 385040 275324 385092 275330
rect 385040 275266 385092 275272
rect 383844 273216 383896 273222
rect 383844 273158 383896 273164
rect 385880 272950 385908 278038
rect 386052 275460 386104 275466
rect 386052 275402 386104 275408
rect 385868 272944 385920 272950
rect 385868 272886 385920 272892
rect 384948 271720 385000 271726
rect 384948 271662 385000 271668
rect 384764 269680 384816 269686
rect 384764 269622 384816 269628
rect 383200 267436 383252 267442
rect 383200 267378 383252 267384
rect 382924 267164 382976 267170
rect 382924 267106 382976 267112
rect 383212 264316 383240 267378
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 384040 264316 384068 266358
rect 384776 264330 384804 269622
rect 384960 266422 384988 271662
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 386064 264330 386092 275402
rect 387352 274106 387380 278052
rect 387340 274100 387392 274106
rect 387340 274042 387392 274048
rect 387432 273964 387484 273970
rect 387432 273906 387484 273912
rect 387444 266422 387472 273906
rect 388548 272542 388576 278052
rect 389192 278038 389758 278066
rect 388536 272536 388588 272542
rect 388536 272478 388588 272484
rect 388996 272400 389048 272406
rect 388996 272342 389048 272348
rect 387616 271584 387668 271590
rect 387616 271526 387668 271532
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 387432 266416 387484 266422
rect 387432 266358 387484 266364
rect 384776 264302 384882 264330
rect 385710 264302 386092 264330
rect 386524 264316 386552 266358
rect 387628 264330 387656 271526
rect 388168 266756 388220 266762
rect 388168 266698 388220 266704
rect 387366 264302 387656 264330
rect 388180 264316 388208 266698
rect 389008 264316 389036 272342
rect 389192 270230 389220 278038
rect 390940 271318 390968 278052
rect 392136 274650 392164 278052
rect 392124 274644 392176 274650
rect 392124 274586 392176 274592
rect 392584 273692 392636 273698
rect 392584 273634 392636 273640
rect 390928 271312 390980 271318
rect 390928 271254 390980 271260
rect 391848 271312 391900 271318
rect 391848 271254 391900 271260
rect 389180 270224 389232 270230
rect 389180 270166 389232 270172
rect 390100 270224 390152 270230
rect 390100 270166 390152 270172
rect 389824 268796 389876 268802
rect 389824 268738 389876 268744
rect 389836 264316 389864 268738
rect 390112 267034 390140 270166
rect 390652 267164 390704 267170
rect 390652 267106 390704 267112
rect 390100 267028 390152 267034
rect 390100 266970 390152 266976
rect 390664 264316 390692 267106
rect 391860 264330 391888 271254
rect 392032 269544 392084 269550
rect 392032 269486 392084 269492
rect 392044 267306 392072 269486
rect 392596 267714 392624 273634
rect 393332 271182 393360 278052
rect 393516 278038 394450 278066
rect 393320 271176 393372 271182
rect 393320 271118 393372 271124
rect 393516 270366 393544 278038
rect 395632 274514 395660 278052
rect 396092 278038 396842 278066
rect 397472 278038 398038 278066
rect 395620 274508 395672 274514
rect 395620 274450 395672 274456
rect 394332 274100 394384 274106
rect 394332 274042 394384 274048
rect 393964 271448 394016 271454
rect 393964 271390 394016 271396
rect 393504 270360 393556 270366
rect 393504 270302 393556 270308
rect 392584 267708 392636 267714
rect 392584 267650 392636 267656
rect 392032 267300 392084 267306
rect 392032 267242 392084 267248
rect 393136 267028 393188 267034
rect 393136 266970 393188 266976
rect 392308 266892 392360 266898
rect 392308 266834 392360 266840
rect 391506 264302 391888 264330
rect 392320 264316 392348 266834
rect 393148 264316 393176 266970
rect 393976 266898 394004 271390
rect 393964 266892 394016 266898
rect 393964 266834 394016 266840
rect 394344 264330 394372 274042
rect 395620 270496 395672 270502
rect 395620 270438 395672 270444
rect 394792 266756 394844 266762
rect 394792 266698 394844 266704
rect 393990 264302 394372 264330
rect 394804 264316 394832 266698
rect 395632 264316 395660 270438
rect 396092 270094 396120 278038
rect 397276 272536 397328 272542
rect 397276 272478 397328 272484
rect 396080 270088 396132 270094
rect 396080 270030 396132 270036
rect 397092 268524 397144 268530
rect 397092 268466 397144 268472
rect 397104 266762 397132 268466
rect 397092 266756 397144 266762
rect 397092 266698 397144 266704
rect 397288 266422 397316 272478
rect 397472 268394 397500 278038
rect 399220 273086 399248 278052
rect 400324 274378 400352 278052
rect 400508 278038 401534 278066
rect 401704 278038 402730 278066
rect 400312 274372 400364 274378
rect 400312 274314 400364 274320
rect 400036 273828 400088 273834
rect 400036 273770 400088 273776
rect 399208 273080 399260 273086
rect 399208 273022 399260 273028
rect 399852 270088 399904 270094
rect 399852 270030 399904 270036
rect 397460 268388 397512 268394
rect 397460 268330 397512 268336
rect 398104 267708 398156 267714
rect 398104 267650 398156 267656
rect 397460 266756 397512 266762
rect 397460 266698 397512 266704
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 396460 264316 396488 266358
rect 397472 266234 397500 266698
rect 397288 266206 397500 266234
rect 397288 264316 397316 266206
rect 398116 264316 398144 267650
rect 399864 267578 399892 270030
rect 399852 267572 399904 267578
rect 399852 267514 399904 267520
rect 400048 266422 400076 273770
rect 400508 269958 400536 278038
rect 401508 273216 401560 273222
rect 401508 273158 401560 273164
rect 400864 270360 400916 270366
rect 400864 270302 400916 270308
rect 400496 269952 400548 269958
rect 400496 269894 400548 269900
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 400036 266416 400088 266422
rect 400036 266358 400088 266364
rect 398944 264316 398972 266358
rect 400036 266280 400088 266286
rect 400036 266222 400088 266228
rect 400048 264330 400076 266222
rect 400876 264330 400904 270302
rect 401520 267734 401548 273158
rect 401704 269550 401732 278038
rect 403912 272814 403940 278052
rect 404372 278038 405122 278066
rect 405752 278038 406318 278066
rect 404176 274644 404228 274650
rect 404176 274586 404228 274592
rect 403900 272808 403952 272814
rect 403900 272750 403952 272756
rect 402612 271176 402664 271182
rect 402612 271118 402664 271124
rect 401876 269952 401928 269958
rect 401876 269894 401928 269900
rect 401692 269544 401744 269550
rect 401692 269486 401744 269492
rect 399786 264302 400076 264330
rect 400614 264302 400904 264330
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401888 267442 401916 269894
rect 401876 267436 401928 267442
rect 401876 267378 401928 267384
rect 402624 264330 402652 271118
rect 403256 268660 403308 268666
rect 403256 268602 403308 268608
rect 403072 267300 403124 267306
rect 403072 267242 403124 267248
rect 402270 264302 402652 264330
rect 403084 264316 403112 267242
rect 403268 266422 403296 268602
rect 403256 266416 403308 266422
rect 403256 266358 403308 266364
rect 404188 264330 404216 274586
rect 404372 269074 404400 278038
rect 405752 270230 405780 278038
rect 406844 272944 406896 272950
rect 406844 272886 406896 272892
rect 405740 270224 405792 270230
rect 405740 270166 405792 270172
rect 404544 269544 404596 269550
rect 404544 269486 404596 269492
rect 404360 269068 404412 269074
rect 404360 269010 404412 269016
rect 404556 266626 404584 269486
rect 405556 267436 405608 267442
rect 405556 267378 405608 267384
rect 404544 266620 404596 266626
rect 404544 266562 404596 266568
rect 404728 266620 404780 266626
rect 404728 266562 404780 266568
rect 403926 264302 404216 264330
rect 404740 264316 404768 266562
rect 405568 264316 405596 267378
rect 406856 264330 406884 272886
rect 407500 271862 407528 278052
rect 408512 278038 408618 278066
rect 408224 273080 408276 273086
rect 408224 273022 408276 273028
rect 407488 271856 407540 271862
rect 407488 271798 407540 271804
rect 407764 271856 407816 271862
rect 407764 271798 407816 271804
rect 407776 266762 407804 271798
rect 408040 268388 408092 268394
rect 408040 268330 408092 268336
rect 407764 266756 407816 266762
rect 407764 266698 407816 266704
rect 407212 266416 407264 266422
rect 407212 266358 407264 266364
rect 406410 264302 406884 264330
rect 407224 264316 407252 266358
rect 408052 264316 408080 268330
rect 408236 266422 408264 273022
rect 408512 269822 408540 278038
rect 409236 274508 409288 274514
rect 409236 274450 409288 274456
rect 408500 269816 408552 269822
rect 408500 269758 408552 269764
rect 408224 266416 408276 266422
rect 408224 266358 408276 266364
rect 409248 264330 409276 274450
rect 409800 273698 409828 278052
rect 410996 274242 411024 278052
rect 411824 278038 412206 278066
rect 412652 278038 413402 278066
rect 410984 274236 411036 274242
rect 410984 274178 411036 274184
rect 409788 273692 409840 273698
rect 409788 273634 409840 273640
rect 411824 271046 411852 278038
rect 412272 272808 412324 272814
rect 412272 272750 412324 272756
rect 411812 271040 411864 271046
rect 411812 270982 411864 270988
rect 409696 270224 409748 270230
rect 409696 270166 409748 270172
rect 408894 264302 409276 264330
rect 409708 264316 409736 270166
rect 410524 267572 410576 267578
rect 410524 267514 410576 267520
rect 410536 264316 410564 267514
rect 412284 266422 412312 272750
rect 412652 270094 412680 278038
rect 413468 274916 413520 274922
rect 413468 274858 413520 274864
rect 412640 270088 412692 270094
rect 412640 270030 412692 270036
rect 412456 269816 412508 269822
rect 412456 269758 412508 269764
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 411364 264316 411392 266358
rect 412468 264330 412496 269758
rect 412640 268116 412692 268122
rect 412640 268058 412692 268064
rect 412652 266626 412680 268058
rect 412640 266620 412692 266626
rect 412640 266562 412692 266568
rect 413480 264330 413508 274858
rect 413836 274372 413888 274378
rect 413836 274314 413888 274320
rect 412206 264302 412496 264330
rect 413034 264302 413508 264330
rect 413848 264316 413876 274314
rect 414584 272678 414612 278052
rect 415412 278038 415794 278066
rect 416792 278038 416898 278066
rect 414572 272672 414624 272678
rect 414572 272614 414624 272620
rect 414480 271040 414532 271046
rect 414480 270982 414532 270988
rect 414492 267714 414520 270982
rect 414664 270088 414716 270094
rect 414664 270030 414716 270036
rect 414480 267708 414532 267714
rect 414480 267650 414532 267656
rect 414676 264316 414704 270030
rect 415412 268938 415440 278038
rect 416412 275324 416464 275330
rect 416412 275266 416464 275272
rect 415400 268932 415452 268938
rect 415400 268874 415452 268880
rect 416424 266422 416452 275266
rect 416596 274236 416648 274242
rect 416596 274178 416648 274184
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 415504 264316 415532 266358
rect 416608 264330 416636 274178
rect 416792 269958 416820 278038
rect 418080 271726 418108 278052
rect 418264 278038 419290 278066
rect 418068 271720 418120 271726
rect 418068 271662 418120 271668
rect 417424 270904 417476 270910
rect 417424 270846 417476 270852
rect 416780 269952 416832 269958
rect 416780 269894 416832 269900
rect 417148 269952 417200 269958
rect 417148 269894 417200 269900
rect 416346 264302 416636 264330
rect 417160 264316 417188 269894
rect 417436 267170 417464 270846
rect 418264 269686 418292 278038
rect 420472 275466 420500 278052
rect 420460 275460 420512 275466
rect 420460 275402 420512 275408
rect 420644 275052 420696 275058
rect 420644 274994 420696 275000
rect 419172 272672 419224 272678
rect 419172 272614 419224 272620
rect 418252 269680 418304 269686
rect 418252 269622 418304 269628
rect 417424 267164 417476 267170
rect 417424 267106 417476 267112
rect 417976 267164 418028 267170
rect 417976 267106 418028 267112
rect 417988 264316 418016 267106
rect 419184 264330 419212 272614
rect 420184 271720 420236 271726
rect 420184 271662 420236 271668
rect 419632 268252 419684 268258
rect 419632 268194 419684 268200
rect 418830 264302 419212 264330
rect 419644 264316 419672 268194
rect 420196 267034 420224 271662
rect 420184 267028 420236 267034
rect 420184 266970 420236 266976
rect 420656 264330 420684 274994
rect 421668 273970 421696 278052
rect 421656 273964 421708 273970
rect 421656 273906 421708 273912
rect 421840 273964 421892 273970
rect 421840 273906 421892 273912
rect 421852 267734 421880 273906
rect 422864 271590 422892 278052
rect 423692 278038 423982 278066
rect 423404 275460 423456 275466
rect 423404 275402 423456 275408
rect 422852 271584 422904 271590
rect 422852 271526 422904 271532
rect 422944 270632 422996 270638
rect 422944 270574 422996 270580
rect 422116 269680 422168 269686
rect 422116 269622 422168 269628
rect 421760 267706 421880 267734
rect 421760 264330 421788 267706
rect 420486 264302 420684 264330
rect 421314 264302 421788 264330
rect 422128 264316 422156 269622
rect 422956 267306 422984 270574
rect 422944 267300 422996 267306
rect 422944 267242 422996 267248
rect 423416 264330 423444 275402
rect 423692 269550 423720 278038
rect 425164 272406 425192 278052
rect 425348 278038 426374 278066
rect 425152 272400 425204 272406
rect 425152 272342 425204 272348
rect 423680 269544 423732 269550
rect 423680 269486 423732 269492
rect 423956 269272 424008 269278
rect 423956 269214 424008 269220
rect 423772 267708 423824 267714
rect 423772 267650 423824 267656
rect 422970 264302 423444 264330
rect 423784 264316 423812 267650
rect 423968 267442 423996 269214
rect 425348 268802 425376 278038
rect 427084 275188 427136 275194
rect 427084 275130 427136 275136
rect 426348 272128 426400 272134
rect 426348 272070 426400 272076
rect 425336 268796 425388 268802
rect 425336 268738 425388 268744
rect 426360 267734 426388 272070
rect 426268 267706 426388 267734
rect 423956 267436 424008 267442
rect 423956 267378 424008 267384
rect 424600 267300 424652 267306
rect 424600 267242 424652 267248
rect 424612 264316 424640 267242
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426268 264316 426296 267706
rect 427096 266422 427124 275130
rect 427556 270910 427584 278052
rect 428752 271318 428780 278052
rect 429948 271454 429976 278052
rect 430212 275596 430264 275602
rect 430212 275538 430264 275544
rect 429936 271448 429988 271454
rect 429936 271390 429988 271396
rect 428740 271312 428792 271318
rect 428740 271254 428792 271260
rect 427544 270904 427596 270910
rect 427544 270846 427596 270852
rect 427452 270768 427504 270774
rect 427452 270710 427504 270716
rect 427084 266416 427136 266422
rect 427084 266358 427136 266364
rect 427464 264330 427492 270710
rect 429108 269408 429160 269414
rect 429108 269350 429160 269356
rect 429120 267578 429148 269350
rect 429108 267572 429160 267578
rect 429108 267514 429160 267520
rect 427912 266892 427964 266898
rect 427912 266834 427964 266840
rect 427110 264302 427492 264330
rect 427924 264316 427952 266834
rect 428740 266756 428792 266762
rect 428740 266698 428792 266704
rect 428752 264316 428780 266698
rect 429568 266416 429620 266422
rect 429568 266358 429620 266364
rect 429580 264316 429608 266358
rect 430224 264330 430252 275538
rect 431144 271726 431172 278052
rect 432248 274106 432276 278052
rect 433444 277394 433472 278052
rect 433352 277366 433472 277394
rect 433628 278038 434654 278066
rect 432236 274100 432288 274106
rect 432236 274042 432288 274048
rect 432604 274100 432656 274106
rect 432604 274042 432656 274048
rect 431132 271720 431184 271726
rect 431132 271662 431184 271668
rect 430396 270904 430448 270910
rect 430396 270846 430448 270852
rect 430408 266422 430436 270846
rect 432236 269544 432288 269550
rect 432236 269486 432288 269492
rect 432052 267436 432104 267442
rect 432052 267378 432104 267384
rect 431224 267028 431276 267034
rect 431224 266970 431276 266976
rect 430396 266416 430448 266422
rect 430396 266358 430448 266364
rect 430224 264302 430422 264330
rect 431236 264316 431264 266970
rect 432064 264316 432092 267378
rect 432248 267170 432276 269486
rect 432236 267164 432288 267170
rect 432236 267106 432288 267112
rect 432616 267034 432644 274042
rect 433352 268530 433380 277366
rect 433628 270502 433656 278038
rect 435640 275732 435692 275738
rect 435640 275674 435692 275680
rect 434628 271720 434680 271726
rect 434628 271662 434680 271668
rect 433616 270496 433668 270502
rect 433616 270438 433668 270444
rect 433708 268932 433760 268938
rect 433708 268874 433760 268880
rect 433340 268524 433392 268530
rect 433340 268466 433392 268472
rect 432880 267164 432932 267170
rect 432880 267106 432932 267112
rect 432604 267028 432656 267034
rect 432604 266970 432656 266976
rect 432892 264316 432920 267106
rect 433720 264316 433748 268874
rect 434640 267734 434668 271662
rect 434548 267706 434668 267734
rect 434548 264316 434576 267706
rect 435652 264330 435680 275674
rect 435836 272542 435864 278052
rect 435824 272536 435876 272542
rect 435824 272478 435876 272484
rect 437032 271862 437060 278052
rect 438136 278038 438242 278066
rect 437020 271856 437072 271862
rect 437020 271798 437072 271804
rect 437204 271856 437256 271862
rect 437204 271798 437256 271804
rect 436192 269068 436244 269074
rect 436192 269010 436244 269016
rect 435390 264302 435680 264330
rect 436204 264316 436232 269010
rect 437216 264330 437244 271798
rect 438136 271046 438164 278038
rect 439332 273834 439360 278052
rect 440252 278038 440542 278066
rect 439320 273828 439372 273834
rect 439320 273770 439372 273776
rect 438768 272536 438820 272542
rect 438768 272478 438820 272484
rect 438124 271040 438176 271046
rect 438124 270982 438176 270988
rect 438308 271040 438360 271046
rect 438308 270982 438360 270988
rect 438320 264330 438348 270982
rect 438780 267734 438808 272478
rect 439964 271584 440016 271590
rect 439964 271526 440016 271532
rect 437046 264302 437244 264330
rect 437874 264302 438348 264330
rect 438688 267706 438808 267734
rect 438688 264316 438716 267706
rect 439976 264330 440004 271526
rect 440252 268666 440280 278038
rect 441724 277394 441752 278052
rect 441632 277366 441752 277394
rect 440884 273692 440936 273698
rect 440884 273634 440936 273640
rect 440240 268660 440292 268666
rect 440240 268602 440292 268608
rect 440896 267714 440924 273634
rect 441632 270366 441660 277366
rect 442264 273828 442316 273834
rect 442264 273770 442316 273776
rect 441620 270360 441672 270366
rect 441620 270302 441672 270308
rect 441160 268796 441212 268802
rect 441160 268738 441212 268744
rect 440884 267708 440936 267714
rect 440884 267650 440936 267656
rect 440332 266756 440384 266762
rect 440332 266698 440384 266704
rect 439530 264302 440004 264330
rect 440344 264316 440372 266698
rect 441172 264316 441200 268738
rect 442276 266626 442304 273770
rect 442920 273222 442948 278052
rect 442908 273216 442960 273222
rect 442908 273158 442960 273164
rect 442908 271448 442960 271454
rect 442908 271390 442960 271396
rect 442724 267708 442776 267714
rect 442724 267650 442776 267656
rect 442264 266620 442316 266626
rect 442264 266562 442316 266568
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 267650
rect 442920 266422 442948 271390
rect 444116 271182 444144 278052
rect 445024 275868 445076 275874
rect 445024 275810 445076 275816
rect 444104 271176 444156 271182
rect 444104 271118 444156 271124
rect 443644 268660 443696 268666
rect 443644 268602 443696 268608
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 442736 264302 442842 264330
rect 443656 264316 443684 268602
rect 445036 266762 445064 275810
rect 445312 270638 445340 278052
rect 446508 274650 446536 278052
rect 447152 278038 447626 278066
rect 448532 278038 448822 278066
rect 446496 274644 446548 274650
rect 446496 274586 446548 274592
rect 446404 273556 446456 273562
rect 446404 273498 446456 273504
rect 445668 271312 445720 271318
rect 445668 271254 445720 271260
rect 445300 270632 445352 270638
rect 445300 270574 445352 270580
rect 445300 267572 445352 267578
rect 445300 267514 445352 267520
rect 445024 266756 445076 266762
rect 445024 266698 445076 266704
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 444484 264316 444512 266358
rect 445312 264316 445340 267514
rect 445680 266422 445708 271254
rect 446416 267306 446444 273498
rect 446956 272264 447008 272270
rect 446956 272206 447008 272212
rect 446404 267300 446456 267306
rect 446404 267242 446456 267248
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446128 266416 446180 266422
rect 446128 266358 446180 266364
rect 446140 264316 446168 266358
rect 446968 264316 446996 272206
rect 447152 268122 447180 278038
rect 447784 271992 447836 271998
rect 447784 271934 447836 271940
rect 447140 268116 447192 268122
rect 447140 268058 447192 268064
rect 447796 266422 447824 271934
rect 448532 269278 448560 278038
rect 450004 272950 450032 278052
rect 450832 278038 451214 278066
rect 451384 278038 452410 278066
rect 450544 274644 450596 274650
rect 450544 274586 450596 274592
rect 449992 272944 450044 272950
rect 449992 272886 450044 272892
rect 449808 272400 449860 272406
rect 449808 272342 449860 272348
rect 448520 269272 448572 269278
rect 448520 269214 448572 269220
rect 448612 268524 448664 268530
rect 448612 268466 448664 268472
rect 448152 267300 448204 267306
rect 448152 267242 448204 267248
rect 447784 266416 447836 266422
rect 447784 266358 447836 266364
rect 448164 264330 448192 267242
rect 447810 264302 448192 264330
rect 448624 264316 448652 268466
rect 449820 264330 449848 272342
rect 450556 267034 450584 274586
rect 450832 273086 450860 278038
rect 451188 273216 451240 273222
rect 451188 273158 451240 273164
rect 450820 273080 450872 273086
rect 450820 273022 450872 273028
rect 451200 267734 451228 273158
rect 451384 268394 451412 278038
rect 453592 274514 453620 278052
rect 454052 278038 454710 278066
rect 455432 278038 455906 278066
rect 453580 274508 453632 274514
rect 453580 274450 453632 274456
rect 453764 274508 453816 274514
rect 453764 274450 453816 274456
rect 453776 273358 453804 274450
rect 453304 273352 453356 273358
rect 453304 273294 453356 273300
rect 453764 273352 453816 273358
rect 453764 273294 453816 273300
rect 452292 273080 452344 273086
rect 452292 273022 452344 273028
rect 451372 268388 451424 268394
rect 451372 268330 451424 268336
rect 451108 267706 451228 267734
rect 450544 267028 450596 267034
rect 450544 266970 450596 266976
rect 450268 266892 450320 266898
rect 450268 266834 450320 266840
rect 449466 264302 449848 264330
rect 450280 264316 450308 266834
rect 451108 264316 451136 267706
rect 452304 264330 452332 273022
rect 453316 267442 453344 273294
rect 453580 270496 453632 270502
rect 453580 270438 453632 270444
rect 453304 267436 453356 267442
rect 453304 267378 453356 267384
rect 452752 266620 452804 266626
rect 452752 266562 452804 266568
rect 451950 264302 452332 264330
rect 452764 264316 452792 266562
rect 453592 264316 453620 270438
rect 454052 270230 454080 278038
rect 454408 276004 454460 276010
rect 454408 275946 454460 275952
rect 454420 275738 454448 275946
rect 454408 275732 454460 275738
rect 454408 275674 454460 275680
rect 455236 272944 455288 272950
rect 455236 272886 455288 272892
rect 454040 270224 454092 270230
rect 454040 270166 454092 270172
rect 455052 267028 455104 267034
rect 455052 266970 455104 266976
rect 454408 266416 454460 266422
rect 454408 266358 454460 266364
rect 454420 264316 454448 266358
rect 455064 264330 455092 266970
rect 455248 266422 455276 272886
rect 455432 269414 455460 278038
rect 457088 272814 457116 278052
rect 457444 276004 457496 276010
rect 457444 275946 457496 275952
rect 457076 272808 457128 272814
rect 457076 272750 457128 272756
rect 456064 270360 456116 270366
rect 456064 270302 456116 270308
rect 455420 269408 455472 269414
rect 455420 269350 455472 269356
rect 455236 266416 455288 266422
rect 455236 266358 455288 266364
rect 455064 264302 455262 264330
rect 456076 264316 456104 270302
rect 457456 267306 457484 275946
rect 458088 273080 458140 273086
rect 458088 273022 458140 273028
rect 457444 267300 457496 267306
rect 457444 267242 457496 267248
rect 457720 266756 457772 266762
rect 457720 266698 457772 266704
rect 456892 266416 456944 266422
rect 456892 266358 456944 266364
rect 456904 264316 456932 266358
rect 457732 264316 457760 266698
rect 458100 266422 458128 273022
rect 458284 269822 458312 278052
rect 459480 274922 459508 278052
rect 459468 274916 459520 274922
rect 459468 274858 459520 274864
rect 460676 274378 460704 278052
rect 460952 278038 461886 278066
rect 460664 274372 460716 274378
rect 460664 274314 460716 274320
rect 460020 273420 460072 273426
rect 460020 273362 460072 273368
rect 459468 271176 459520 271182
rect 459468 271118 459520 271124
rect 458548 270224 458600 270230
rect 458548 270166 458600 270172
rect 458272 269816 458324 269822
rect 458272 269758 458324 269764
rect 458088 266416 458140 266422
rect 458088 266358 458140 266364
rect 458560 264316 458588 270166
rect 459480 267734 459508 271118
rect 459388 267706 459508 267734
rect 459388 264316 459416 267706
rect 460032 267170 460060 273362
rect 460952 270094 460980 278038
rect 462976 275330 463004 278052
rect 462964 275324 463016 275330
rect 462964 275266 463016 275272
rect 463148 275324 463200 275330
rect 463148 275266 463200 275272
rect 462226 272368 462282 272377
rect 462226 272303 462282 272312
rect 460940 270088 460992 270094
rect 460940 270030 460992 270036
rect 461400 270088 461452 270094
rect 461400 270030 461452 270036
rect 460204 267436 460256 267442
rect 460204 267378 460256 267384
rect 460020 267164 460072 267170
rect 460020 267106 460072 267112
rect 460216 264316 460244 267378
rect 461412 264330 461440 270030
rect 462240 264330 462268 272303
rect 463160 264330 463188 275266
rect 464172 274242 464200 278052
rect 465092 278038 465382 278066
rect 464160 274236 464212 274242
rect 464160 274178 464212 274184
rect 465092 269958 465120 278038
rect 466564 277394 466592 278052
rect 466472 277366 466592 277394
rect 467392 278038 467774 278066
rect 467944 278038 468970 278066
rect 465724 274372 465776 274378
rect 465724 274314 465776 274320
rect 465736 273426 465764 274314
rect 465724 273420 465776 273426
rect 465724 273362 465776 273368
rect 465540 273080 465592 273086
rect 465540 273022 465592 273028
rect 465724 273080 465776 273086
rect 465724 273022 465776 273028
rect 465552 272678 465580 273022
rect 465736 272814 465764 273022
rect 465724 272808 465776 272814
rect 465724 272750 465776 272756
rect 465356 272672 465408 272678
rect 465356 272614 465408 272620
rect 465540 272672 465592 272678
rect 466092 272672 466144 272678
rect 465540 272614 465592 272620
rect 465736 272620 466092 272626
rect 465736 272614 466144 272620
rect 465368 272490 465396 272614
rect 465736 272598 466132 272614
rect 465736 272490 465764 272598
rect 465368 272462 465764 272490
rect 465080 269952 465132 269958
rect 465080 269894 465132 269900
rect 463516 269816 463568 269822
rect 463516 269758 463568 269764
rect 461058 264302 461440 264330
rect 461886 264302 462268 264330
rect 462714 264302 463188 264330
rect 463528 264316 463556 269758
rect 466472 269550 466500 277366
rect 467392 272678 467420 278038
rect 467564 273420 467616 273426
rect 467564 273362 467616 273368
rect 467380 272672 467432 272678
rect 467380 272614 467432 272620
rect 466460 269544 466512 269550
rect 466460 269486 466512 269492
rect 466000 269408 466052 269414
rect 466000 269350 466052 269356
rect 464344 268388 464396 268394
rect 464344 268330 464396 268336
rect 464356 264316 464384 268330
rect 465172 267164 465224 267170
rect 465172 267106 465224 267112
rect 465184 264316 465212 267106
rect 466012 264316 466040 269350
rect 466828 266416 466880 266422
rect 466828 266358 466880 266364
rect 466840 264316 466868 266358
rect 467576 264330 467604 273362
rect 467748 272672 467800 272678
rect 467748 272614 467800 272620
rect 467760 266422 467788 272614
rect 467944 268258 467972 278038
rect 470152 275058 470180 278052
rect 470140 275052 470192 275058
rect 470140 274994 470192 275000
rect 469864 274780 469916 274786
rect 469864 274722 469916 274728
rect 468484 269952 468536 269958
rect 468484 269894 468536 269900
rect 467932 268252 467984 268258
rect 467932 268194 467984 268200
rect 467748 266416 467800 266422
rect 467748 266358 467800 266364
rect 467576 264302 467682 264330
rect 468496 264316 468524 269894
rect 469876 266626 469904 274722
rect 471256 273970 471284 278052
rect 471992 278038 472466 278066
rect 473372 278038 473662 278066
rect 471612 276276 471664 276282
rect 471612 276218 471664 276224
rect 471244 273964 471296 273970
rect 471244 273906 471296 273912
rect 470416 272672 470468 272678
rect 470414 272640 470416 272649
rect 470600 272672 470652 272678
rect 470468 272640 470470 272649
rect 470414 272575 470470 272584
rect 470598 272640 470600 272649
rect 470652 272640 470654 272649
rect 470598 272575 470654 272584
rect 470428 272462 470824 272490
rect 470428 272377 470456 272462
rect 470414 272368 470470 272377
rect 470414 272303 470470 272312
rect 470796 272134 470824 272462
rect 470554 272128 470606 272134
rect 470784 272128 470836 272134
rect 470606 272076 470640 272082
rect 470554 272070 470640 272076
rect 470784 272070 470836 272076
rect 470566 272054 470640 272070
rect 470612 271969 470640 272054
rect 470598 271960 470654 271969
rect 470598 271895 470654 271904
rect 470968 269272 471020 269278
rect 470968 269214 471020 269220
rect 470140 267300 470192 267306
rect 470140 267242 470192 267248
rect 469864 266620 469916 266626
rect 469864 266562 469916 266568
rect 469312 265124 469364 265130
rect 469312 265066 469364 265072
rect 469324 264316 469352 265066
rect 470152 264316 470180 267242
rect 470980 264316 471008 269214
rect 471624 264330 471652 276218
rect 471992 269686 472020 278038
rect 473372 275466 473400 278038
rect 473360 275460 473412 275466
rect 473360 275402 473412 275408
rect 473360 274916 473412 274922
rect 473360 274858 473412 274864
rect 473372 269686 473400 274858
rect 474648 274236 474700 274242
rect 474648 274178 474700 274184
rect 471980 269680 472032 269686
rect 471980 269622 472032 269628
rect 472624 269680 472676 269686
rect 472624 269622 472676 269628
rect 473360 269680 473412 269686
rect 473360 269622 473412 269628
rect 471624 264302 471822 264330
rect 472636 264316 472664 269622
rect 474280 269408 474332 269414
rect 474280 269350 474332 269356
rect 473452 266416 473504 266422
rect 473452 266358 473504 266364
rect 473464 264316 473492 266358
rect 474292 264316 474320 269350
rect 474660 266422 474688 274178
rect 474844 273698 474872 278052
rect 476040 277394 476068 278052
rect 475948 277366 476068 277394
rect 475384 275868 475436 275874
rect 475384 275810 475436 275816
rect 475396 275466 475424 275810
rect 475384 275460 475436 275466
rect 475384 275402 475436 275408
rect 475752 273964 475804 273970
rect 475752 273906 475804 273912
rect 474832 273692 474884 273698
rect 474832 273634 474884 273640
rect 474648 266416 474700 266422
rect 474648 266358 474700 266364
rect 475108 265260 475160 265266
rect 475108 265202 475160 265208
rect 475120 264316 475148 265202
rect 475764 264330 475792 273906
rect 475948 273562 475976 277366
rect 477040 276548 477092 276554
rect 477040 276490 477092 276496
rect 476120 275052 476172 275058
rect 476120 274994 476172 275000
rect 475936 273556 475988 273562
rect 475936 273498 475988 273504
rect 476132 273426 476160 274994
rect 476120 273420 476172 273426
rect 476120 273362 476172 273368
rect 477052 264330 477080 276490
rect 477236 275194 477264 278052
rect 478064 278038 478354 278066
rect 479168 278038 479550 278066
rect 477224 275188 477276 275194
rect 477224 275130 477276 275136
rect 478064 271969 478092 278038
rect 478512 276412 478564 276418
rect 478512 276354 478564 276360
rect 478050 271960 478106 271969
rect 478050 271895 478106 271904
rect 478524 266422 478552 276354
rect 478696 273420 478748 273426
rect 478696 273362 478748 273368
rect 477592 266416 477644 266422
rect 477592 266358 477644 266364
rect 478512 266416 478564 266422
rect 478512 266358 478564 266364
rect 475764 264302 475962 264330
rect 476790 264302 477080 264330
rect 477604 264316 477632 266358
rect 478708 264330 478736 273362
rect 479168 270774 479196 278038
rect 479524 275868 479576 275874
rect 479524 275810 479576 275816
rect 479156 270768 479208 270774
rect 479156 270710 479208 270716
rect 479536 266762 479564 275810
rect 480732 274650 480760 278052
rect 480720 274644 480772 274650
rect 480720 274586 480772 274592
rect 481928 273834 481956 278052
rect 482836 277364 482888 277370
rect 482836 277306 482888 277312
rect 481916 273828 481968 273834
rect 481916 273770 481968 273776
rect 481364 273692 481416 273698
rect 481364 273634 481416 273640
rect 479524 266756 479576 266762
rect 479524 266698 479576 266704
rect 480076 265532 480128 265538
rect 480076 265474 480128 265480
rect 479248 265396 479300 265402
rect 479248 265338 479300 265344
rect 478446 264302 478736 264330
rect 479260 264316 479288 265338
rect 480088 264316 480116 265474
rect 481376 264330 481404 273634
rect 482560 266552 482612 266558
rect 482560 266494 482612 266500
rect 481732 266416 481784 266422
rect 481732 266358 481784 266364
rect 480930 264302 481404 264330
rect 481744 264316 481772 266358
rect 482572 264316 482600 266494
rect 482848 266422 482876 277306
rect 483124 270910 483152 278052
rect 484320 275602 484348 278052
rect 484308 275596 484360 275602
rect 484308 275538 484360 275544
rect 485044 275460 485096 275466
rect 485044 275402 485096 275408
rect 485228 275460 485280 275466
rect 485228 275402 485280 275408
rect 485056 275194 485084 275402
rect 485044 275188 485096 275194
rect 485044 275130 485096 275136
rect 485240 275058 485268 275402
rect 485228 275052 485280 275058
rect 485228 274994 485280 275000
rect 485516 274106 485544 278052
rect 485688 277228 485740 277234
rect 485688 277170 485740 277176
rect 485504 274100 485556 274106
rect 485504 274042 485556 274048
rect 484308 273556 484360 273562
rect 484308 273498 484360 273504
rect 483112 270904 483164 270910
rect 483112 270846 483164 270852
rect 484320 266422 484348 273498
rect 485228 271720 485280 271726
rect 485228 271662 485280 271668
rect 485412 271720 485464 271726
rect 485412 271662 485464 271668
rect 485240 271046 485268 271662
rect 485228 271040 485280 271046
rect 485228 270982 485280 270988
rect 485424 269770 485452 271662
rect 485056 269742 485452 269770
rect 485056 266558 485084 269742
rect 485700 267734 485728 277170
rect 486620 274514 486648 278052
rect 486608 274508 486660 274514
rect 486608 274450 486660 274456
rect 487816 274378 487844 278052
rect 488552 278038 489026 278066
rect 488356 274644 488408 274650
rect 488356 274586 488408 274592
rect 487804 274372 487856 274378
rect 487804 274314 487856 274320
rect 487068 273828 487120 273834
rect 487068 273770 487120 273776
rect 486884 270768 486936 270774
rect 486884 270710 486936 270716
rect 485424 267706 485728 267734
rect 485044 266552 485096 266558
rect 485044 266494 485096 266500
rect 482836 266416 482888 266422
rect 482836 266358 482888 266364
rect 483388 266416 483440 266422
rect 483388 266358 483440 266364
rect 484308 266416 484360 266422
rect 484308 266358 484360 266364
rect 483400 264316 483428 266358
rect 484216 266280 484268 266286
rect 484216 266222 484268 266228
rect 484228 264316 484256 266222
rect 485424 264330 485452 267706
rect 485872 266416 485924 266422
rect 485872 266358 485924 266364
rect 485070 264302 485452 264330
rect 485884 264316 485912 266358
rect 486896 264330 486924 270710
rect 487080 266422 487108 273770
rect 487068 266416 487120 266422
rect 487068 266358 487120 266364
rect 487528 266212 487580 266218
rect 487528 266154 487580 266160
rect 486726 264302 486924 264330
rect 487540 264316 487568 266154
rect 488368 264316 488396 274586
rect 488552 268938 488580 278038
rect 489918 272776 489974 272785
rect 489918 272711 489974 272720
rect 489932 272626 489960 272711
rect 489886 272598 489960 272626
rect 489886 272542 489914 272598
rect 489874 272536 489926 272542
rect 489874 272478 489926 272484
rect 490012 272536 490064 272542
rect 490012 272478 490064 272484
rect 490024 272218 490052 272478
rect 489886 272190 490052 272218
rect 489886 272134 489914 272190
rect 489874 272128 489926 272134
rect 489874 272070 489926 272076
rect 490012 272128 490064 272134
rect 490012 272070 490064 272076
rect 490024 271726 490052 272070
rect 490012 271720 490064 271726
rect 490012 271662 490064 271668
rect 490208 271046 490236 278052
rect 491404 275194 491432 278052
rect 491772 278038 492614 278066
rect 491392 275188 491444 275194
rect 491392 275130 491444 275136
rect 491208 274100 491260 274106
rect 491208 274042 491260 274048
rect 490196 271040 490248 271046
rect 490196 270982 490248 270988
rect 489644 270632 489696 270638
rect 489644 270574 489696 270580
rect 488540 268932 488592 268938
rect 488540 268874 488592 268880
rect 489656 264330 489684 270574
rect 490012 266756 490064 266762
rect 490012 266698 490064 266704
rect 489210 264302 489684 264330
rect 490024 264316 490052 266698
rect 491220 264330 491248 274042
rect 491772 269074 491800 278038
rect 493324 275188 493376 275194
rect 493324 275130 493376 275136
rect 492404 275052 492456 275058
rect 492404 274994 492456 275000
rect 492416 270910 492444 274994
rect 492404 270904 492456 270910
rect 492404 270846 492456 270852
rect 492588 270904 492640 270910
rect 492588 270846 492640 270852
rect 491760 269068 491812 269074
rect 491760 269010 491812 269016
rect 492600 266490 492628 270846
rect 493336 267714 493364 275130
rect 493704 271862 493732 278052
rect 494900 275058 494928 278052
rect 495728 278038 496110 278066
rect 495072 277092 495124 277098
rect 495072 277034 495124 277040
rect 494888 275052 494940 275058
rect 494888 274994 494940 275000
rect 493692 271856 493744 271862
rect 493692 271798 493744 271804
rect 493600 268252 493652 268258
rect 493600 268194 493652 268200
rect 493324 267708 493376 267714
rect 493324 267650 493376 267656
rect 491668 266484 491720 266490
rect 491668 266426 491720 266432
rect 492588 266484 492640 266490
rect 492588 266426 492640 266432
rect 490866 264302 491248 264330
rect 491680 264316 491708 266426
rect 492496 266076 492548 266082
rect 492496 266018 492548 266024
rect 492508 264316 492536 266018
rect 493612 264330 493640 268194
rect 495084 267734 495112 277034
rect 495728 272785 495756 278038
rect 495714 272776 495770 272785
rect 495714 272711 495770 272720
rect 496544 271856 496596 271862
rect 496544 271798 496596 271804
rect 495256 271040 495308 271046
rect 495256 270982 495308 270988
rect 494992 267706 495112 267734
rect 494152 266484 494204 266490
rect 494152 266426 494204 266432
rect 493350 264302 493640 264330
rect 494164 264316 494192 266426
rect 494992 264316 495020 267706
rect 495268 266490 495296 270982
rect 495808 268116 495860 268122
rect 495808 268058 495860 268064
rect 495256 266484 495308 266490
rect 495256 266426 495308 266432
rect 495820 264316 495848 268058
rect 496556 264330 496584 271798
rect 497292 271590 497320 278052
rect 498488 275738 498516 278052
rect 499684 277394 499712 278052
rect 499592 277366 499712 277394
rect 498476 275732 498528 275738
rect 498476 275674 498528 275680
rect 497464 275188 497516 275194
rect 497464 275130 497516 275136
rect 497280 271584 497332 271590
rect 497280 271526 497332 271532
rect 497476 267578 497504 275130
rect 499304 271584 499356 271590
rect 499304 271526 499356 271532
rect 498292 269068 498344 269074
rect 498292 269010 498344 269016
rect 497832 267708 497884 267714
rect 497832 267650 497884 267656
rect 497464 267572 497516 267578
rect 497464 267514 497516 267520
rect 497844 264330 497872 267650
rect 496556 264302 496662 264330
rect 497490 264302 497872 264330
rect 498304 264316 498332 269010
rect 499316 264330 499344 271526
rect 499592 268802 499620 277366
rect 500880 271454 500908 278052
rect 501604 275596 501656 275602
rect 501604 275538 501656 275544
rect 500868 271448 500920 271454
rect 500868 271390 500920 271396
rect 500776 268932 500828 268938
rect 500776 268874 500828 268880
rect 499580 268796 499632 268802
rect 499580 268738 499632 268744
rect 499948 266484 500000 266490
rect 499948 266426 500000 266432
rect 499146 264302 499344 264330
rect 499960 264316 499988 266426
rect 500788 264316 500816 268874
rect 501616 266626 501644 275538
rect 501984 275058 502012 278052
rect 502352 278038 503194 278066
rect 501972 275052 502024 275058
rect 501972 274994 502024 275000
rect 501972 271720 502024 271726
rect 501972 271662 502024 271668
rect 501604 266620 501656 266626
rect 501604 266562 501656 266568
rect 501984 264330 502012 271662
rect 502352 268666 502380 278038
rect 503444 275052 503496 275058
rect 503444 274994 503496 275000
rect 503260 268796 503312 268802
rect 503260 268738 503312 268744
rect 502340 268660 502392 268666
rect 502340 268602 502392 268608
rect 502432 266484 502484 266490
rect 502432 266426 502484 266432
rect 501630 264302 502012 264330
rect 502444 264316 502472 266426
rect 503272 264316 503300 268738
rect 503456 266490 503484 274994
rect 504376 271318 504404 278052
rect 505572 275194 505600 278052
rect 505560 275188 505612 275194
rect 505560 275130 505612 275136
rect 506768 271998 506796 278052
rect 507964 277394 507992 278052
rect 507964 277366 508084 277394
rect 507860 275732 507912 275738
rect 507860 275674 507912 275680
rect 507492 275188 507544 275194
rect 507492 275130 507544 275136
rect 506756 271992 506808 271998
rect 506756 271934 506808 271940
rect 507124 271992 507176 271998
rect 507124 271934 507176 271940
rect 505008 271448 505060 271454
rect 505008 271390 505060 271396
rect 504364 271312 504416 271318
rect 504364 271254 504416 271260
rect 504824 266892 504876 266898
rect 504824 266834 504876 266840
rect 503444 266484 503496 266490
rect 503444 266426 503496 266432
rect 504088 266484 504140 266490
rect 504088 266426 504140 266432
rect 504100 264316 504128 266426
rect 504836 264330 504864 266834
rect 505020 266490 505048 271390
rect 505744 268660 505796 268666
rect 505744 268602 505796 268608
rect 505008 266484 505060 266490
rect 505008 266426 505060 266432
rect 504836 264302 504942 264330
rect 505756 264316 505784 268602
rect 507136 266762 507164 271934
rect 507504 267734 507532 275130
rect 507872 274242 507900 275674
rect 507860 274236 507912 274242
rect 507860 274178 507912 274184
rect 508056 272270 508084 277366
rect 509068 276010 509096 278052
rect 509252 278038 510278 278066
rect 509056 276004 509108 276010
rect 509056 275946 509108 275952
rect 508596 274372 508648 274378
rect 508596 274314 508648 274320
rect 508044 272264 508096 272270
rect 508044 272206 508096 272212
rect 507676 271312 507728 271318
rect 507676 271254 507728 271260
rect 507412 267706 507532 267734
rect 507124 266756 507176 266762
rect 507124 266698 507176 266704
rect 506572 266484 506624 266490
rect 506572 266426 506624 266432
rect 506584 264316 506612 266426
rect 507412 264316 507440 267706
rect 507688 266490 507716 271254
rect 507676 266484 507728 266490
rect 507676 266426 507728 266432
rect 508608 264330 508636 274314
rect 509056 269544 509108 269550
rect 509056 269486 509108 269492
rect 508254 264302 508636 264330
rect 509068 264316 509096 269486
rect 509252 268530 509280 278038
rect 511460 272406 511488 278052
rect 511632 276956 511684 276962
rect 511632 276898 511684 276904
rect 511448 272400 511500 272406
rect 511448 272342 511500 272348
rect 509240 268524 509292 268530
rect 509240 268466 509292 268472
rect 511644 267734 511672 276898
rect 512656 275602 512684 278052
rect 512644 275596 512696 275602
rect 512644 275538 512696 275544
rect 511816 274236 511868 274242
rect 511816 274178 511868 274184
rect 511552 267706 511672 267734
rect 509884 266756 509936 266762
rect 509884 266698 509936 266704
rect 509896 264316 509924 266698
rect 510712 266620 510764 266626
rect 510712 266562 510764 266568
rect 510724 264316 510752 266562
rect 511552 264316 511580 267706
rect 511828 266626 511856 274178
rect 513852 273222 513880 278052
rect 514484 276820 514536 276826
rect 514484 276762 514536 276768
rect 513840 273216 513892 273222
rect 513840 273158 513892 273164
rect 514024 273216 514076 273222
rect 514024 273158 514076 273164
rect 514036 272406 514064 273158
rect 512644 272400 512696 272406
rect 512644 272342 512696 272348
rect 514024 272400 514076 272406
rect 514024 272342 514076 272348
rect 512656 267034 512684 272342
rect 513196 268524 513248 268530
rect 513196 268466 513248 268472
rect 512644 267028 512696 267034
rect 512644 266970 512696 266976
rect 511816 266620 511868 266626
rect 511816 266562 511868 266568
rect 512368 265940 512420 265946
rect 512368 265882 512420 265888
rect 512380 264316 512408 265882
rect 513208 264316 513236 268466
rect 513932 266892 513984 266898
rect 513932 266834 513984 266840
rect 513944 266626 513972 266834
rect 513932 266620 513984 266626
rect 513932 266562 513984 266568
rect 514496 264330 514524 276762
rect 515048 272950 515076 278052
rect 515404 275596 515456 275602
rect 515404 275538 515456 275544
rect 515036 272944 515088 272950
rect 515036 272886 515088 272892
rect 514852 267572 514904 267578
rect 514852 267514 514904 267520
rect 514050 264302 514524 264330
rect 514864 264316 514892 267514
rect 515416 267442 515444 275538
rect 516244 274786 516272 278052
rect 516796 278038 517362 278066
rect 516232 274780 516284 274786
rect 516232 274722 516284 274728
rect 516796 270502 516824 278038
rect 517152 276004 517204 276010
rect 517152 275946 517204 275952
rect 516784 270496 516836 270502
rect 516784 270438 516836 270444
rect 515404 267436 515456 267442
rect 515404 267378 515456 267384
rect 516508 266756 516560 266762
rect 516508 266698 516560 266704
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266698
rect 517164 264330 517192 275946
rect 518544 273086 518572 278052
rect 518716 276684 518768 276690
rect 518716 276626 518768 276632
rect 518532 273080 518584 273086
rect 518532 273022 518584 273028
rect 517336 272400 517388 272406
rect 517336 272342 517388 272348
rect 517348 266762 517376 272342
rect 517520 270496 517572 270502
rect 517520 270438 517572 270444
rect 517532 267714 517560 270438
rect 518728 267734 518756 276626
rect 519740 273222 519768 278052
rect 520292 278038 520950 278066
rect 519728 273216 519780 273222
rect 519728 273158 519780 273164
rect 520096 272264 520148 272270
rect 520096 272206 520148 272212
rect 517520 267708 517572 267714
rect 517520 267650 517572 267656
rect 518544 267706 518756 267734
rect 517336 266756 517388 266762
rect 517336 266698 517388 266704
rect 518544 264330 518572 267706
rect 519820 267436 519872 267442
rect 519820 267378 519872 267384
rect 518992 266892 519044 266898
rect 518992 266834 519044 266840
rect 517164 264302 517362 264330
rect 518190 264302 518572 264330
rect 519004 264316 519032 266834
rect 519832 264316 519860 267378
rect 520108 266898 520136 272206
rect 520292 270366 520320 278038
rect 521476 273216 521528 273222
rect 521476 273158 521528 273164
rect 520280 270360 520332 270366
rect 520280 270302 520332 270308
rect 520096 266892 520148 266898
rect 520096 266834 520148 266840
rect 520648 265668 520700 265674
rect 520648 265610 520700 265616
rect 520660 264316 520688 265610
rect 521488 264316 521516 273158
rect 522132 272814 522160 278052
rect 523328 275874 523356 278052
rect 524432 278038 524538 278066
rect 525352 278038 525642 278066
rect 523316 275868 523368 275874
rect 523316 275810 523368 275816
rect 524144 275868 524196 275874
rect 524144 275810 524196 275816
rect 524156 272814 524184 275810
rect 522120 272808 522172 272814
rect 522120 272750 522172 272756
rect 522764 272808 522816 272814
rect 522764 272750 522816 272756
rect 524144 272808 524196 272814
rect 524144 272750 524196 272756
rect 522776 264330 522804 272750
rect 523868 271176 523920 271182
rect 523866 271144 523868 271153
rect 524052 271176 524104 271182
rect 523920 271144 523922 271153
rect 524052 271118 524104 271124
rect 523866 271079 523922 271088
rect 523132 270224 523184 270230
rect 523132 270166 523184 270172
rect 522330 264302 522804 264330
rect 523144 264316 523172 270166
rect 524064 267734 524092 271118
rect 524432 270366 524460 278038
rect 525352 271153 525380 278038
rect 526824 275602 526852 278052
rect 527192 278038 528034 278066
rect 526812 275596 526864 275602
rect 526812 275538 526864 275544
rect 526444 274780 526496 274786
rect 526444 274722 526496 274728
rect 525338 271144 525394 271153
rect 525338 271079 525394 271088
rect 524420 270360 524472 270366
rect 524420 270302 524472 270308
rect 525616 270360 525668 270366
rect 525616 270302 525668 270308
rect 523972 267706 524092 267734
rect 523972 264316 524000 267706
rect 524788 267028 524840 267034
rect 524788 266970 524840 266976
rect 524800 264316 524828 266970
rect 525628 264316 525656 270302
rect 526456 267170 526484 274722
rect 526812 273080 526864 273086
rect 526812 273022 526864 273028
rect 526444 267164 526496 267170
rect 526444 267106 526496 267112
rect 526824 264330 526852 273022
rect 527192 270094 527220 278038
rect 528192 275596 528244 275602
rect 528192 275538 528244 275544
rect 527180 270088 527232 270094
rect 527180 270030 527232 270036
rect 528204 266898 528232 275538
rect 529216 272542 529244 278052
rect 530412 275330 530440 278052
rect 531332 278038 531622 278066
rect 530400 275324 530452 275330
rect 530400 275266 530452 275272
rect 529848 272944 529900 272950
rect 529848 272886 529900 272892
rect 529204 272536 529256 272542
rect 529204 272478 529256 272484
rect 528376 270088 528428 270094
rect 528376 270030 528428 270036
rect 527272 266892 527324 266898
rect 527272 266834 527324 266840
rect 528192 266892 528244 266898
rect 528192 266834 528244 266840
rect 526470 264302 526852 264330
rect 527284 264316 527312 266834
rect 528388 264330 528416 270030
rect 529664 267708 529716 267714
rect 529664 267650 529716 267656
rect 528928 266892 528980 266898
rect 528928 266834 528980 266840
rect 528126 264302 528416 264330
rect 528940 264316 528968 266834
rect 529676 264330 529704 267650
rect 529860 266898 529888 272886
rect 530398 270192 530454 270201
rect 530398 270127 530454 270136
rect 530412 269686 530440 270127
rect 531332 269822 531360 278038
rect 532332 275324 532384 275330
rect 532332 275266 532384 275272
rect 531964 269952 532016 269958
rect 531964 269894 532016 269900
rect 531320 269816 531372 269822
rect 531320 269758 531372 269764
rect 531976 269686 532004 269894
rect 530400 269680 530452 269686
rect 530400 269622 530452 269628
rect 530584 269680 530636 269686
rect 530584 269622 530636 269628
rect 531964 269680 532016 269686
rect 531964 269622 532016 269628
rect 529848 266892 529900 266898
rect 529848 266834 529900 266840
rect 529676 264302 529782 264330
rect 530596 264316 530624 269622
rect 532344 267734 532372 275266
rect 532516 272808 532568 272814
rect 532516 272750 532568 272756
rect 532252 267706 532372 267734
rect 531412 266892 531464 266898
rect 531412 266834 531464 266840
rect 531424 264316 531452 266834
rect 532252 264316 532280 267706
rect 532528 266898 532556 272750
rect 532712 268394 532740 278052
rect 533908 274786 533936 278052
rect 534092 278038 535118 278066
rect 533896 274780 533948 274786
rect 533896 274722 533948 274728
rect 533712 272536 533764 272542
rect 533712 272478 533764 272484
rect 533528 270360 533580 270366
rect 533528 270302 533580 270308
rect 533160 270224 533212 270230
rect 533160 270166 533212 270172
rect 533172 269686 533200 270166
rect 533540 269958 533568 270302
rect 533528 269952 533580 269958
rect 533528 269894 533580 269900
rect 533160 269680 533212 269686
rect 533160 269622 533212 269628
rect 532700 268388 532752 268394
rect 532700 268330 532752 268336
rect 532516 266892 532568 266898
rect 532516 266834 532568 266840
rect 533068 266892 533120 266898
rect 533068 266834 533120 266840
rect 533080 264316 533108 266834
rect 533724 264330 533752 272478
rect 534092 270201 534120 278038
rect 534724 274780 534776 274786
rect 534724 274722 534776 274728
rect 534078 270192 534134 270201
rect 534078 270127 534134 270136
rect 533988 269952 534040 269958
rect 533988 269894 534040 269900
rect 534000 266898 534028 269894
rect 534736 267306 534764 274722
rect 536300 272678 536328 278052
rect 537496 275466 537524 278052
rect 538508 278038 538706 278066
rect 537484 275460 537536 275466
rect 537484 275402 537536 275408
rect 537300 275324 537352 275330
rect 537300 275266 537352 275272
rect 537576 275324 537628 275330
rect 537576 275266 537628 275272
rect 537944 275324 537996 275330
rect 537944 275266 537996 275272
rect 537312 275097 537340 275266
rect 537298 275088 537354 275097
rect 537298 275023 537354 275032
rect 536748 274508 536800 274514
rect 536748 274450 536800 274456
rect 536288 272672 536340 272678
rect 536288 272614 536340 272620
rect 536564 272672 536616 272678
rect 536564 272614 536616 272620
rect 534724 267300 534776 267306
rect 534724 267242 534776 267248
rect 534724 267164 534776 267170
rect 534724 267106 534776 267112
rect 533988 266892 534040 266898
rect 533988 266834 534040 266840
rect 533724 264302 533922 264330
rect 534736 264316 534764 267106
rect 535552 266892 535604 266898
rect 535552 266834 535604 266840
rect 535564 264316 535592 266834
rect 536576 264330 536604 272614
rect 536760 266898 536788 274450
rect 536748 266892 536800 266898
rect 536748 266834 536800 266840
rect 537588 264330 537616 275266
rect 537956 274786 537984 275266
rect 538126 275088 538182 275097
rect 538126 275023 538182 275032
rect 538140 274786 538168 275023
rect 537944 274780 537996 274786
rect 537944 274722 537996 274728
rect 538128 274780 538180 274786
rect 538128 274722 538180 274728
rect 537760 269952 537812 269958
rect 537758 269920 537760 269929
rect 537944 269952 537996 269958
rect 537812 269920 537814 269929
rect 537944 269894 537996 269900
rect 538310 269920 538366 269929
rect 537758 269855 537814 269864
rect 536406 264302 536604 264330
rect 537234 264302 537616 264330
rect 537956 264330 537984 269894
rect 538310 269855 538366 269864
rect 538324 269414 538352 269855
rect 538508 269822 538536 278038
rect 539888 277394 539916 278052
rect 539888 277366 540008 277394
rect 539322 274544 539378 274553
rect 539322 274479 539378 274488
rect 538496 269816 538548 269822
rect 538496 269758 538548 269764
rect 538680 269816 538732 269822
rect 538680 269758 538732 269764
rect 538692 269634 538720 269758
rect 538508 269606 538720 269634
rect 538128 269408 538180 269414
rect 538128 269350 538180 269356
rect 538312 269408 538364 269414
rect 538312 269350 538364 269356
rect 538140 269226 538168 269350
rect 538508 269226 538536 269606
rect 538140 269198 538536 269226
rect 539336 264330 539364 274479
rect 539692 266892 539744 266898
rect 539692 266834 539744 266840
rect 537956 264302 538062 264330
rect 538890 264302 539364 264330
rect 539704 264316 539732 266834
rect 539980 265130 540008 277366
rect 540992 275330 541020 278052
rect 541176 278038 542202 278066
rect 540980 275324 541032 275330
rect 540980 275266 541032 275272
rect 541176 269362 541204 278038
rect 543384 276282 543412 278052
rect 543372 276276 543424 276282
rect 543372 276218 543424 276224
rect 543372 276140 543424 276146
rect 543372 276082 543424 276088
rect 543004 275324 543056 275330
rect 543004 275266 543056 275272
rect 542266 274816 542322 274825
rect 543016 274786 543044 275266
rect 543186 274816 543242 274825
rect 542266 274751 542322 274760
rect 543004 274780 543056 274786
rect 540624 269334 541204 269362
rect 540624 269278 540652 269334
rect 540612 269272 540664 269278
rect 540612 269214 540664 269220
rect 540796 269272 540848 269278
rect 540796 269214 540848 269220
rect 539968 265124 540020 265130
rect 539968 265066 540020 265072
rect 540808 264330 540836 269214
rect 541348 268388 541400 268394
rect 541348 268330 541400 268336
rect 540546 264302 540836 264330
rect 541360 264316 541388 268330
rect 542280 267734 542308 274751
rect 543186 274751 543188 274760
rect 543004 274722 543056 274728
rect 543240 274751 543242 274760
rect 543188 274722 543240 274728
rect 543384 273970 543412 276082
rect 544580 274922 544608 278052
rect 545776 275738 545804 278052
rect 546512 278038 546986 278066
rect 547984 278038 548090 278066
rect 545764 275732 545816 275738
rect 545764 275674 545816 275680
rect 544568 274916 544620 274922
rect 544568 274858 544620 274864
rect 543830 274544 543886 274553
rect 543694 274508 543746 274514
rect 543830 274479 543832 274488
rect 543694 274450 543746 274456
rect 543884 274479 543886 274488
rect 543832 274450 543884 274456
rect 543706 274394 543734 274450
rect 543706 274366 543872 274394
rect 543844 273970 543872 274366
rect 543372 273964 543424 273970
rect 543372 273906 543424 273912
rect 543832 273964 543884 273970
rect 543832 273906 543884 273912
rect 543694 273420 543746 273426
rect 543694 273362 543746 273368
rect 543706 273306 543734 273362
rect 544014 273320 544070 273329
rect 543706 273278 544014 273306
rect 544014 273255 544070 273264
rect 543188 269952 543240 269958
rect 543188 269894 543240 269900
rect 542820 269816 542872 269822
rect 542820 269758 542872 269764
rect 542832 269090 542860 269758
rect 543200 269278 543228 269894
rect 543188 269272 543240 269278
rect 543188 269214 543240 269220
rect 546512 269210 546540 278038
rect 543372 269204 543424 269210
rect 543372 269146 543424 269152
rect 546500 269204 546552 269210
rect 546500 269146 546552 269152
rect 543384 269090 543412 269146
rect 542832 269062 543412 269090
rect 542188 267706 542308 267734
rect 542188 264316 542216 267706
rect 543004 267300 543056 267306
rect 543004 267242 543056 267248
rect 543016 264316 543044 267242
rect 547984 265266 548012 278038
rect 549272 276146 549300 278052
rect 550468 276554 550496 278052
rect 550456 276548 550508 276554
rect 550456 276490 550508 276496
rect 551664 276418 551692 278052
rect 552584 278038 552874 278066
rect 553412 278038 554070 278066
rect 554792 278038 555266 278066
rect 551652 276412 551704 276418
rect 551652 276354 551704 276360
rect 549260 276140 549312 276146
rect 549260 276082 549312 276088
rect 549904 273556 549956 273562
rect 549904 273498 549956 273504
rect 549916 266490 549944 273498
rect 552584 273329 552612 278038
rect 552570 273320 552626 273329
rect 552570 273255 552626 273264
rect 549904 266484 549956 266490
rect 549904 266426 549956 266432
rect 553412 265402 553440 278038
rect 554792 265538 554820 278038
rect 556356 273698 556384 278052
rect 557552 277370 557580 278052
rect 557540 277364 557592 277370
rect 557540 277306 557592 277312
rect 556344 273692 556396 273698
rect 556344 273634 556396 273640
rect 556804 273556 556856 273562
rect 556804 273498 556856 273504
rect 556816 266626 556844 273498
rect 558748 272134 558776 278052
rect 559944 273426 559972 278052
rect 560496 278038 561154 278066
rect 560300 273828 560352 273834
rect 560300 273770 560352 273776
rect 560312 273426 560340 273770
rect 559932 273420 559984 273426
rect 559932 273362 559984 273368
rect 560300 273420 560352 273426
rect 560300 273362 560352 273368
rect 558736 272128 558788 272134
rect 558736 272070 558788 272076
rect 556804 266620 556856 266626
rect 556804 266562 556856 266568
rect 560496 266354 560524 278038
rect 562336 277234 562364 278052
rect 562324 277228 562376 277234
rect 562324 277170 562376 277176
rect 563440 273426 563468 278052
rect 563704 273556 563756 273562
rect 563704 273498 563756 273504
rect 563428 273420 563480 273426
rect 563428 273362 563480 273368
rect 563716 266762 563744 273498
rect 564636 270774 564664 278052
rect 564624 270768 564676 270774
rect 564624 270710 564676 270716
rect 563704 266756 563756 266762
rect 563704 266698 563756 266704
rect 560484 266348 560536 266354
rect 560484 266290 560536 266296
rect 565832 266218 565860 278052
rect 567028 274650 567056 278052
rect 567016 274644 567068 274650
rect 567016 274586 567068 274592
rect 568224 270638 568252 278052
rect 569420 271998 569448 278052
rect 569972 278038 570630 278066
rect 571628 278038 571734 278066
rect 572732 278038 572930 278066
rect 569972 274106 570000 278038
rect 569960 274100 570012 274106
rect 569960 274042 570012 274048
rect 569408 271992 569460 271998
rect 569408 271934 569460 271940
rect 571628 270910 571656 278038
rect 571800 274100 571852 274106
rect 571800 274042 571852 274048
rect 571812 273834 571840 274042
rect 571800 273828 571852 273834
rect 571800 273770 571852 273776
rect 571984 273828 572036 273834
rect 571984 273770 572036 273776
rect 571996 273562 572024 273770
rect 571984 273556 572036 273562
rect 571984 273498 572036 273504
rect 571616 270904 571668 270910
rect 571616 270846 571668 270852
rect 571984 270904 572036 270910
rect 571984 270846 572036 270852
rect 568212 270632 568264 270638
rect 568212 270574 568264 270580
rect 571996 267578 572024 270846
rect 571984 267572 572036 267578
rect 571984 267514 572036 267520
rect 565820 266212 565872 266218
rect 565820 266154 565872 266160
rect 572732 266082 572760 278038
rect 574112 268258 574140 278052
rect 575308 271046 575336 278052
rect 576504 277098 576532 278052
rect 576872 278038 577714 278066
rect 578528 278038 578910 278066
rect 579632 278038 580014 278066
rect 581012 278038 581210 278066
rect 576492 277092 576544 277098
rect 576492 277034 576544 277040
rect 575296 271040 575348 271046
rect 575296 270982 575348 270988
rect 574100 268252 574152 268258
rect 574100 268194 574152 268200
rect 576872 268122 576900 278038
rect 578528 271862 578556 278038
rect 578516 271856 578568 271862
rect 578516 271798 578568 271804
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 576860 268116 576912 268122
rect 576860 268058 576912 268064
rect 578896 267442 578924 271798
rect 579632 270502 579660 278038
rect 579620 270496 579672 270502
rect 579620 270438 579672 270444
rect 581012 269074 581040 278038
rect 582392 271590 582420 278052
rect 583588 274106 583616 278052
rect 583772 278038 584798 278066
rect 583576 274100 583628 274106
rect 583576 274042 583628 274048
rect 582380 271584 582432 271590
rect 582380 271526 582432 271532
rect 581644 270496 581696 270502
rect 581644 270438 581696 270444
rect 581656 269414 581684 270438
rect 581644 269408 581696 269414
rect 581644 269350 581696 269356
rect 581000 269068 581052 269074
rect 581000 269010 581052 269016
rect 583772 268938 583800 278038
rect 585980 271726 586008 278052
rect 587084 275058 587112 278052
rect 587912 278038 588294 278066
rect 587072 275052 587124 275058
rect 587072 274994 587124 275000
rect 585968 271720 586020 271726
rect 585968 271662 586020 271668
rect 585784 271584 585836 271590
rect 585784 271526 585836 271532
rect 583760 268932 583812 268938
rect 583760 268874 583812 268880
rect 585796 267714 585824 271526
rect 587912 268802 587940 278038
rect 589476 271454 589504 278052
rect 590672 273698 590700 278052
rect 590856 278038 591882 278066
rect 590660 273692 590712 273698
rect 590660 273634 590712 273640
rect 589464 271448 589516 271454
rect 589464 271390 589516 271396
rect 587900 268796 587952 268802
rect 587900 268738 587952 268744
rect 590856 268666 590884 278038
rect 593064 271318 593092 278052
rect 594260 275194 594288 278052
rect 595088 278038 595378 278066
rect 596192 278038 596574 278066
rect 594248 275188 594300 275194
rect 594248 275130 594300 275136
rect 595088 274378 595116 278038
rect 595076 274372 595128 274378
rect 595076 274314 595128 274320
rect 595444 274372 595496 274378
rect 595444 274314 595496 274320
rect 593052 271312 593104 271318
rect 593052 271254 593104 271260
rect 590844 268660 590896 268666
rect 590844 268602 590896 268608
rect 585784 267708 585836 267714
rect 585784 267650 585836 267656
rect 578884 267436 578936 267442
rect 578884 267378 578936 267384
rect 595456 266898 595484 274314
rect 596192 269550 596220 278038
rect 597756 273834 597784 278052
rect 598952 274242 598980 278052
rect 600148 276962 600176 278052
rect 600332 278038 601358 278066
rect 601712 278038 602462 278066
rect 600136 276956 600188 276962
rect 600136 276898 600188 276904
rect 598940 274236 598992 274242
rect 598940 274178 598992 274184
rect 597744 273828 597796 273834
rect 597744 273770 597796 273776
rect 596180 269544 596232 269550
rect 596180 269486 596232 269492
rect 595444 266892 595496 266898
rect 595444 266834 595496 266840
rect 572720 266076 572772 266082
rect 572720 266018 572772 266024
rect 600332 265946 600360 278038
rect 601712 268530 601740 278038
rect 603644 276826 603672 278052
rect 603632 276820 603684 276826
rect 603632 276762 603684 276768
rect 604840 270910 604868 278052
rect 605852 278038 606050 278066
rect 604828 270904 604880 270910
rect 604828 270846 604880 270852
rect 601700 268524 601752 268530
rect 601700 268466 601752 268472
rect 600320 265940 600372 265946
rect 600320 265882 600372 265888
rect 605852 265810 605880 278038
rect 607232 272406 607260 278052
rect 608428 276010 608456 278052
rect 609624 276690 609652 278052
rect 609612 276684 609664 276690
rect 609612 276626 609664 276632
rect 608416 276004 608468 276010
rect 608416 275946 608468 275952
rect 607220 272400 607272 272406
rect 607220 272342 607272 272348
rect 610728 272270 610756 278052
rect 610716 272264 610768 272270
rect 610716 272206 610768 272212
rect 611924 271862 611952 278052
rect 612752 278038 613134 278066
rect 611912 271856 611964 271862
rect 611912 271798 611964 271804
rect 612004 271312 612056 271318
rect 612004 271254 612056 271260
rect 612016 267034 612044 271254
rect 612004 267028 612056 267034
rect 612004 266970 612056 266976
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 612752 265674 612780 278038
rect 614316 273222 614344 278052
rect 615512 275874 615540 278052
rect 616156 278038 616722 278066
rect 615500 275868 615552 275874
rect 615500 275810 615552 275816
rect 614304 273216 614356 273222
rect 614304 273158 614356 273164
rect 616156 269686 616184 278038
rect 617812 271182 617840 278052
rect 618640 278038 619022 278066
rect 619652 278038 620218 278066
rect 618640 271318 618668 278038
rect 618628 271312 618680 271318
rect 618628 271254 618680 271260
rect 618904 271312 618956 271318
rect 618904 271254 618956 271260
rect 617800 271176 617852 271182
rect 617800 271118 617852 271124
rect 616144 269680 616196 269686
rect 616144 269622 616196 269628
rect 618916 267170 618944 271254
rect 619652 270230 619680 278038
rect 621400 273086 621428 278052
rect 622596 275602 622624 278052
rect 623806 278038 624004 278066
rect 622584 275596 622636 275602
rect 622584 275538 622636 275544
rect 621388 273080 621440 273086
rect 621388 273022 621440 273028
rect 620284 270496 620336 270502
rect 620284 270438 620336 270444
rect 619640 270224 619692 270230
rect 619640 270166 619692 270172
rect 620296 270094 620324 270438
rect 623976 270230 624004 278038
rect 624988 272950 625016 278052
rect 624976 272944 625028 272950
rect 624976 272886 625028 272892
rect 626092 271590 626120 278052
rect 626552 278038 627302 278066
rect 626080 271584 626132 271590
rect 626080 271526 626132 271532
rect 625804 271176 625856 271182
rect 625804 271118 625856 271124
rect 623964 270224 624016 270230
rect 623964 270166 624016 270172
rect 620284 270088 620336 270094
rect 620284 270030 620336 270036
rect 625816 267306 625844 271118
rect 626552 270366 626580 278038
rect 628484 272814 628512 278052
rect 629680 275330 629708 278052
rect 630692 278038 630890 278066
rect 629668 275324 629720 275330
rect 629668 275266 629720 275272
rect 628472 272808 628524 272814
rect 628472 272750 628524 272756
rect 626540 270360 626592 270366
rect 626540 270302 626592 270308
rect 630692 270094 630720 278038
rect 632072 272542 632100 278052
rect 632060 272536 632112 272542
rect 632060 272478 632112 272484
rect 633268 271318 633296 278052
rect 634372 273970 634400 278052
rect 634360 273964 634412 273970
rect 634360 273906 634412 273912
rect 635568 272678 635596 278052
rect 636764 275466 636792 278052
rect 637592 278038 637974 278066
rect 636752 275460 636804 275466
rect 636752 275402 636804 275408
rect 635556 272672 635608 272678
rect 635556 272614 635608 272620
rect 633256 271312 633308 271318
rect 633256 271254 633308 271260
rect 630680 270088 630732 270094
rect 630680 270030 630732 270036
rect 637592 269822 637620 278038
rect 639156 274514 639184 278052
rect 639144 274508 639196 274514
rect 639144 274450 639196 274456
rect 640352 274378 640380 278052
rect 640536 278038 641470 278066
rect 641732 278038 642666 278066
rect 640340 274372 640392 274378
rect 640340 274314 640392 274320
rect 640536 269958 640564 278038
rect 640524 269952 640576 269958
rect 640524 269894 640576 269900
rect 637580 269816 637632 269822
rect 637580 269758 637632 269764
rect 641732 268394 641760 278038
rect 643848 274786 643876 278052
rect 643836 274780 643888 274786
rect 643836 274722 643888 274728
rect 645044 271182 645072 278052
rect 645872 278038 646254 278066
rect 647252 278038 647450 278066
rect 645032 271176 645084 271182
rect 645032 271118 645084 271124
rect 641720 268388 641772 268394
rect 641720 268330 641772 268336
rect 625804 267300 625856 267306
rect 625804 267242 625856 267248
rect 618904 267164 618956 267170
rect 618904 267106 618956 267112
rect 612740 265668 612792 265674
rect 612740 265610 612792 265616
rect 554780 265532 554832 265538
rect 554780 265474 554832 265480
rect 553400 265396 553452 265402
rect 553400 265338 553452 265344
rect 547972 265260 548024 265266
rect 547972 265202 548024 265208
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 645872 261526 645900 278038
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 560944 259480 560996 259486
rect 560944 259422 560996 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 553490 255640 553546 255649
rect 553490 255575 553492 255584
rect 553544 255575 553546 255584
rect 555424 255604 555476 255610
rect 553492 255546 553544 255552
rect 555424 255546 555476 255552
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 554136 251194 554188 251200
rect 554042 249112 554098 249121
rect 554042 249047 554098 249056
rect 553858 246936 553914 246945
rect 553858 246871 553914 246880
rect 553872 245682 553900 246871
rect 553860 245676 553912 245682
rect 553860 245618 553912 245624
rect 553674 242584 553730 242593
rect 553674 242519 553730 242528
rect 553688 241534 553716 242519
rect 553676 241528 553728 241534
rect 553676 241470 553728 241476
rect 137928 231328 137980 231334
rect 137928 231270 137980 231276
rect 91744 231192 91796 231198
rect 91744 231134 91796 231140
rect 86224 229900 86276 229906
rect 86224 229842 86276 229848
rect 68284 229764 68336 229770
rect 68284 229706 68336 229712
rect 67548 228676 67600 228682
rect 67548 228618 67600 228624
rect 64788 227724 64840 227730
rect 64788 227666 64840 227672
rect 62946 225584 63002 225593
rect 62946 225519 63002 225528
rect 64604 220380 64656 220386
rect 64604 220322 64656 220328
rect 64616 219434 64644 220322
rect 64800 219434 64828 227666
rect 66168 225752 66220 225758
rect 66168 225694 66220 225700
rect 63960 219428 64012 219434
rect 64616 219406 64736 219434
rect 64800 219428 64932 219434
rect 64800 219406 64880 219428
rect 63960 219370 64012 219376
rect 63132 219156 63184 219162
rect 63132 219098 63184 219104
rect 62764 218884 62816 218890
rect 62764 218826 62816 218832
rect 63144 217138 63172 219098
rect 63972 217138 64000 219370
rect 64708 217274 64736 219406
rect 64880 219370 64932 219376
rect 66180 218074 66208 225694
rect 67272 218204 67324 218210
rect 67272 218146 67324 218152
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 66444 218068 66496 218074
rect 66444 218010 66496 218016
rect 64708 217246 64782 217274
rect 61442 217110 61516 217138
rect 62270 217110 62344 217138
rect 63098 217110 63172 217138
rect 63926 217110 64000 217138
rect 61442 216988 61470 217110
rect 62270 216988 62298 217110
rect 63098 216988 63126 217110
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217138 66484 218010
rect 67284 217138 67312 218146
rect 67560 218074 67588 228618
rect 68296 218210 68324 229706
rect 82084 229628 82136 229634
rect 82084 229570 82136 229576
rect 72424 226160 72476 226166
rect 72424 226102 72476 226108
rect 68928 224256 68980 224262
rect 68928 224198 68980 224204
rect 68744 223168 68796 223174
rect 68744 223110 68796 223116
rect 68284 218204 68336 218210
rect 68284 218146 68336 218152
rect 68756 218074 68784 223110
rect 67548 218068 67600 218074
rect 67548 218010 67600 218016
rect 68100 218068 68152 218074
rect 68100 218010 68152 218016
rect 68744 218068 68796 218074
rect 68744 218010 68796 218016
rect 68112 217138 68140 218010
rect 68940 217274 68968 224198
rect 71412 222896 71464 222902
rect 71412 222838 71464 222844
rect 69756 220108 69808 220114
rect 69756 220050 69808 220056
rect 69768 217274 69796 220050
rect 70584 219156 70636 219162
rect 70584 219098 70636 219104
rect 65582 217110 65656 217138
rect 66410 217110 66484 217138
rect 67238 217110 67312 217138
rect 68066 217110 68140 217138
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217110
rect 67238 216988 67266 217110
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 219098
rect 71424 217274 71452 222838
rect 72436 219026 72464 226102
rect 76564 225888 76616 225894
rect 76564 225830 76616 225836
rect 73712 224392 73764 224398
rect 73712 224334 73764 224340
rect 73068 220244 73120 220250
rect 73068 220186 73120 220192
rect 72424 219020 72476 219026
rect 72424 218962 72476 218968
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220186
rect 73724 218074 73752 224334
rect 75828 223032 75880 223038
rect 75828 222974 75880 222980
rect 73896 221604 73948 221610
rect 73896 221546 73948 221552
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221546
rect 75552 218204 75604 218210
rect 75552 218146 75604 218152
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75564 217138 75592 218146
rect 75840 218074 75868 222974
rect 76380 220652 76432 220658
rect 76380 220594 76432 220600
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220594
rect 76576 218210 76604 225830
rect 79968 224664 80020 224670
rect 79968 224606 80020 224612
rect 78588 222624 78640 222630
rect 78588 222566 78640 222572
rect 77208 219020 77260 219026
rect 77208 218962 77260 218968
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218962
rect 78600 218074 78628 222566
rect 79692 220516 79744 220522
rect 79692 220458 79744 220464
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217274 79732 220458
rect 79980 218074 80008 224606
rect 81348 223304 81400 223310
rect 81348 223246 81400 223252
rect 80520 220856 80572 220862
rect 80520 220798 80572 220804
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217274 80560 220798
rect 81360 217274 81388 223246
rect 82096 221610 82124 229570
rect 86236 229094 86264 229842
rect 86144 229066 86264 229094
rect 83464 226024 83516 226030
rect 83464 225966 83516 225972
rect 82084 221604 82136 221610
rect 82084 221546 82136 221552
rect 83004 220992 83056 220998
rect 83004 220934 83056 220940
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217246 79732 217274
rect 80486 217246 80560 217274
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217246
rect 80486 216988 80514 217246
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220934
rect 83476 218074 83504 225966
rect 85488 224528 85540 224534
rect 85488 224470 85540 224476
rect 85304 222760 85356 222766
rect 85304 222702 85356 222708
rect 83832 218884 83884 218890
rect 83832 218826 83884 218832
rect 83464 218068 83516 218074
rect 83464 218010 83516 218016
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218826
rect 85316 218074 85344 222702
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 85304 218068 85356 218074
rect 85304 218010 85356 218016
rect 84672 217138 84700 218010
rect 85500 217274 85528 224470
rect 86144 220862 86172 229066
rect 88248 227860 88300 227866
rect 88248 227802 88300 227808
rect 87972 223576 88024 223582
rect 87972 223518 88024 223524
rect 86316 221604 86368 221610
rect 86316 221546 86368 221552
rect 86132 220856 86184 220862
rect 86132 220798 86184 220804
rect 86328 217274 86356 221546
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87156 217138 87184 218010
rect 87984 217274 88012 223518
rect 88260 218074 88288 227802
rect 89628 227180 89680 227186
rect 89628 227122 89680 227128
rect 89444 224800 89496 224806
rect 89444 224742 89496 224748
rect 88892 223440 88944 223446
rect 88892 223382 88944 223388
rect 88904 222630 88932 223382
rect 88892 222624 88944 222630
rect 88892 222566 88944 222572
rect 89456 218074 89484 224742
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227122
rect 91284 222012 91336 222018
rect 91284 221954 91336 221960
rect 90456 218068 90508 218074
rect 90456 218010 90508 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90468 217138 90496 218010
rect 91296 217274 91324 221954
rect 91756 218074 91784 231134
rect 128268 231056 128320 231062
rect 128268 230998 128320 231004
rect 118608 230920 118660 230926
rect 118608 230862 118660 230868
rect 110328 230784 110380 230790
rect 110328 230726 110380 230732
rect 97908 230648 97960 230654
rect 97908 230590 97960 230596
rect 95240 230172 95292 230178
rect 95240 230114 95292 230120
rect 93768 228812 93820 228818
rect 93768 228754 93820 228760
rect 93780 218074 93808 228754
rect 95252 227866 95280 230114
rect 95240 227860 95292 227866
rect 95240 227802 95292 227808
rect 96436 227316 96488 227322
rect 96436 227258 96488 227264
rect 96252 224936 96304 224942
rect 96252 224878 96304 224884
rect 94596 221876 94648 221882
rect 94596 221818 94648 221824
rect 91744 218068 91796 218074
rect 91744 218010 91796 218016
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 93768 218068 93820 218074
rect 93768 218010 93820 218016
rect 90422 217110 90496 217138
rect 91250 217246 91324 217274
rect 92066 217252 92118 217258
rect 90422 216988 90450 217110
rect 91250 216988 91278 217246
rect 92066 217194 92118 217200
rect 92078 216988 92106 217194
rect 92952 217138 92980 218010
rect 93768 217456 93820 217462
rect 93768 217398 93820 217404
rect 93780 217138 93808 217398
rect 94608 217274 94636 221818
rect 96264 218074 96292 224878
rect 95424 218068 95476 218074
rect 95424 218010 95476 218016
rect 96252 218068 96304 218074
rect 96252 218010 96304 218016
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 94562 217246 94636 217274
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217246
rect 95436 217138 95464 218010
rect 96448 217274 96476 227258
rect 97724 221740 97776 221746
rect 97724 221682 97776 221688
rect 97736 219434 97764 221682
rect 97736 219406 97856 219434
rect 97080 218068 97132 218074
rect 97080 218010 97132 218016
rect 95390 217110 95464 217138
rect 96218 217246 96476 217274
rect 95390 216988 95418 217110
rect 96218 216988 96246 217246
rect 97092 217138 97120 218010
rect 97828 217274 97856 219406
rect 97920 218090 97948 230590
rect 102140 229492 102192 229498
rect 102140 229434 102192 229440
rect 100668 229084 100720 229090
rect 100668 229026 100720 229032
rect 99288 222624 99340 222630
rect 99288 222566 99340 222572
rect 97920 218074 98040 218090
rect 99300 218074 99328 222566
rect 100392 218612 100444 218618
rect 100392 218554 100444 218560
rect 97920 218068 98052 218074
rect 97920 218062 98000 218068
rect 98000 218010 98052 218016
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97828 217246 97902 217274
rect 97046 217110 97120 217138
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218554
rect 100680 218074 100708 229026
rect 102152 227458 102180 229434
rect 106188 229084 106240 229090
rect 106188 229026 106240 229032
rect 102140 227452 102192 227458
rect 102140 227394 102192 227400
rect 103428 227452 103480 227458
rect 103428 227394 103480 227400
rect 102048 224120 102100 224126
rect 102048 224062 102100 224068
rect 101220 220788 101272 220794
rect 101220 220730 101272 220736
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101232 217274 101260 220730
rect 102060 217274 102088 224062
rect 103440 218074 103468 227394
rect 106004 223984 106056 223990
rect 106004 223926 106056 223932
rect 104532 221332 104584 221338
rect 104532 221274 104584 221280
rect 102876 218068 102928 218074
rect 102876 218010 102928 218016
rect 103428 218068 103480 218074
rect 103428 218010 103480 218016
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217246 101260 217274
rect 102014 217246 102088 217274
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217246
rect 102014 216988 102042 217246
rect 102888 217138 102916 218010
rect 103704 217592 103756 217598
rect 103704 217534 103756 217540
rect 103716 217138 103744 217534
rect 104544 217274 104572 221274
rect 105820 219496 105872 219502
rect 105820 219438 105872 219444
rect 105832 218618 105860 219438
rect 105820 218612 105872 218618
rect 105820 218554 105872 218560
rect 106016 218074 106044 223926
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106004 218068 106056 218074
rect 106004 218010 106056 218016
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106200 217274 106228 229026
rect 110144 227588 110196 227594
rect 110144 227530 110196 227536
rect 106924 226500 106976 226506
rect 106924 226442 106976 226448
rect 106936 219298 106964 226442
rect 108672 223848 108724 223854
rect 108672 223790 108724 223796
rect 107660 223440 107712 223446
rect 107660 223382 107712 223388
rect 108304 223440 108356 223446
rect 108304 223382 108356 223388
rect 107672 222630 107700 223382
rect 107660 222624 107712 222630
rect 107660 222566 107712 222572
rect 108316 222494 108344 223382
rect 108304 222488 108356 222494
rect 108304 222430 108356 222436
rect 107844 219972 107896 219978
rect 107844 219914 107896 219920
rect 106924 219292 106976 219298
rect 106924 219234 106976 219240
rect 107016 218476 107068 218482
rect 107016 218418 107068 218424
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218418
rect 107856 217274 107884 219914
rect 108684 217274 108712 223790
rect 110156 218074 110184 227530
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 110144 218068 110196 218074
rect 110144 218010 110196 218016
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110340 217274 110368 230726
rect 111064 229356 111116 229362
rect 111064 229298 111116 229304
rect 111076 227730 111104 229298
rect 112812 228268 112864 228274
rect 112812 228210 112864 228216
rect 111064 227724 111116 227730
rect 111064 227666 111116 227672
rect 111984 222148 112036 222154
rect 111984 222090 112036 222096
rect 111156 221196 111208 221202
rect 111156 221138 111208 221144
rect 111168 217274 111196 221138
rect 111996 217274 112024 222090
rect 112824 217274 112852 228210
rect 117228 227724 117280 227730
rect 117228 227666 117280 227672
rect 115296 223712 115348 223718
rect 115296 223654 115348 223660
rect 114468 219836 114520 219842
rect 114468 219778 114520 219784
rect 113640 219292 113692 219298
rect 113640 219234 113692 219240
rect 109466 217110 109540 217138
rect 110294 217246 110368 217274
rect 111122 217246 111196 217274
rect 111950 217246 112024 217274
rect 112778 217246 112852 217274
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111122 216988 111150 217246
rect 111950 216988 111978 217246
rect 112778 216988 112806 217246
rect 113652 217138 113680 219234
rect 114480 217274 114508 219778
rect 115308 217274 115336 223654
rect 117240 218074 117268 227666
rect 118424 222488 118476 222494
rect 118424 222430 118476 222436
rect 118436 219434 118464 222430
rect 118436 219406 118556 219434
rect 117964 219156 118016 219162
rect 117964 219098 118016 219104
rect 117976 218346 118004 219098
rect 117964 218340 118016 218346
rect 117964 218282 118016 218288
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 117780 218068 117832 218074
rect 117780 218010 117832 218016
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 115262 217246 115336 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115262 216988 115290 217246
rect 116136 217138 116164 218010
rect 116952 217728 117004 217734
rect 116952 217670 117004 217676
rect 116964 217138 116992 217670
rect 117792 217138 117820 218010
rect 118528 217274 118556 219406
rect 118620 218090 118648 230862
rect 126888 230036 126940 230042
rect 126888 229978 126940 229984
rect 123484 229220 123536 229226
rect 123484 229162 123536 229168
rect 119988 228132 120040 228138
rect 119988 228074 120040 228080
rect 118620 218074 118740 218090
rect 120000 218074 120028 228074
rect 122748 226908 122800 226914
rect 122748 226850 122800 226856
rect 122564 226296 122616 226302
rect 122564 226238 122616 226244
rect 121092 219700 121144 219706
rect 121092 219642 121144 219648
rect 120264 218612 120316 218618
rect 120264 218554 120316 218560
rect 118620 218068 118752 218074
rect 118620 218062 118700 218068
rect 118700 218010 118752 218016
rect 119436 218068 119488 218074
rect 119436 218010 119488 218016
rect 119988 218068 120040 218074
rect 119988 218010 120040 218016
rect 118528 217246 118602 217274
rect 116090 217110 116164 217138
rect 116918 217110 116992 217138
rect 117746 217110 117820 217138
rect 116090 216988 116118 217110
rect 116918 216988 116946 217110
rect 117746 216988 117774 217110
rect 118574 216988 118602 217246
rect 119448 217138 119476 218010
rect 120276 217138 120304 218554
rect 121104 217274 121132 219642
rect 122576 218074 122604 226238
rect 121920 218068 121972 218074
rect 121920 218010 121972 218016
rect 122564 218068 122616 218074
rect 122564 218010 122616 218016
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 218010
rect 122760 217274 122788 226850
rect 123496 218346 123524 229162
rect 126704 227996 126756 228002
rect 126704 227938 126756 227944
rect 125232 225480 125284 225486
rect 125232 225422 125284 225428
rect 124404 221060 124456 221066
rect 124404 221002 124456 221008
rect 123484 218340 123536 218346
rect 123484 218282 123536 218288
rect 123576 218204 123628 218210
rect 123576 218146 123628 218152
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 218146
rect 124416 217274 124444 221002
rect 125244 217274 125272 225422
rect 126520 222624 126572 222630
rect 126520 222566 126572 222572
rect 126532 222358 126560 222566
rect 126520 222352 126572 222358
rect 126520 222294 126572 222300
rect 126716 218074 126744 227938
rect 126060 218068 126112 218074
rect 126060 218010 126112 218016
rect 126704 218068 126756 218074
rect 126704 218010 126756 218016
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 218010
rect 126900 217274 126928 229978
rect 127624 219972 127676 219978
rect 127624 219914 127676 219920
rect 127808 219972 127860 219978
rect 127808 219914 127860 219920
rect 127636 219706 127664 219914
rect 127624 219700 127676 219706
rect 127624 219642 127676 219648
rect 127820 219570 127848 219914
rect 127808 219564 127860 219570
rect 127808 219506 127860 219512
rect 128280 218074 128308 230998
rect 130384 230444 130436 230450
rect 130384 230386 130436 230392
rect 129556 226772 129608 226778
rect 129556 226714 129608 226720
rect 129372 225344 129424 225350
rect 129372 225286 129424 225292
rect 129384 218074 129412 225286
rect 127716 218068 127768 218074
rect 127716 218010 127768 218016
rect 128268 218068 128320 218074
rect 128268 218010 128320 218016
rect 128544 218068 128596 218074
rect 128544 218010 128596 218016
rect 129372 218068 129424 218074
rect 129372 218010 129424 218016
rect 126026 217110 126100 217138
rect 126854 217246 126928 217274
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 218010
rect 128556 217138 128584 218010
rect 129568 217274 129596 226714
rect 130396 225214 130424 230386
rect 133788 230308 133840 230314
rect 133788 230250 133840 230256
rect 133512 227860 133564 227866
rect 133512 227802 133564 227808
rect 130384 225208 130436 225214
rect 130384 225150 130436 225156
rect 132408 225072 132460 225078
rect 132408 225014 132460 225020
rect 132420 218346 132448 225014
rect 132592 219156 132644 219162
rect 132592 219098 132644 219104
rect 131856 218340 131908 218346
rect 131856 218282 131908 218288
rect 132408 218340 132460 218346
rect 132408 218282 132460 218288
rect 130200 218068 130252 218074
rect 130200 218010 130252 218016
rect 127682 217110 127756 217138
rect 128510 217110 128584 217138
rect 129338 217246 129596 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 218010
rect 131028 217864 131080 217870
rect 131028 217806 131080 217812
rect 131040 217138 131068 217806
rect 131868 217138 131896 218282
rect 132604 218226 132632 219098
rect 132512 218198 132632 218226
rect 132512 218074 132540 218198
rect 133524 218074 133552 227802
rect 133800 219434 133828 230250
rect 136548 226636 136600 226642
rect 136548 226578 136600 226584
rect 135076 225208 135128 225214
rect 135076 225150 135128 225156
rect 134340 219564 134392 219570
rect 134340 219506 134392 219512
rect 133708 219406 133828 219434
rect 132500 218068 132552 218074
rect 132500 218010 132552 218016
rect 132684 218068 132736 218074
rect 132684 218010 132736 218016
rect 133512 218068 133564 218074
rect 133512 218010 133564 218016
rect 132696 217138 132724 218010
rect 133708 217274 133736 219406
rect 134352 217274 134380 219506
rect 130166 217110 130240 217138
rect 130994 217110 131068 217138
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133736 217274
rect 134306 217246 134380 217274
rect 135088 217274 135116 225150
rect 136560 218074 136588 226578
rect 137940 219434 137968 231270
rect 140042 229120 140098 229129
rect 140042 229055 140098 229064
rect 139306 228304 139362 228313
rect 139306 228239 139362 228248
rect 139124 222352 139176 222358
rect 139124 222294 139176 222300
rect 137664 219406 137968 219434
rect 136824 218340 136876 218346
rect 136824 218282 136876 218288
rect 135996 218068 136048 218074
rect 135996 218010 136048 218016
rect 136548 218068 136600 218074
rect 136548 218010 136600 218016
rect 135088 217246 135162 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217110
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135134 216988 135162 217246
rect 136008 217138 136036 218010
rect 136836 217138 136864 218282
rect 137664 217274 137692 219406
rect 139136 218074 139164 222294
rect 138480 218068 138532 218074
rect 138480 218010 138532 218016
rect 139124 218068 139176 218074
rect 139124 218010 139176 218016
rect 135962 217110 136036 217138
rect 136790 217110 136864 217138
rect 137618 217246 137692 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217110
rect 137618 216988 137646 217246
rect 138492 217138 138520 218010
rect 139320 217274 139348 228239
rect 140056 219026 140084 229055
rect 141160 228410 141188 231676
rect 141344 231662 141818 231690
rect 142172 231662 142462 231690
rect 142816 231662 143106 231690
rect 141148 228404 141200 228410
rect 141148 228346 141200 228352
rect 141148 226160 141200 226166
rect 141146 226128 141148 226137
rect 141200 226128 141202 226137
rect 141146 226063 141202 226072
rect 141344 221474 141372 231662
rect 142172 227050 142200 231662
rect 142434 230480 142490 230489
rect 142434 230415 142436 230424
rect 142488 230415 142490 230424
rect 142620 230444 142672 230450
rect 142436 230386 142488 230392
rect 142620 230386 142672 230392
rect 142632 229770 142660 230386
rect 142620 229764 142672 229770
rect 142620 229706 142672 229712
rect 142816 228698 142844 231662
rect 142988 229084 143040 229090
rect 142988 229026 143040 229032
rect 143448 229084 143500 229090
rect 143448 229026 143500 229032
rect 142632 228670 142844 228698
rect 143000 228682 143028 229026
rect 142988 228676 143040 228682
rect 142632 228546 142660 228670
rect 142988 228618 143040 228624
rect 142620 228540 142672 228546
rect 142620 228482 142672 228488
rect 142988 228540 143040 228546
rect 142988 228482 143040 228488
rect 143000 228313 143028 228482
rect 142986 228304 143042 228313
rect 142986 228239 143042 228248
rect 142160 227044 142212 227050
rect 142160 226986 142212 226992
rect 143264 227044 143316 227050
rect 143264 226986 143316 226992
rect 141516 226160 141568 226166
rect 141516 226102 141568 226108
rect 141528 225622 141556 226102
rect 141516 225616 141568 225622
rect 141516 225558 141568 225564
rect 141792 225616 141844 225622
rect 141792 225558 141844 225564
rect 141332 221468 141384 221474
rect 141332 221410 141384 221416
rect 140778 220416 140834 220425
rect 140778 220351 140834 220360
rect 140792 219706 140820 220351
rect 140780 219700 140832 219706
rect 140780 219642 140832 219648
rect 140964 219700 141016 219706
rect 140964 219642 141016 219648
rect 140044 219020 140096 219026
rect 140044 218962 140096 218968
rect 139492 218340 139544 218346
rect 139492 218282 139544 218288
rect 140136 218340 140188 218346
rect 140136 218282 140188 218288
rect 139504 218074 139532 218282
rect 139492 218068 139544 218074
rect 139492 218010 139544 218016
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218282
rect 140976 217274 141004 219642
rect 141804 217274 141832 225558
rect 142342 220416 142398 220425
rect 141976 220380 142028 220386
rect 142342 220351 142398 220360
rect 141976 220322 142028 220328
rect 141988 219745 142016 220322
rect 142356 220182 142384 220351
rect 142344 220176 142396 220182
rect 142158 220144 142214 220153
rect 142344 220118 142396 220124
rect 142158 220079 142160 220088
rect 142212 220079 142214 220088
rect 142160 220050 142212 220056
rect 141974 219736 142030 219745
rect 141974 219671 142030 219680
rect 143276 218754 143304 226986
rect 142620 218748 142672 218754
rect 142620 218690 142672 218696
rect 143264 218748 143316 218754
rect 143264 218690 143316 218696
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218690
rect 143460 217274 143488 229026
rect 143736 218890 143764 231676
rect 144104 231662 144394 231690
rect 144104 230489 144132 231662
rect 144090 230480 144146 230489
rect 144090 230415 144146 230424
rect 143998 229528 144054 229537
rect 143998 229463 144000 229472
rect 144052 229463 144054 229472
rect 144184 229492 144236 229498
rect 144000 229434 144052 229440
rect 144184 229434 144236 229440
rect 144196 219745 144224 229434
rect 145024 226166 145052 231676
rect 145392 231662 145682 231690
rect 146326 231662 146616 231690
rect 145392 229537 145420 231662
rect 146208 231600 146260 231606
rect 146208 231542 146260 231548
rect 146220 230450 146248 231542
rect 146208 230444 146260 230450
rect 146208 230386 146260 230392
rect 145378 229528 145434 229537
rect 145378 229463 145434 229472
rect 146206 229392 146262 229401
rect 146206 229327 146262 229336
rect 146220 229090 146248 229327
rect 146208 229084 146260 229090
rect 146208 229026 146260 229032
rect 146392 229084 146444 229090
rect 146392 229026 146444 229032
rect 146404 228970 146432 229026
rect 145944 228942 146432 228970
rect 145944 228546 145972 228942
rect 145932 228540 145984 228546
rect 145932 228482 145984 228488
rect 146116 228540 146168 228546
rect 146116 228482 146168 228488
rect 145012 226160 145064 226166
rect 145196 226160 145248 226166
rect 145012 226102 145064 226108
rect 145194 226128 145196 226137
rect 145248 226128 145250 226137
rect 145194 226063 145250 226072
rect 145930 222320 145986 222329
rect 145930 222255 145986 222264
rect 144826 220416 144882 220425
rect 144826 220351 144882 220360
rect 144182 219736 144238 219745
rect 144182 219671 144238 219680
rect 143724 218884 143776 218890
rect 143724 218826 143776 218832
rect 144840 218754 144868 220351
rect 145944 218754 145972 222255
rect 144276 218748 144328 218754
rect 144276 218690 144328 218696
rect 144828 218748 144880 218754
rect 144828 218690 144880 218696
rect 145104 218748 145156 218754
rect 145104 218690 145156 218696
rect 145932 218748 145984 218754
rect 145932 218690 145984 218696
rect 142586 217110 142660 217138
rect 143414 217246 143488 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144288 217138 144316 218690
rect 145116 217138 145144 218690
rect 146128 217274 146156 228482
rect 146588 226506 146616 231662
rect 146760 231464 146812 231470
rect 146760 231406 146812 231412
rect 146576 226500 146628 226506
rect 146576 226442 146628 226448
rect 146772 226166 146800 231406
rect 146956 229498 146984 231676
rect 147232 231662 147614 231690
rect 147968 231662 148258 231690
rect 147232 231470 147260 231662
rect 147220 231464 147272 231470
rect 147220 231406 147272 231412
rect 147634 230444 147686 230450
rect 147634 230386 147686 230392
rect 147646 230194 147674 230386
rect 147324 230166 147674 230194
rect 147128 229560 147180 229566
rect 147128 229502 147180 229508
rect 146944 229492 146996 229498
rect 146944 229434 146996 229440
rect 147140 229129 147168 229502
rect 147126 229120 147182 229129
rect 147126 229055 147182 229064
rect 146760 226160 146812 226166
rect 146760 226102 146812 226108
rect 147324 224954 147352 230166
rect 147968 229809 147996 231662
rect 147586 229800 147642 229809
rect 147954 229800 148010 229809
rect 147586 229735 147642 229744
rect 147772 229764 147824 229770
rect 147600 229362 147628 229735
rect 147954 229735 148010 229744
rect 147772 229706 147824 229712
rect 147784 229650 147812 229706
rect 147784 229634 148180 229650
rect 147784 229628 148192 229634
rect 147784 229622 148140 229628
rect 148140 229570 148192 229576
rect 147770 229392 147826 229401
rect 147588 229356 147640 229362
rect 147770 229327 147772 229336
rect 147588 229298 147640 229304
rect 147824 229327 147826 229336
rect 147772 229298 147824 229304
rect 148888 228410 148916 231676
rect 149532 230450 149560 231676
rect 149808 231662 150190 231690
rect 150544 231662 150834 231690
rect 151004 231662 151478 231690
rect 149520 230444 149572 230450
rect 149520 230386 149572 230392
rect 148876 228404 148928 228410
rect 148876 228346 148928 228352
rect 148968 226160 149020 226166
rect 148968 226102 149020 226108
rect 146588 224926 147352 224954
rect 146588 223258 146616 224926
rect 146496 223230 146616 223258
rect 146496 223174 146524 223230
rect 146484 223168 146536 223174
rect 146484 223110 146536 223116
rect 146668 223168 146720 223174
rect 146668 223110 146720 223116
rect 146680 222494 146708 223110
rect 147310 223000 147366 223009
rect 147310 222935 147366 222944
rect 146668 222488 146720 222494
rect 146668 222430 146720 222436
rect 147128 222352 147180 222358
rect 147126 222320 147128 222329
rect 147180 222320 147182 222329
rect 147126 222255 147182 222264
rect 147324 219434 147352 222935
rect 147588 221468 147640 221474
rect 147588 221410 147640 221416
rect 147128 219428 147352 219434
rect 147180 219406 147352 219428
rect 147128 219370 147180 219376
rect 146760 218884 146812 218890
rect 146760 218826 146812 218832
rect 144242 217110 144316 217138
rect 145070 217110 145144 217138
rect 145898 217246 146156 217274
rect 144242 216988 144270 217110
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218826
rect 147600 217274 147628 221410
rect 148980 218754 149008 226102
rect 149808 225758 149836 231662
rect 150544 231606 150572 231662
rect 150532 231600 150584 231606
rect 150532 231542 150584 231548
rect 150346 229392 150402 229401
rect 150346 229327 150402 229336
rect 150072 226500 150124 226506
rect 150072 226442 150124 226448
rect 149796 225752 149848 225758
rect 149796 225694 149848 225700
rect 150084 218754 150112 226442
rect 150360 219434 150388 229327
rect 151004 224954 151032 231662
rect 151176 229356 151228 229362
rect 151176 229298 151228 229304
rect 151188 225842 151216 229298
rect 150912 224926 151032 224954
rect 151096 225814 151216 225842
rect 150912 220153 150940 224926
rect 151096 220930 151124 225814
rect 151268 225752 151320 225758
rect 151268 225694 151320 225700
rect 151084 220924 151136 220930
rect 151084 220866 151136 220872
rect 151084 220312 151136 220318
rect 151084 220254 151136 220260
rect 151280 220266 151308 225694
rect 151912 223304 151964 223310
rect 151912 223246 151964 223252
rect 151924 223145 151952 223246
rect 151910 223136 151966 223145
rect 151910 223071 151966 223080
rect 151450 223000 151506 223009
rect 151506 222958 151814 222986
rect 151450 222935 151506 222944
rect 151786 222902 151814 222958
rect 151636 222896 151688 222902
rect 151636 222838 151688 222844
rect 151774 222896 151826 222902
rect 151774 222838 151826 222844
rect 151648 222737 151676 222838
rect 152108 222737 152136 231676
rect 152464 231328 152516 231334
rect 152464 231270 152516 231276
rect 152476 230518 152504 231270
rect 152464 230512 152516 230518
rect 152464 230454 152516 230460
rect 152464 228676 152516 228682
rect 152464 228618 152516 228624
rect 152476 228410 152504 228618
rect 152464 228404 152516 228410
rect 152464 228346 152516 228352
rect 152752 224262 152780 231676
rect 153396 229226 153424 231676
rect 153580 231662 154054 231690
rect 154698 231662 154988 231690
rect 153384 229220 153436 229226
rect 153384 229162 153436 229168
rect 153108 228676 153160 228682
rect 153108 228618 153160 228624
rect 152740 224256 152792 224262
rect 152740 224198 152792 224204
rect 152372 223032 152424 223038
rect 152372 222974 152424 222980
rect 151634 222728 151690 222737
rect 151634 222663 151690 222672
rect 152094 222728 152150 222737
rect 152094 222663 152150 222672
rect 151726 220552 151782 220561
rect 151726 220487 151728 220496
rect 151780 220487 151782 220496
rect 151912 220516 151964 220522
rect 151728 220458 151780 220464
rect 151912 220458 151964 220464
rect 151450 220416 151506 220425
rect 151506 220386 151814 220402
rect 151506 220380 151826 220386
rect 151506 220374 151774 220380
rect 151450 220351 151506 220360
rect 151774 220322 151826 220328
rect 151096 220153 151124 220254
rect 151280 220238 151676 220266
rect 150898 220144 150954 220153
rect 150898 220079 150954 220088
rect 151082 220144 151138 220153
rect 151082 220079 151138 220088
rect 151452 220108 151504 220114
rect 151452 220050 151504 220056
rect 151464 219434 151492 220050
rect 150268 219406 150388 219434
rect 150912 219406 151492 219434
rect 148416 218748 148468 218754
rect 148416 218690 148468 218696
rect 148968 218748 149020 218754
rect 148968 218690 149020 218696
rect 149244 218748 149296 218754
rect 149244 218690 149296 218696
rect 150072 218748 150124 218754
rect 150072 218690 150124 218696
rect 146726 217110 146800 217138
rect 147554 217246 147628 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217246
rect 148428 217138 148456 218690
rect 149256 217138 149284 218690
rect 150268 217274 150296 219406
rect 150912 217274 150940 219406
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150296 217274
rect 150866 217246 150940 217274
rect 151648 217274 151676 220238
rect 151924 220153 151952 220458
rect 151910 220144 151966 220153
rect 151910 220079 151966 220088
rect 152384 218482 152412 222974
rect 153120 218482 153148 228618
rect 153580 220522 153608 231662
rect 153844 229356 153896 229362
rect 153844 229298 153896 229304
rect 153568 220516 153620 220522
rect 153568 220458 153620 220464
rect 153856 219026 153884 229298
rect 154960 223174 154988 231662
rect 155328 224398 155356 231676
rect 155972 229634 156000 231676
rect 156156 231662 156630 231690
rect 156892 231662 157274 231690
rect 157918 231662 158300 231690
rect 155960 229628 156012 229634
rect 155960 229570 156012 229576
rect 155316 224392 155368 224398
rect 155316 224334 155368 224340
rect 155868 224392 155920 224398
rect 155868 224334 155920 224340
rect 154948 223168 155000 223174
rect 154948 223110 155000 223116
rect 155040 220924 155092 220930
rect 155040 220866 155092 220872
rect 154212 220516 154264 220522
rect 154212 220458 154264 220464
rect 153844 219020 153896 219026
rect 153844 218962 153896 218968
rect 153384 218884 153436 218890
rect 153384 218826 153436 218832
rect 152372 218476 152424 218482
rect 152372 218418 152424 218424
rect 152556 218476 152608 218482
rect 152556 218418 152608 218424
rect 153108 218476 153160 218482
rect 153108 218418 153160 218424
rect 151648 217246 151722 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150866 216988 150894 217246
rect 151694 216988 151722 217246
rect 152568 217138 152596 218418
rect 153396 217138 153424 218826
rect 154224 217274 154252 220458
rect 155052 217274 155080 220866
rect 155880 217274 155908 224334
rect 156156 220658 156184 231662
rect 156512 231328 156564 231334
rect 156512 231270 156564 231276
rect 156524 229362 156552 231270
rect 156694 229936 156750 229945
rect 156694 229871 156696 229880
rect 156748 229871 156750 229880
rect 156696 229842 156748 229848
rect 156512 229356 156564 229362
rect 156512 229298 156564 229304
rect 156694 227488 156750 227497
rect 156694 227423 156750 227432
rect 156708 227186 156736 227423
rect 156696 227180 156748 227186
rect 156696 227122 156748 227128
rect 156892 224954 156920 231662
rect 157294 230172 157346 230178
rect 157294 230114 157346 230120
rect 157432 230172 157484 230178
rect 157432 230114 157484 230120
rect 157306 229770 157334 230114
rect 157444 229945 157472 230114
rect 157430 229936 157486 229945
rect 157430 229871 157486 229880
rect 157294 229764 157346 229770
rect 157294 229706 157346 229712
rect 157340 229628 157392 229634
rect 157340 229570 157392 229576
rect 157062 229392 157118 229401
rect 157062 229327 157064 229336
rect 157116 229327 157118 229336
rect 157064 229298 157116 229304
rect 156432 224926 156920 224954
rect 156432 223310 156460 224926
rect 156420 223304 156472 223310
rect 156420 223246 156472 223252
rect 156604 223304 156656 223310
rect 156604 223246 156656 223252
rect 156420 223168 156472 223174
rect 156420 223110 156472 223116
rect 156432 222902 156460 223110
rect 156420 222896 156472 222902
rect 156420 222838 156472 222844
rect 156616 222766 156644 223246
rect 156786 223136 156842 223145
rect 156786 223071 156842 223080
rect 156800 222766 156828 223071
rect 156604 222760 156656 222766
rect 156604 222702 156656 222708
rect 156788 222760 156840 222766
rect 156788 222702 156840 222708
rect 157352 222194 157380 229570
rect 158272 225894 158300 231662
rect 158548 229906 158576 231676
rect 158916 231662 159206 231690
rect 158536 229900 158588 229906
rect 158536 229842 158588 229848
rect 158260 225888 158312 225894
rect 158260 225830 158312 225836
rect 157524 223032 157576 223038
rect 157524 222974 157576 222980
rect 157260 222166 157380 222194
rect 156144 220652 156196 220658
rect 156144 220594 156196 220600
rect 156604 220652 156656 220658
rect 156604 220594 156656 220600
rect 156616 220250 156644 220594
rect 156970 220552 157026 220561
rect 156788 220516 156840 220522
rect 156970 220487 156972 220496
rect 156788 220458 156840 220464
rect 157024 220487 157026 220496
rect 156972 220458 157024 220464
rect 156800 220250 156828 220458
rect 156604 220244 156656 220250
rect 156604 220186 156656 220192
rect 156788 220244 156840 220250
rect 156788 220186 156840 220192
rect 156328 219292 156380 219298
rect 156328 219234 156380 219240
rect 156340 218890 156368 219234
rect 156328 218884 156380 218890
rect 156328 218826 156380 218832
rect 157260 218482 157288 222166
rect 156696 218476 156748 218482
rect 156696 218418 156748 218424
rect 157248 218476 157300 218482
rect 157248 218418 157300 218424
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217246 154252 217274
rect 155006 217246 155080 217274
rect 155834 217246 155908 217274
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217246
rect 155006 216988 155034 217246
rect 155834 216988 155862 217246
rect 156708 217138 156736 218418
rect 157536 217138 157564 222974
rect 158350 220960 158406 220969
rect 158350 220895 158406 220904
rect 158364 217138 158392 220895
rect 158916 220522 158944 231662
rect 159640 227180 159692 227186
rect 159640 227122 159692 227128
rect 159652 224398 159680 227122
rect 159640 224392 159692 224398
rect 159640 224334 159692 224340
rect 159836 222766 159864 231676
rect 160006 228168 160062 228177
rect 160006 228103 160062 228112
rect 159824 222760 159876 222766
rect 159824 222702 159876 222708
rect 158904 220516 158956 220522
rect 158904 220458 158956 220464
rect 160020 219434 160048 228103
rect 160480 224670 160508 231676
rect 161124 230178 161152 231676
rect 161112 230172 161164 230178
rect 161112 230114 161164 230120
rect 161768 229226 161796 231676
rect 161952 231662 162426 231690
rect 161756 229220 161808 229226
rect 161756 229162 161808 229168
rect 160468 224664 160520 224670
rect 160468 224606 160520 224612
rect 161664 224392 161716 224398
rect 161664 224334 161716 224340
rect 160836 220516 160888 220522
rect 160836 220458 160888 220464
rect 159180 219428 159232 219434
rect 159180 219370 159232 219376
rect 160008 219428 160060 219434
rect 160008 219370 160060 219376
rect 159192 217138 159220 219370
rect 160008 219292 160060 219298
rect 160008 219234 160060 219240
rect 160020 217138 160048 219234
rect 160848 217138 160876 220458
rect 161676 217138 161704 224334
rect 161952 223310 161980 231662
rect 163056 226030 163084 231676
rect 163700 231334 163728 231676
rect 163688 231328 163740 231334
rect 163688 231270 163740 231276
rect 163964 229900 164016 229906
rect 163964 229842 164016 229848
rect 163044 226024 163096 226030
rect 163044 225966 163096 225972
rect 161940 223304 161992 223310
rect 161940 223246 161992 223252
rect 162308 223304 162360 223310
rect 162308 223246 162360 223252
rect 161938 221640 161994 221649
rect 161938 221575 161940 221584
rect 161992 221575 161994 221584
rect 162124 221604 162176 221610
rect 161940 221546 161992 221552
rect 162124 221546 162176 221552
rect 162136 220930 162164 221546
rect 162124 220924 162176 220930
rect 162124 220866 162176 220872
rect 162320 218890 162348 223246
rect 163780 220924 163832 220930
rect 163780 220866 163832 220872
rect 163792 220522 163820 220866
rect 163780 220516 163832 220522
rect 163780 220458 163832 220464
rect 163976 219434 164004 229842
rect 164344 221649 164372 231676
rect 164988 223582 165016 231676
rect 165160 224664 165212 224670
rect 165160 224606 165212 224612
rect 164976 223576 165028 223582
rect 164976 223518 165028 223524
rect 164330 221640 164386 221649
rect 164330 221575 164386 221584
rect 164148 220516 164200 220522
rect 164148 220458 164200 220464
rect 163320 219428 163372 219434
rect 163320 219370 163372 219376
rect 163964 219428 164016 219434
rect 163964 219370 164016 219376
rect 162308 218884 162360 218890
rect 162308 218826 162360 218832
rect 162492 218884 162544 218890
rect 162492 218826 162544 218832
rect 162504 217138 162532 218826
rect 163332 217138 163360 219370
rect 164160 217138 164188 220458
rect 165172 217274 165200 224606
rect 165632 224534 165660 231676
rect 166276 229770 166304 231676
rect 166552 231662 166934 231690
rect 167196 231662 167578 231690
rect 166264 229764 166316 229770
rect 166264 229706 166316 229712
rect 166552 227497 166580 231662
rect 166814 228848 166870 228857
rect 166814 228783 166816 228792
rect 166868 228783 166870 228792
rect 166816 228754 166868 228760
rect 166814 228440 166870 228449
rect 166814 228375 166816 228384
rect 166868 228375 166870 228384
rect 166954 228404 167006 228410
rect 166816 228346 166868 228352
rect 166954 228346 167006 228352
rect 166966 228290 166994 228346
rect 166828 228262 166994 228290
rect 166828 228177 166856 228262
rect 166814 228168 166870 228177
rect 166814 228103 166870 228112
rect 166538 227488 166594 227497
rect 166538 227423 166594 227432
rect 165620 224528 165672 224534
rect 165620 224470 165672 224476
rect 165988 224528 166040 224534
rect 165988 224470 166040 224476
rect 165620 222760 165672 222766
rect 165620 222702 165672 222708
rect 165632 218482 165660 222702
rect 165804 218748 165856 218754
rect 165804 218690 165856 218696
rect 165620 218476 165672 218482
rect 165620 218418 165672 218424
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217110 158392 217138
rect 159146 217110 159220 217138
rect 159974 217110 160048 217138
rect 160802 217110 160876 217138
rect 161630 217110 161704 217138
rect 162458 217110 162532 217138
rect 163286 217110 163360 217138
rect 164114 217110 164188 217138
rect 164942 217246 165200 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217110
rect 159146 216988 159174 217110
rect 159974 216988 160002 217110
rect 160802 216988 160830 217110
rect 161630 216988 161658 217110
rect 162458 216988 162486 217110
rect 163286 216988 163314 217110
rect 164114 216988 164142 217110
rect 164942 216988 164970 217246
rect 165816 217138 165844 218690
rect 166000 218210 166028 224470
rect 167196 222018 167224 231662
rect 168208 224806 168236 231676
rect 168852 231198 168880 231676
rect 169128 231662 169510 231690
rect 169864 231662 170154 231690
rect 170324 231662 170798 231690
rect 168840 231192 168892 231198
rect 168840 231134 168892 231140
rect 169128 228857 169156 231662
rect 169298 228984 169354 228993
rect 169298 228919 169300 228928
rect 169352 228919 169354 228928
rect 169300 228890 169352 228896
rect 169114 228848 169170 228857
rect 169114 228783 169170 228792
rect 169482 227352 169538 227361
rect 169482 227287 169484 227296
rect 169536 227287 169538 227296
rect 169484 227258 169536 227264
rect 169668 225888 169720 225894
rect 169668 225830 169720 225836
rect 168196 224800 168248 224806
rect 168196 224742 168248 224748
rect 168012 224256 168064 224262
rect 168012 224198 168064 224204
rect 167184 222012 167236 222018
rect 167184 221954 167236 221960
rect 167460 222012 167512 222018
rect 167460 221954 167512 221960
rect 167472 221746 167500 221954
rect 167460 221740 167512 221746
rect 167460 221682 167512 221688
rect 167644 221740 167696 221746
rect 167644 221682 167696 221688
rect 167656 221202 167684 221682
rect 167828 221604 167880 221610
rect 167828 221546 167880 221552
rect 167840 221202 167868 221546
rect 167644 221196 167696 221202
rect 167644 221138 167696 221144
rect 167828 221196 167880 221202
rect 167828 221138 167880 221144
rect 166736 221054 167132 221082
rect 166736 220969 166764 221054
rect 166722 220960 166778 220969
rect 166722 220895 166778 220904
rect 166906 220960 166962 220969
rect 167104 220930 167132 221054
rect 166906 220895 166962 220904
rect 167092 220924 167144 220930
rect 166448 220788 166500 220794
rect 166920 220776 166948 220895
rect 167092 220866 167144 220872
rect 166500 220748 166948 220776
rect 167184 220788 167236 220794
rect 166448 220730 166500 220736
rect 167184 220730 167236 220736
rect 167196 220674 167224 220730
rect 166460 220658 167224 220674
rect 166448 220652 167224 220658
rect 166500 220646 167224 220652
rect 166448 220594 166500 220600
rect 166908 220516 166960 220522
rect 166908 220458 166960 220464
rect 167092 220516 167144 220522
rect 167092 220458 167144 220464
rect 166920 220289 166948 220458
rect 167104 220289 167132 220458
rect 166906 220280 166962 220289
rect 166906 220215 166962 220224
rect 167090 220280 167146 220289
rect 167090 220215 167146 220224
rect 167460 219292 167512 219298
rect 167460 219234 167512 219240
rect 166632 218476 166684 218482
rect 166632 218418 166684 218424
rect 165988 218204 166040 218210
rect 165988 218146 166040 218152
rect 166644 217138 166672 218418
rect 167472 217138 167500 219234
rect 168024 217274 168052 224198
rect 168196 221740 168248 221746
rect 168196 221682 168248 221688
rect 168208 219298 168236 221682
rect 169680 219298 169708 225830
rect 169864 221882 169892 231662
rect 169852 221876 169904 221882
rect 169852 221818 169904 221824
rect 168196 219292 168248 219298
rect 168196 219234 168248 219240
rect 169116 219292 169168 219298
rect 169116 219234 169168 219240
rect 169668 219292 169720 219298
rect 169668 219234 169720 219240
rect 169944 219292 169996 219298
rect 169944 219234 169996 219240
rect 168024 217246 168282 217274
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217246
rect 169128 217138 169156 219234
rect 169956 217138 169984 219234
rect 170324 217326 170352 231662
rect 171048 229764 171100 229770
rect 171048 229706 171100 229712
rect 171060 219298 171088 229706
rect 171230 227624 171286 227633
rect 171230 227559 171286 227568
rect 171244 227458 171272 227559
rect 171232 227452 171284 227458
rect 171232 227394 171284 227400
rect 171428 226930 171456 231676
rect 171704 231662 172086 231690
rect 171704 227361 171732 231662
rect 172150 228984 172206 228993
rect 172150 228919 172206 228928
rect 172336 228948 172388 228954
rect 172164 228818 172192 228919
rect 172336 228890 172388 228896
rect 172152 228812 172204 228818
rect 172152 228754 172204 228760
rect 172348 228449 172376 228890
rect 172334 228440 172390 228449
rect 172334 228375 172390 228384
rect 172150 227624 172206 227633
rect 172150 227559 172206 227568
rect 172164 227458 172192 227559
rect 172152 227452 172204 227458
rect 172152 227394 172204 227400
rect 171690 227352 171746 227361
rect 171690 227287 171746 227296
rect 171600 227180 171652 227186
rect 171600 227122 171652 227128
rect 171244 226902 171456 226930
rect 171048 219292 171100 219298
rect 171048 219234 171100 219240
rect 171046 218648 171102 218657
rect 171046 218583 171048 218592
rect 171100 218583 171102 218592
rect 171048 218554 171100 218560
rect 170772 218068 170824 218074
rect 170772 218010 170824 218016
rect 170312 217320 170364 217326
rect 170312 217262 170364 217268
rect 170784 217138 170812 218010
rect 171244 217462 171272 226902
rect 171612 225894 171640 227122
rect 171600 225888 171652 225894
rect 171600 225830 171652 225836
rect 171784 225888 171836 225894
rect 171784 225830 171836 225836
rect 171796 224954 171824 225830
rect 171428 224926 171824 224954
rect 171428 218210 171456 224926
rect 171968 224800 172020 224806
rect 171968 224742 172020 224748
rect 171784 223576 171836 223582
rect 171784 223518 171836 223524
rect 171796 222902 171824 223518
rect 171784 222896 171836 222902
rect 171784 222838 171836 222844
rect 171600 218884 171652 218890
rect 171600 218826 171652 218832
rect 171612 218618 171640 218826
rect 171600 218612 171652 218618
rect 171600 218554 171652 218560
rect 171416 218204 171468 218210
rect 171416 218146 171468 218152
rect 171232 217456 171284 217462
rect 171232 217398 171284 217404
rect 171980 217274 172008 224742
rect 172716 222018 172744 231676
rect 172992 231662 173374 231690
rect 172992 224942 173020 231662
rect 174004 230654 174032 231676
rect 173992 230648 174044 230654
rect 173992 230590 174044 230596
rect 173162 228848 173218 228857
rect 174648 228818 174676 231676
rect 175306 231662 175504 231690
rect 174818 228848 174874 228857
rect 173162 228783 173218 228792
rect 174636 228812 174688 228818
rect 172980 224936 173032 224942
rect 172980 224878 173032 224884
rect 172888 222896 172940 222902
rect 172888 222838 172940 222844
rect 172704 222012 172756 222018
rect 172704 221954 172756 221960
rect 172428 219292 172480 219298
rect 172428 219234 172480 219240
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217110 170812 217138
rect 171566 217246 172008 217274
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217110
rect 171566 216988 171594 217246
rect 172440 217138 172468 219234
rect 172900 218657 172928 222838
rect 173176 219298 173204 228783
rect 174818 228783 174820 228792
rect 174636 228754 174688 228760
rect 174872 228783 174874 228792
rect 174820 228754 174872 228760
rect 174084 221876 174136 221882
rect 174084 221818 174136 221824
rect 173164 219292 173216 219298
rect 173164 219234 173216 219240
rect 172886 218648 172942 218657
rect 172886 218583 172942 218592
rect 173256 218204 173308 218210
rect 173256 218146 173308 218152
rect 173268 217138 173296 218146
rect 174096 217138 174124 221818
rect 174912 221740 174964 221746
rect 174912 221682 174964 221688
rect 174924 217138 174952 221682
rect 175476 220969 175504 231662
rect 175936 223446 175964 231676
rect 176488 231662 176594 231690
rect 176488 224954 176516 231662
rect 176752 230172 176804 230178
rect 176752 230114 176804 230120
rect 176764 229094 176792 230114
rect 176120 224926 176516 224954
rect 176672 229066 176792 229094
rect 175924 223440 175976 223446
rect 175924 223382 175976 223388
rect 176120 223174 176148 224926
rect 176672 223530 176700 229066
rect 177224 227458 177252 231676
rect 177408 231662 177882 231690
rect 177212 227452 177264 227458
rect 177212 227394 177264 227400
rect 177408 225026 177436 231662
rect 176304 223502 176700 223530
rect 177316 224998 177436 225026
rect 176108 223168 176160 223174
rect 176108 223110 176160 223116
rect 175462 220960 175518 220969
rect 175462 220895 175518 220904
rect 175740 218748 175792 218754
rect 175740 218690 175792 218696
rect 175752 217138 175780 218690
rect 176304 217274 176332 223502
rect 177316 221377 177344 224998
rect 177488 224936 177540 224942
rect 177488 224878 177540 224884
rect 176474 221368 176530 221377
rect 176474 221303 176476 221312
rect 176528 221303 176530 221312
rect 177302 221368 177358 221377
rect 177302 221303 177358 221312
rect 176476 221274 176528 221280
rect 177304 221196 177356 221202
rect 177304 221138 177356 221144
rect 176474 220824 176530 220833
rect 176474 220759 176476 220768
rect 176528 220759 176530 220768
rect 176614 220788 176666 220794
rect 176476 220730 176528 220736
rect 176614 220730 176666 220736
rect 176626 220674 176654 220730
rect 176488 220646 176654 220674
rect 176488 218074 176516 220646
rect 176476 218068 176528 218074
rect 176476 218010 176528 218016
rect 177316 217274 177344 221138
rect 177500 219162 177528 224878
rect 178512 224126 178540 231676
rect 178788 231662 179170 231690
rect 178500 224120 178552 224126
rect 178500 224062 178552 224068
rect 178788 219434 178816 231662
rect 179800 229094 179828 231676
rect 179984 231662 180458 231690
rect 179984 229094 180012 231662
rect 179708 229066 179828 229094
rect 179892 229066 180012 229094
rect 179708 228954 179736 229066
rect 179696 228948 179748 228954
rect 179696 228890 179748 228896
rect 179328 224120 179380 224126
rect 179328 224062 179380 224068
rect 178420 219406 178816 219434
rect 177488 219156 177540 219162
rect 177488 219098 177540 219104
rect 178224 218068 178276 218074
rect 178224 218010 178276 218016
rect 176304 217246 176562 217274
rect 177316 217246 177390 217274
rect 172394 217110 172468 217138
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217110 174952 217138
rect 175706 217110 175780 217138
rect 172394 216988 172422 217110
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217110
rect 175706 216988 175734 217110
rect 176534 216988 176562 217246
rect 177362 216988 177390 217246
rect 178236 217138 178264 218010
rect 178420 217598 178448 219406
rect 179052 219156 179104 219162
rect 179052 219098 179104 219104
rect 178408 217592 178460 217598
rect 178408 217534 178460 217540
rect 179064 217138 179092 219098
rect 179340 218074 179368 224062
rect 179892 220833 179920 229066
rect 180064 228948 180116 228954
rect 180064 228890 180116 228896
rect 179878 220824 179934 220833
rect 179878 220759 179934 220768
rect 180076 218890 180104 228890
rect 181088 223990 181116 231676
rect 181352 227452 181404 227458
rect 181352 227394 181404 227400
rect 181076 223984 181128 223990
rect 181076 223926 181128 223932
rect 180524 220788 180576 220794
rect 180524 220730 180576 220736
rect 180708 220788 180760 220794
rect 180708 220730 180760 220736
rect 180536 220153 180564 220730
rect 180522 220144 180578 220153
rect 180522 220079 180578 220088
rect 180064 218884 180116 218890
rect 180064 218826 180116 218832
rect 179880 218204 179932 218210
rect 179880 218146 179932 218152
rect 179328 218068 179380 218074
rect 179328 218010 179380 218016
rect 179892 217138 179920 218146
rect 180720 217274 180748 220730
rect 181168 218748 181220 218754
rect 181168 218690 181220 218696
rect 181180 218346 181208 218690
rect 181364 218618 181392 227394
rect 181732 223582 181760 231676
rect 182376 227594 182404 231676
rect 182652 231662 183034 231690
rect 182364 227588 182416 227594
rect 182364 227530 182416 227536
rect 181720 223576 181772 223582
rect 181720 223518 181772 223524
rect 181996 223168 182048 223174
rect 181996 223110 182048 223116
rect 181352 218612 181404 218618
rect 181352 218554 181404 218560
rect 182008 218346 182036 223110
rect 182652 221610 182680 231662
rect 183664 223854 183692 231676
rect 184308 230790 184336 231676
rect 184296 230784 184348 230790
rect 184296 230726 184348 230732
rect 184664 229220 184716 229226
rect 184664 229162 184716 229168
rect 183652 223848 183704 223854
rect 183652 223790 183704 223796
rect 184388 223848 184440 223854
rect 184388 223790 184440 223796
rect 183192 223576 183244 223582
rect 183192 223518 183244 223524
rect 182640 221604 182692 221610
rect 182640 221546 182692 221552
rect 182364 219292 182416 219298
rect 182364 219234 182416 219240
rect 181168 218340 181220 218346
rect 181168 218282 181220 218288
rect 181536 218340 181588 218346
rect 181536 218282 181588 218288
rect 181996 218340 182048 218346
rect 181996 218282 182048 218288
rect 178190 217110 178264 217138
rect 179018 217110 179092 217138
rect 179846 217110 179920 217138
rect 180674 217246 180748 217274
rect 178190 216988 178218 217110
rect 179018 216988 179046 217110
rect 179846 216988 179874 217110
rect 180674 216988 180702 217246
rect 181548 217138 181576 218282
rect 182376 217138 182404 219234
rect 183204 217274 183232 223518
rect 184400 218754 184428 223790
rect 184676 223582 184704 229162
rect 184952 228274 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 184940 228268 184992 228274
rect 184940 228210 184992 228216
rect 184664 223576 184716 223582
rect 184664 223518 184716 223524
rect 184848 223440 184900 223446
rect 184848 223382 184900 223388
rect 184662 221776 184718 221785
rect 184662 221711 184718 221720
rect 184676 219434 184704 221711
rect 184676 219406 184796 219434
rect 184388 218748 184440 218754
rect 184388 218690 184440 218696
rect 184020 218340 184072 218346
rect 184020 218282 184072 218288
rect 181502 217110 181576 217138
rect 182330 217110 182404 217138
rect 183158 217246 183232 217274
rect 181502 216988 181530 217110
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 218282
rect 184768 217274 184796 219406
rect 184860 218362 184888 223382
rect 185136 219842 185164 231662
rect 185400 227588 185452 227594
rect 185400 227530 185452 227536
rect 185412 226914 185440 227530
rect 185584 227316 185636 227322
rect 185584 227258 185636 227264
rect 185596 226914 185624 227258
rect 185400 226908 185452 226914
rect 185400 226850 185452 226856
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185400 224528 185452 224534
rect 185400 224470 185452 224476
rect 185584 224528 185636 224534
rect 185584 224470 185636 224476
rect 185412 223990 185440 224470
rect 185596 224126 185624 224470
rect 185584 224120 185636 224126
rect 185584 224062 185636 224068
rect 185400 223984 185452 223990
rect 185400 223926 185452 223932
rect 185872 222154 185900 231662
rect 186136 227452 186188 227458
rect 186136 227394 186188 227400
rect 185860 222148 185912 222154
rect 185860 222090 185912 222096
rect 185766 221776 185822 221785
rect 185766 221711 185768 221720
rect 185820 221711 185822 221720
rect 185768 221682 185820 221688
rect 185860 221332 185912 221338
rect 185860 221274 185912 221280
rect 185872 221218 185900 221274
rect 185320 221202 185900 221218
rect 185308 221196 185900 221202
rect 185360 221190 185900 221196
rect 185308 221138 185360 221144
rect 185766 220144 185822 220153
rect 185766 220079 185822 220088
rect 185780 219978 185808 220079
rect 185768 219972 185820 219978
rect 185768 219914 185820 219920
rect 185124 219836 185176 219842
rect 185124 219778 185176 219784
rect 184860 218346 184980 218362
rect 186148 218346 186176 227394
rect 186884 223310 186912 231676
rect 187528 227730 187556 231676
rect 188172 230926 188200 231676
rect 188160 230920 188212 230926
rect 188160 230862 188212 230868
rect 187516 227724 187568 227730
rect 187516 227666 187568 227672
rect 187700 227724 187752 227730
rect 187700 227666 187752 227672
rect 187712 227458 187740 227666
rect 187700 227452 187752 227458
rect 187700 227394 187752 227400
rect 188816 223718 188844 231676
rect 189092 231662 189474 231690
rect 189092 229094 189120 231662
rect 189092 229066 189304 229094
rect 188804 223712 188856 223718
rect 188804 223654 188856 223660
rect 187332 223576 187384 223582
rect 187332 223518 187384 223524
rect 186872 223304 186924 223310
rect 186872 223246 186924 223252
rect 186504 218612 186556 218618
rect 186504 218554 186556 218560
rect 184860 218340 184992 218346
rect 184860 218334 184940 218340
rect 184940 218282 184992 218288
rect 185676 218340 185728 218346
rect 185676 218282 185728 218288
rect 186136 218340 186188 218346
rect 186136 218282 186188 218288
rect 184768 217246 184842 217274
rect 183986 217110 184060 217138
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218282
rect 186516 217138 186544 218554
rect 187344 217138 187372 223518
rect 188160 223304 188212 223310
rect 188160 223246 188212 223252
rect 188172 217138 188200 223246
rect 188988 218884 189040 218890
rect 188988 218826 189040 218832
rect 189000 217138 189028 218826
rect 189276 217734 189304 229066
rect 189724 228268 189776 228274
rect 189724 228210 189776 228216
rect 189736 219298 189764 228210
rect 190104 228138 190132 231676
rect 190656 231662 190762 231690
rect 190656 229094 190684 231662
rect 190472 229066 190684 229094
rect 190092 228132 190144 228138
rect 190092 228074 190144 228080
rect 189908 227452 189960 227458
rect 189908 227394 189960 227400
rect 189724 219292 189776 219298
rect 189724 219234 189776 219240
rect 189920 219178 189948 227394
rect 190472 219858 190500 229066
rect 191392 222630 191420 231676
rect 191564 223712 191616 223718
rect 191564 223654 191616 223660
rect 191380 222624 191432 222630
rect 191380 222566 191432 222572
rect 190644 219972 190696 219978
rect 190644 219914 190696 219920
rect 190104 219842 190500 219858
rect 190092 219836 190500 219842
rect 190144 219830 190500 219836
rect 190092 219778 190144 219784
rect 189644 219150 189948 219178
rect 189644 218754 189672 219150
rect 189632 218748 189684 218754
rect 189632 218690 189684 218696
rect 189816 218748 189868 218754
rect 189816 218690 189868 218696
rect 189264 217728 189316 217734
rect 189264 217670 189316 217676
rect 189828 217138 189856 218690
rect 190656 217138 190684 219914
rect 191576 217274 191604 223654
rect 192036 222766 192064 231676
rect 192680 227594 192708 231676
rect 192944 228132 192996 228138
rect 192944 228074 192996 228080
rect 192668 227588 192720 227594
rect 192668 227530 192720 227536
rect 192024 222760 192076 222766
rect 192024 222702 192076 222708
rect 192956 219298 192984 228074
rect 193324 221066 193352 231676
rect 193968 226302 193996 231676
rect 193956 226296 194008 226302
rect 193956 226238 194008 226244
rect 194140 226296 194192 226302
rect 194140 226238 194192 226244
rect 193956 222760 194008 222766
rect 193956 222702 194008 222708
rect 193312 221060 193364 221066
rect 193312 221002 193364 221008
rect 192300 219292 192352 219298
rect 192300 219234 192352 219240
rect 192944 219292 192996 219298
rect 192944 219234 192996 219240
rect 193128 219292 193180 219298
rect 193128 219234 193180 219240
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217110 187372 217138
rect 188126 217110 188200 217138
rect 188954 217110 189028 217138
rect 189782 217110 189856 217138
rect 190610 217110 190684 217138
rect 191438 217246 191604 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217110
rect 188126 216988 188154 217110
rect 188954 216988 188982 217110
rect 189782 216988 189810 217110
rect 190610 216988 190638 217110
rect 191438 216988 191466 217246
rect 192312 217138 192340 219234
rect 193140 217138 193168 219234
rect 193968 217138 193996 222702
rect 194152 218890 194180 226238
rect 194612 223990 194640 231676
rect 195060 230648 195112 230654
rect 195060 230590 195112 230596
rect 195072 230042 195100 230590
rect 195060 230036 195112 230042
rect 195060 229978 195112 229984
rect 195256 228002 195284 231676
rect 195900 231062 195928 231676
rect 196176 231662 196558 231690
rect 196912 231662 197202 231690
rect 197464 231662 197846 231690
rect 198016 231662 198490 231690
rect 195888 231056 195940 231062
rect 195888 230998 195940 231004
rect 195428 230036 195480 230042
rect 195428 229978 195480 229984
rect 195244 227996 195296 228002
rect 195244 227938 195296 227944
rect 194784 224120 194836 224126
rect 194784 224062 194836 224068
rect 194600 223984 194652 223990
rect 194600 223926 194652 223932
rect 194140 218884 194192 218890
rect 194140 218826 194192 218832
rect 194324 218884 194376 218890
rect 194324 218826 194376 218832
rect 194336 218618 194364 218826
rect 194324 218612 194376 218618
rect 194324 218554 194376 218560
rect 194796 217138 194824 224062
rect 194968 223984 195020 223990
rect 194968 223926 195020 223932
rect 194980 223718 195008 223926
rect 194968 223712 195020 223718
rect 194968 223654 195020 223660
rect 195440 218754 195468 229978
rect 196176 225486 196204 231662
rect 196912 230654 196940 231662
rect 196900 230648 196952 230654
rect 196900 230590 196952 230596
rect 197464 226778 197492 231662
rect 198016 229094 198044 231662
rect 197740 229066 198044 229094
rect 197452 226772 197504 226778
rect 197452 226714 197504 226720
rect 196624 226024 196676 226030
rect 196624 225966 196676 225972
rect 196164 225480 196216 225486
rect 196164 225422 196216 225428
rect 196636 219162 196664 225966
rect 197176 222624 197228 222630
rect 197176 222566 197228 222572
rect 196624 219156 196676 219162
rect 196624 219098 196676 219104
rect 195428 218748 195480 218754
rect 195428 218690 195480 218696
rect 195612 218748 195664 218754
rect 195612 218690 195664 218696
rect 195624 217138 195652 218690
rect 196440 218340 196492 218346
rect 196440 218282 196492 218288
rect 196452 217138 196480 218282
rect 197188 217274 197216 222566
rect 197740 217870 197768 229066
rect 198004 225480 198056 225486
rect 198004 225422 198056 225428
rect 198016 218754 198044 225422
rect 199120 225350 199148 231676
rect 199108 225344 199160 225350
rect 199108 225286 199160 225292
rect 199764 224942 199792 231676
rect 200408 227866 200436 231676
rect 200592 231662 201066 231690
rect 200592 229094 200620 231662
rect 200592 229066 200804 229094
rect 200396 227860 200448 227866
rect 200396 227802 200448 227808
rect 200028 227724 200080 227730
rect 200028 227666 200080 227672
rect 200040 225026 200068 227666
rect 200040 224998 200160 225026
rect 199752 224936 199804 224942
rect 199752 224878 199804 224884
rect 199936 224936 199988 224942
rect 199936 224878 199988 224884
rect 199948 224074 199976 224878
rect 200132 224754 200160 224998
rect 199856 224046 199976 224074
rect 200040 224726 200160 224754
rect 199856 223990 199884 224046
rect 199844 223984 199896 223990
rect 199844 223926 199896 223932
rect 200040 219298 200068 224726
rect 200396 222148 200448 222154
rect 200396 222090 200448 222096
rect 198188 219292 198240 219298
rect 198188 219234 198240 219240
rect 198924 219292 198976 219298
rect 198924 219234 198976 219240
rect 200028 219292 200080 219298
rect 200028 219234 200080 219240
rect 198200 218754 198228 219234
rect 198004 218748 198056 218754
rect 198004 218690 198056 218696
rect 198188 218748 198240 218754
rect 198188 218690 198240 218696
rect 198096 218612 198148 218618
rect 198096 218554 198148 218560
rect 197728 217864 197780 217870
rect 197728 217806 197780 217812
rect 197188 217246 197262 217274
rect 192266 217110 192340 217138
rect 193094 217110 193168 217138
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217110 195652 217138
rect 196406 217110 196480 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217110
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217110
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198108 217138 198136 218554
rect 198936 217138 198964 219234
rect 199752 219156 199804 219162
rect 199752 219098 199804 219104
rect 199764 217138 199792 219098
rect 200408 218618 200436 222090
rect 200776 219570 200804 229066
rect 201696 225078 201724 231676
rect 202340 230314 202368 231676
rect 202998 231662 203196 231690
rect 202328 230308 202380 230314
rect 202328 230250 202380 230256
rect 202420 228540 202472 228546
rect 202420 228482 202472 228488
rect 202432 228138 202460 228482
rect 202420 228132 202472 228138
rect 202420 228074 202472 228080
rect 203168 226642 203196 231662
rect 203628 230518 203656 231676
rect 203616 230512 203668 230518
rect 203616 230454 203668 230460
rect 203524 227860 203576 227866
rect 203524 227802 203576 227808
rect 203156 226636 203208 226642
rect 203156 226578 203208 226584
rect 202602 226264 202658 226273
rect 202602 226199 202658 226208
rect 201684 225072 201736 225078
rect 201684 225014 201736 225020
rect 201408 223984 201460 223990
rect 201408 223926 201460 223932
rect 201132 219700 201184 219706
rect 201132 219642 201184 219648
rect 200764 219564 200816 219570
rect 200764 219506 200816 219512
rect 201144 219434 201172 219642
rect 200592 219406 201172 219434
rect 200396 218612 200448 218618
rect 200396 218554 200448 218560
rect 200592 217274 200620 219406
rect 201420 217274 201448 223926
rect 202420 220380 202472 220386
rect 202420 220322 202472 220328
rect 202432 219881 202460 220322
rect 202418 219872 202474 219881
rect 202418 219807 202474 219816
rect 202616 219434 202644 226199
rect 203156 225616 203208 225622
rect 203156 225558 203208 225564
rect 203168 225350 203196 225558
rect 203156 225344 203208 225350
rect 203156 225286 203208 225292
rect 202788 220380 202840 220386
rect 202788 220322 202840 220328
rect 202800 219842 202828 220322
rect 203154 219872 203210 219881
rect 202788 219836 202840 219842
rect 203154 219807 203210 219816
rect 202788 219778 202840 219784
rect 203168 219706 203196 219807
rect 203156 219700 203208 219706
rect 203156 219642 203208 219648
rect 202616 219406 202828 219434
rect 201868 219292 201920 219298
rect 201868 219234 201920 219240
rect 201880 218482 201908 219234
rect 201868 218476 201920 218482
rect 201868 218418 201920 218424
rect 202800 218346 202828 219406
rect 203536 219026 203564 227802
rect 204076 227044 204128 227050
rect 204076 226986 204128 226992
rect 204088 226642 204116 226986
rect 204076 226636 204128 226642
rect 204076 226578 204128 226584
rect 204272 225214 204300 231676
rect 204916 229094 204944 231676
rect 204548 229066 204944 229094
rect 205560 229090 205588 231676
rect 205836 231662 206218 231690
rect 205548 229084 205600 229090
rect 204548 225894 204576 229066
rect 205548 229026 205600 229032
rect 205456 227860 205508 227866
rect 205456 227802 205508 227808
rect 204904 227724 204956 227730
rect 204904 227666 204956 227672
rect 204916 227458 204944 227666
rect 204720 227452 204772 227458
rect 204720 227394 204772 227400
rect 204904 227452 204956 227458
rect 204904 227394 204956 227400
rect 204732 226778 204760 227394
rect 204720 226772 204772 226778
rect 204720 226714 204772 226720
rect 204904 226296 204956 226302
rect 205088 226296 205140 226302
rect 204904 226238 204956 226244
rect 205086 226264 205088 226273
rect 205140 226264 205142 226273
rect 204916 225894 204944 226238
rect 205086 226199 205142 226208
rect 204536 225888 204588 225894
rect 204536 225830 204588 225836
rect 204904 225888 204956 225894
rect 204904 225830 204956 225836
rect 204904 225752 204956 225758
rect 204904 225694 204956 225700
rect 204916 225486 204944 225694
rect 204904 225480 204956 225486
rect 204904 225422 204956 225428
rect 204260 225208 204312 225214
rect 204260 225150 204312 225156
rect 204536 225208 204588 225214
rect 204536 225150 204588 225156
rect 203892 225072 203944 225078
rect 203892 225014 203944 225020
rect 203524 219020 203576 219026
rect 203524 218962 203576 218968
rect 203064 218612 203116 218618
rect 203064 218554 203116 218560
rect 202236 218340 202288 218346
rect 202236 218282 202288 218288
rect 202788 218340 202840 218346
rect 202788 218282 202840 218288
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217246 200620 217274
rect 201374 217246 201448 217274
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217246
rect 201374 216988 201402 217246
rect 202248 217138 202276 218282
rect 203076 217138 203104 218554
rect 203904 217274 203932 225014
rect 204548 219434 204576 225150
rect 204904 221468 204956 221474
rect 204904 221410 204956 221416
rect 205088 221468 205140 221474
rect 205088 221410 205140 221416
rect 204916 221202 204944 221410
rect 204904 221196 204956 221202
rect 204904 221138 204956 221144
rect 205100 221066 205128 221410
rect 205088 221060 205140 221066
rect 205088 221002 205140 221008
rect 204536 219428 204588 219434
rect 204536 219370 204588 219376
rect 204720 218340 204772 218346
rect 204720 218282 204772 218288
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218282
rect 205468 217274 205496 227802
rect 205836 219570 205864 231662
rect 206284 230444 206336 230450
rect 206284 230386 206336 230392
rect 206008 229084 206060 229090
rect 206008 229026 206060 229032
rect 206020 228002 206048 229026
rect 206008 227996 206060 228002
rect 206008 227938 206060 227944
rect 205824 219564 205876 219570
rect 205824 219506 205876 219512
rect 206296 219434 206324 230386
rect 206848 222494 206876 231676
rect 207492 223854 207520 231676
rect 208136 226642 208164 231676
rect 208596 231662 208794 231690
rect 208124 226636 208176 226642
rect 208124 226578 208176 226584
rect 207480 223848 207532 223854
rect 207480 223790 207532 223796
rect 207664 223712 207716 223718
rect 207664 223654 207716 223660
rect 206836 222488 206888 222494
rect 206836 222430 206888 222436
rect 207204 219700 207256 219706
rect 207204 219642 207256 219648
rect 206204 219406 206324 219434
rect 206204 218618 206232 219406
rect 206376 219020 206428 219026
rect 206376 218962 206428 218968
rect 206192 218612 206244 218618
rect 206192 218554 206244 218560
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206388 217138 206416 218962
rect 207216 217274 207244 219642
rect 207676 219298 207704 223654
rect 207848 222488 207900 222494
rect 207848 222430 207900 222436
rect 207664 219292 207716 219298
rect 207664 219234 207716 219240
rect 207860 218346 207888 222430
rect 208596 219570 208624 231662
rect 209424 225350 209452 231676
rect 210068 229498 210096 231676
rect 210424 230308 210476 230314
rect 210424 230250 210476 230256
rect 210056 229492 210108 229498
rect 210056 229434 210108 229440
rect 209596 225480 209648 225486
rect 209596 225422 209648 225428
rect 209412 225344 209464 225350
rect 209412 225286 209464 225292
rect 209608 219586 209636 225422
rect 208584 219564 208636 219570
rect 208584 219506 208636 219512
rect 209516 219558 209636 219586
rect 208032 218612 208084 218618
rect 208032 218554 208084 218560
rect 207848 218340 207900 218346
rect 207848 218282 207900 218288
rect 206342 217110 206416 217138
rect 207170 217246 207244 217274
rect 206342 216988 206370 217110
rect 207170 216988 207198 217246
rect 208044 217138 208072 218554
rect 209516 218346 209544 219558
rect 210436 219434 210464 230250
rect 210712 228138 210740 231676
rect 210700 228132 210752 228138
rect 210700 228074 210752 228080
rect 210976 227860 211028 227866
rect 210976 227802 211028 227808
rect 209688 219428 209740 219434
rect 209688 219370 209740 219376
rect 210424 219428 210476 219434
rect 210424 219370 210476 219376
rect 208860 218340 208912 218346
rect 208860 218282 208912 218288
rect 209504 218340 209556 218346
rect 209504 218282 209556 218288
rect 208872 217138 208900 218282
rect 209700 217138 209728 219370
rect 210332 218340 210384 218346
rect 210332 218282 210384 218288
rect 210344 218074 210372 218282
rect 210988 218074 211016 227802
rect 211356 221202 211384 231676
rect 212000 222358 212028 231676
rect 212172 226636 212224 226642
rect 212172 226578 212224 226584
rect 211988 222352 212040 222358
rect 211988 222294 212040 222300
rect 211344 221196 211396 221202
rect 211344 221138 211396 221144
rect 211528 221196 211580 221202
rect 211528 221138 211580 221144
rect 211344 219292 211396 219298
rect 211344 219234 211396 219240
rect 210332 218068 210384 218074
rect 210332 218010 210384 218016
rect 210516 218068 210568 218074
rect 210516 218010 210568 218016
rect 210976 218068 211028 218074
rect 210976 218010 211028 218016
rect 210528 217138 210556 218010
rect 211356 217138 211384 219234
rect 211540 218618 211568 221138
rect 211528 218612 211580 218618
rect 211528 218554 211580 218560
rect 212184 217274 212212 226578
rect 212644 222902 212672 231676
rect 213288 226506 213316 231676
rect 213946 231662 214144 231690
rect 214116 229094 214144 231662
rect 214116 229066 214236 229094
rect 213920 228132 213972 228138
rect 213920 228074 213972 228080
rect 213276 226500 213328 226506
rect 213276 226442 213328 226448
rect 213932 226250 213960 228074
rect 214208 227202 214236 229066
rect 214380 229084 214432 229090
rect 214380 229026 214432 229032
rect 214392 228682 214420 229026
rect 214380 228676 214432 228682
rect 214380 228618 214432 228624
rect 214576 228562 214604 231676
rect 214748 230036 214800 230042
rect 214748 229978 214800 229984
rect 214760 229634 214788 229978
rect 214748 229628 214800 229634
rect 214748 229570 214800 229576
rect 215220 229362 215248 231676
rect 215208 229356 215260 229362
rect 215208 229298 215260 229304
rect 214748 229084 214800 229090
rect 214748 229026 214800 229032
rect 214392 228534 214604 228562
rect 214392 228138 214420 228534
rect 214564 228404 214616 228410
rect 214564 228346 214616 228352
rect 214576 228138 214604 228346
rect 214380 228132 214432 228138
rect 214380 228074 214432 228080
rect 214564 228132 214616 228138
rect 214564 228074 214616 228080
rect 214760 228002 214788 229026
rect 215864 228546 215892 231676
rect 216048 231662 216522 231690
rect 215852 228540 215904 228546
rect 215852 228482 215904 228488
rect 214748 227996 214800 228002
rect 214748 227938 214800 227944
rect 214748 227588 214800 227594
rect 214748 227530 214800 227536
rect 214932 227588 214984 227594
rect 214932 227530 214984 227536
rect 214208 227174 214328 227202
rect 214104 227044 214156 227050
rect 214104 226986 214156 226992
rect 214116 226778 214144 226986
rect 214104 226772 214156 226778
rect 214104 226714 214156 226720
rect 213472 226222 213960 226250
rect 213472 226166 213500 226222
rect 213460 226160 213512 226166
rect 213460 226102 213512 226108
rect 213644 226160 213696 226166
rect 213644 226102 213696 226108
rect 213656 225894 213684 226102
rect 213644 225888 213696 225894
rect 213644 225830 213696 225836
rect 212632 222896 212684 222902
rect 212632 222838 212684 222844
rect 213184 222896 213236 222902
rect 213184 222838 213236 222844
rect 212908 220244 212960 220250
rect 212908 220186 212960 220192
rect 212920 219570 212948 220186
rect 212908 219564 212960 219570
rect 212908 219506 212960 219512
rect 213000 218476 213052 218482
rect 213000 218418 213052 218424
rect 207998 217110 208072 217138
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217110 210556 217138
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 207998 216988 208026 217110
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217110
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 218418
rect 213196 218346 213224 222838
rect 213828 220244 213880 220250
rect 213828 220186 213880 220192
rect 213184 218340 213236 218346
rect 213184 218282 213236 218288
rect 213840 217274 213868 220186
rect 214300 220114 214328 227174
rect 214760 226914 214788 227530
rect 214748 226908 214800 226914
rect 214748 226850 214800 226856
rect 214944 226642 214972 227530
rect 214932 226636 214984 226642
rect 214932 226578 214984 226584
rect 215208 225208 215260 225214
rect 215208 225150 215260 225156
rect 214564 220380 214616 220386
rect 214564 220322 214616 220328
rect 214576 220114 214604 220322
rect 214288 220108 214340 220114
rect 214288 220050 214340 220056
rect 214564 220108 214616 220114
rect 214564 220050 214616 220056
rect 215220 218074 215248 225150
rect 216048 224954 216076 231662
rect 216220 228540 216272 228546
rect 216220 228482 216272 228488
rect 216232 224954 216260 228482
rect 216404 226500 216456 226506
rect 216404 226442 216456 226448
rect 216416 224954 216444 226442
rect 217152 225622 217180 231676
rect 217508 228404 217560 228410
rect 217508 228346 217560 228352
rect 217140 225616 217192 225622
rect 217140 225558 217192 225564
rect 215956 224926 216076 224954
rect 216140 224926 216260 224954
rect 216324 224926 216444 224954
rect 215956 219570 215984 224926
rect 215944 219564 215996 219570
rect 215944 219506 215996 219512
rect 216140 218074 216168 224926
rect 214656 218068 214708 218074
rect 214656 218010 214708 218016
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 216128 218068 216180 218074
rect 216128 218010 216180 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 218010
rect 215496 217138 215524 218010
rect 216324 217274 216352 224926
rect 217140 220244 217192 220250
rect 217140 220186 217192 220192
rect 217152 217274 217180 220186
rect 217520 219434 217548 228346
rect 217796 227730 217824 231676
rect 217784 227724 217836 227730
rect 217784 227666 217836 227672
rect 218440 226778 218468 231676
rect 218428 226772 218480 226778
rect 218428 226714 218480 226720
rect 217876 225616 217928 225622
rect 217876 225558 217928 225564
rect 217888 225214 217916 225558
rect 217876 225208 217928 225214
rect 217876 225150 217928 225156
rect 219084 223038 219112 231676
rect 219742 231662 220216 231690
rect 219992 230036 220044 230042
rect 219992 229978 220044 229984
rect 220004 229770 220032 229978
rect 219992 229764 220044 229770
rect 219992 229706 220044 229712
rect 219808 228812 219860 228818
rect 219808 228754 219860 228760
rect 219622 228712 219678 228721
rect 219622 228647 219678 228656
rect 219636 228546 219664 228647
rect 219624 228540 219676 228546
rect 219624 228482 219676 228488
rect 219820 228138 219848 228754
rect 219992 228540 220044 228546
rect 219992 228482 220044 228488
rect 219808 228132 219860 228138
rect 219808 228074 219860 228080
rect 220004 227866 220032 228482
rect 219992 227860 220044 227866
rect 219992 227802 220044 227808
rect 219808 227724 219860 227730
rect 219808 227666 219860 227672
rect 219532 227316 219584 227322
rect 219532 227258 219584 227264
rect 219348 226772 219400 226778
rect 219348 226714 219400 226720
rect 219072 223032 219124 223038
rect 219072 222974 219124 222980
rect 218152 221060 218204 221066
rect 218152 221002 218204 221008
rect 217336 219406 217548 219434
rect 217968 219428 218020 219434
rect 217336 218618 217364 219406
rect 217968 219370 218020 219376
rect 217324 218612 217376 218618
rect 217324 218554 217376 218560
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217246 216352 217274
rect 217106 217246 217180 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217246
rect 217106 216988 217134 217246
rect 217980 217138 218008 219370
rect 218164 219298 218192 221002
rect 218152 219292 218204 219298
rect 218152 219234 218204 219240
rect 219360 218074 219388 226714
rect 219544 226642 219572 227258
rect 219820 227186 219848 227666
rect 219992 227316 220044 227322
rect 219992 227258 220044 227264
rect 219808 227180 219860 227186
rect 219808 227122 219860 227128
rect 220004 226914 220032 227258
rect 219992 226908 220044 226914
rect 219992 226850 220044 226856
rect 219532 226636 219584 226642
rect 219532 226578 219584 226584
rect 219992 226160 220044 226166
rect 219992 226102 220044 226108
rect 220004 225894 220032 226102
rect 219992 225888 220044 225894
rect 219992 225830 220044 225836
rect 220188 221474 220216 231662
rect 220372 229498 220400 231676
rect 220360 229492 220412 229498
rect 220360 229434 220412 229440
rect 220728 229492 220780 229498
rect 220728 229434 220780 229440
rect 220360 228948 220412 228954
rect 220360 228890 220412 228896
rect 220372 228682 220400 228890
rect 220542 228712 220598 228721
rect 220360 228676 220412 228682
rect 220542 228647 220544 228656
rect 220360 228618 220412 228624
rect 220596 228647 220598 228656
rect 220544 228618 220596 228624
rect 220740 226624 220768 229434
rect 221016 228002 221044 231676
rect 221292 231662 221674 231690
rect 221004 227996 221056 228002
rect 221004 227938 221056 227944
rect 220556 226596 220768 226624
rect 220556 226506 220584 226596
rect 220544 226500 220596 226506
rect 220544 226442 220596 226448
rect 220728 226500 220780 226506
rect 220728 226442 220780 226448
rect 220176 221468 220228 221474
rect 220176 221410 220228 221416
rect 220740 219434 220768 226442
rect 221004 221468 221056 221474
rect 221004 221410 221056 221416
rect 221016 221066 221044 221410
rect 221004 221060 221056 221066
rect 221004 221002 221056 221008
rect 221292 220658 221320 231662
rect 221464 228404 221516 228410
rect 221464 228346 221516 228352
rect 221476 228002 221504 228346
rect 221464 227996 221516 228002
rect 221464 227938 221516 227944
rect 221832 227044 221884 227050
rect 221832 226986 221884 226992
rect 221280 220652 221332 220658
rect 221280 220594 221332 220600
rect 221648 219496 221700 219502
rect 221648 219438 221700 219444
rect 220464 219406 220768 219434
rect 219624 218612 219676 218618
rect 219624 218554 219676 218560
rect 218796 218068 218848 218074
rect 218796 218010 218848 218016
rect 219348 218068 219400 218074
rect 219348 218010 219400 218016
rect 218808 217138 218836 218010
rect 219636 217138 219664 218554
rect 220464 217274 220492 219406
rect 221660 218482 221688 219438
rect 221648 218476 221700 218482
rect 221648 218418 221700 218424
rect 221844 218074 221872 226986
rect 222016 226160 222068 226166
rect 222016 226102 222068 226108
rect 221280 218068 221332 218074
rect 221280 218010 221332 218016
rect 221832 218068 221884 218074
rect 221832 218010 221884 218016
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218010
rect 222028 217274 222056 226102
rect 222304 220930 222332 231676
rect 222948 225350 222976 231676
rect 223592 226642 223620 231676
rect 223776 231662 224250 231690
rect 223580 226636 223632 226642
rect 223580 226578 223632 226584
rect 222936 225344 222988 225350
rect 222936 225286 222988 225292
rect 223488 221060 223540 221066
rect 223488 221002 223540 221008
rect 222292 220924 222344 220930
rect 222292 220866 222344 220872
rect 223500 219298 223528 221002
rect 223776 220658 223804 231662
rect 224592 228404 224644 228410
rect 224592 228346 224644 228352
rect 223764 220652 223816 220658
rect 223764 220594 223816 220600
rect 223764 220516 223816 220522
rect 223764 220458 223816 220464
rect 223488 219292 223540 219298
rect 223488 219234 223540 219240
rect 222936 218340 222988 218346
rect 222936 218282 222988 218288
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218282
rect 223776 217274 223804 220458
rect 224604 217274 224632 228346
rect 224880 224398 224908 231676
rect 225524 229906 225552 231676
rect 225512 229900 225564 229906
rect 225512 229842 225564 229848
rect 226168 228818 226196 231676
rect 226536 231662 226826 231690
rect 226156 228812 226208 228818
rect 226156 228754 226208 228760
rect 226156 227860 226208 227866
rect 226156 227802 226208 227808
rect 225604 226636 225656 226642
rect 225604 226578 225656 226584
rect 224868 224392 224920 224398
rect 224868 224334 224920 224340
rect 225616 218210 225644 226578
rect 225972 218476 226024 218482
rect 225972 218418 226024 218424
rect 225604 218204 225656 218210
rect 225604 218146 225656 218152
rect 225420 218068 225472 218074
rect 225420 218010 225472 218016
rect 222902 217110 222976 217138
rect 223730 217246 223804 217274
rect 224558 217246 224632 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217246
rect 224558 216988 224586 217246
rect 225432 217138 225460 218010
rect 225984 217274 226012 218418
rect 226168 218074 226196 227802
rect 226536 222018 226564 231662
rect 227456 224670 227484 231676
rect 227444 224664 227496 224670
rect 227444 224606 227496 224612
rect 227536 223848 227588 223854
rect 227536 223790 227588 223796
rect 226524 222012 226576 222018
rect 226524 221954 226576 221960
rect 227548 218074 227576 223790
rect 228100 223718 228128 231676
rect 228744 227730 228772 231676
rect 229296 231662 229402 231690
rect 228732 227724 228784 227730
rect 228732 227666 228784 227672
rect 228916 227724 228968 227730
rect 228916 227666 228968 227672
rect 228928 226506 228956 227666
rect 228916 226500 228968 226506
rect 228916 226442 228968 226448
rect 228732 224664 228784 224670
rect 228732 224606 228784 224612
rect 228088 223712 228140 223718
rect 228088 223654 228140 223660
rect 227904 220924 227956 220930
rect 227904 220866 227956 220872
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227076 218068 227128 218074
rect 227076 218010 227128 218016
rect 227536 218068 227588 218074
rect 227536 218010 227588 218016
rect 225984 217246 226242 217274
rect 225386 217110 225460 217138
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227088 217138 227116 218010
rect 227916 217274 227944 220866
rect 228744 217274 228772 224606
rect 229296 220114 229324 231662
rect 230032 224262 230060 231676
rect 230676 230042 230704 231676
rect 230664 230036 230716 230042
rect 230664 229978 230716 229984
rect 230480 229900 230532 229906
rect 230480 229842 230532 229848
rect 230020 224256 230072 224262
rect 230492 224210 230520 229842
rect 231124 229492 231176 229498
rect 231124 229434 231176 229440
rect 230020 224198 230072 224204
rect 230400 224182 230520 224210
rect 229284 220108 229336 220114
rect 229284 220050 229336 220056
rect 230204 220108 230256 220114
rect 230204 220050 230256 220056
rect 230216 219434 230244 220050
rect 230216 219406 230336 219434
rect 229560 218068 229612 218074
rect 229560 218010 229612 218016
rect 227042 217110 227116 217138
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 227042 216988 227070 217110
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 218010
rect 230308 217274 230336 219406
rect 230400 218090 230428 224182
rect 231136 219434 231164 229434
rect 231320 228138 231348 231676
rect 231308 228132 231360 228138
rect 231308 228074 231360 228080
rect 231676 224256 231728 224262
rect 231676 224198 231728 224204
rect 231044 219406 231164 219434
rect 231044 218346 231072 219406
rect 231032 218340 231084 218346
rect 231032 218282 231084 218288
rect 230400 218074 230520 218090
rect 231688 218074 231716 224198
rect 231964 221882 231992 231676
rect 232608 224806 232636 231676
rect 233252 229094 233280 231676
rect 233896 229094 233924 231676
rect 233252 229066 233372 229094
rect 232596 224800 232648 224806
rect 232596 224742 232648 224748
rect 233148 224392 233200 224398
rect 233148 224334 233200 224340
rect 232136 222012 232188 222018
rect 232136 221954 232188 221960
rect 231952 221876 232004 221882
rect 231952 221818 232004 221824
rect 232148 221610 232176 221954
rect 232136 221604 232188 221610
rect 232136 221546 232188 221552
rect 232872 218340 232924 218346
rect 232872 218282 232924 218288
rect 230400 218068 230532 218074
rect 230400 218062 230480 218068
rect 230480 218010 230532 218016
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 230308 217246 230382 217274
rect 229526 217110 229600 217138
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217138 232912 218282
rect 233160 218074 233188 224334
rect 233344 222902 233372 229066
rect 233712 229066 233924 229094
rect 234172 231662 234554 231690
rect 234724 231662 235198 231690
rect 234172 229094 234200 231662
rect 234172 229066 234292 229094
rect 233712 227186 233740 229066
rect 233884 228132 233936 228138
rect 233884 228074 233936 228080
rect 233896 227866 233924 228074
rect 233884 227860 233936 227866
rect 233884 227802 233936 227808
rect 233700 227180 233752 227186
rect 233700 227122 233752 227128
rect 233332 222896 233384 222902
rect 233332 222838 233384 222844
rect 233700 221876 233752 221882
rect 233700 221818 233752 221824
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233712 217274 233740 221818
rect 234068 221468 234120 221474
rect 234068 221410 234120 221416
rect 234080 220930 234108 221410
rect 234264 221338 234292 229066
rect 234528 222896 234580 222902
rect 234528 222838 234580 222844
rect 234252 221332 234304 221338
rect 234252 221274 234304 221280
rect 234068 220924 234120 220930
rect 234068 220866 234120 220872
rect 234540 217274 234568 222838
rect 234724 222018 234752 231662
rect 235828 230178 235856 231676
rect 235816 230172 235868 230178
rect 235816 230114 235868 230120
rect 235816 226772 235868 226778
rect 235816 226714 235868 226720
rect 234712 222012 234764 222018
rect 234712 221954 234764 221960
rect 235828 218074 235856 226714
rect 236472 226030 236500 231676
rect 236748 231662 237130 231690
rect 236460 226024 236512 226030
rect 236460 225966 236512 225972
rect 236748 220794 236776 231662
rect 237760 224534 237788 231676
rect 238404 226642 238432 231676
rect 238576 228812 238628 228818
rect 238576 228754 238628 228760
rect 238392 226636 238444 226642
rect 238392 226578 238444 226584
rect 237748 224528 237800 224534
rect 237748 224470 237800 224476
rect 237012 222352 237064 222358
rect 237012 222294 237064 222300
rect 236736 220788 236788 220794
rect 236736 220730 236788 220736
rect 236184 220652 236236 220658
rect 236184 220594 236236 220600
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235816 218068 235868 218074
rect 235816 218010 235868 218016
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217110 232912 217138
rect 233666 217246 233740 217274
rect 234494 217246 234568 217274
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217110
rect 233666 216988 233694 217246
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217274 236224 220594
rect 237024 217274 237052 222294
rect 237840 221332 237892 221338
rect 237840 221274 237892 221280
rect 237852 217274 237880 221274
rect 235322 217110 235396 217138
rect 236150 217246 236224 217274
rect 236978 217246 237052 217274
rect 237806 217246 237880 217274
rect 238588 217274 238616 228754
rect 239048 228274 239076 231676
rect 239036 228268 239088 228274
rect 239036 228210 239088 228216
rect 239312 227860 239364 227866
rect 239312 227802 239364 227808
rect 239324 218890 239352 227802
rect 239692 223446 239720 231676
rect 239680 223440 239732 223446
rect 239680 223382 239732 223388
rect 240336 223174 240364 231676
rect 240980 229226 241008 231676
rect 240968 229220 241020 229226
rect 240968 229162 241020 229168
rect 241624 227322 241652 231676
rect 241612 227316 241664 227322
rect 241612 227258 241664 227264
rect 241152 227180 241204 227186
rect 241152 227122 241204 227128
rect 240324 223168 240376 223174
rect 240324 223110 240376 223116
rect 239496 219292 239548 219298
rect 239496 219234 239548 219240
rect 239312 218884 239364 218890
rect 239312 218826 239364 218832
rect 238588 217246 238662 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217246
rect 236978 216988 237006 217246
rect 237806 216988 237834 217246
rect 238634 216988 238662 217246
rect 239508 217138 239536 219234
rect 240324 218068 240376 218074
rect 240324 218010 240376 218016
rect 240336 217138 240364 218010
rect 241164 217274 241192 227122
rect 242268 223582 242296 231676
rect 242926 231662 243124 231690
rect 242532 230036 242584 230042
rect 242532 229978 242584 229984
rect 242544 229094 242572 229978
rect 242544 229066 242756 229094
rect 242256 223576 242308 223582
rect 242256 223518 242308 223524
rect 241336 223168 241388 223174
rect 241336 223110 241388 223116
rect 241348 218074 241376 223110
rect 241980 218204 242032 218210
rect 241980 218146 242032 218152
rect 241336 218068 241388 218074
rect 241336 218010 241388 218016
rect 239462 217110 239536 217138
rect 240290 217110 240364 217138
rect 241118 217246 241192 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217110
rect 241118 216988 241146 217246
rect 241992 217138 242020 218146
rect 242728 217274 242756 229066
rect 242900 225344 242952 225350
rect 242820 225292 242900 225298
rect 242820 225286 242952 225292
rect 242820 225270 242940 225286
rect 242820 218226 242848 225270
rect 243096 221746 243124 231662
rect 243556 227866 243584 231676
rect 243544 227860 243596 227866
rect 243544 227802 243596 227808
rect 244200 225894 244228 231676
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 244188 225888 244240 225894
rect 244188 225830 244240 225836
rect 244096 223440 244148 223446
rect 244096 223382 244148 223388
rect 243084 221740 243136 221746
rect 243084 221682 243136 221688
rect 243728 221604 243780 221610
rect 243728 221546 243780 221552
rect 243740 221338 243768 221546
rect 243728 221332 243780 221338
rect 243728 221274 243780 221280
rect 243544 219156 243596 219162
rect 243544 219098 243596 219104
rect 242820 218210 242940 218226
rect 243556 218210 243584 219098
rect 242820 218204 242952 218210
rect 242820 218198 242900 218204
rect 242900 218146 242952 218152
rect 243544 218204 243596 218210
rect 243544 218146 243596 218152
rect 244108 218074 244136 223382
rect 244476 219978 244504 231662
rect 245120 223310 245148 231662
rect 246132 229770 246160 231676
rect 246120 229764 246172 229770
rect 246120 229706 246172 229712
rect 246488 229356 246540 229362
rect 246488 229298 246540 229304
rect 246304 227860 246356 227866
rect 246304 227802 246356 227808
rect 245476 224800 245528 224806
rect 245476 224742 245528 224748
rect 245108 223304 245160 223310
rect 245108 223246 245160 223252
rect 245292 223032 245344 223038
rect 245292 222974 245344 222980
rect 244464 219972 244516 219978
rect 244464 219914 244516 219920
rect 245304 218074 245332 222974
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244096 218068 244148 218074
rect 244096 218010 244148 218016
rect 244464 218068 244516 218074
rect 244464 218010 244516 218016
rect 245292 218068 245344 218074
rect 245292 218010 245344 218016
rect 242728 217246 242802 217274
rect 241946 217110 242020 217138
rect 241946 216988 241974 217110
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217138 244504 218010
rect 245488 217274 245516 224742
rect 246120 218884 246172 218890
rect 246120 218826 246172 218832
rect 243602 217110 243676 217138
rect 244430 217110 244504 217138
rect 245258 217246 245516 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246132 217138 246160 218826
rect 246316 218754 246344 227802
rect 246500 220658 246528 229298
rect 246776 228954 246804 231676
rect 246764 228948 246816 228954
rect 246764 228890 246816 228896
rect 247420 222766 247448 231676
rect 248064 224942 248092 231676
rect 248708 227866 248736 231676
rect 248984 231662 249366 231690
rect 248984 229094 249012 231662
rect 248892 229066 249012 229094
rect 248696 227860 248748 227866
rect 248696 227802 248748 227808
rect 248892 225758 248920 229066
rect 249064 227860 249116 227866
rect 249064 227802 249116 227808
rect 248880 225752 248932 225758
rect 248880 225694 248932 225700
rect 248052 224936 248104 224942
rect 248052 224878 248104 224884
rect 248328 224528 248380 224534
rect 248328 224470 248380 224476
rect 247408 222760 247460 222766
rect 247408 222702 247460 222708
rect 246488 220652 246540 220658
rect 246488 220594 246540 220600
rect 246948 220652 247000 220658
rect 246948 220594 247000 220600
rect 246304 218748 246356 218754
rect 246304 218690 246356 218696
rect 246960 217274 246988 220594
rect 248340 218074 248368 224470
rect 249076 218210 249104 227802
rect 249248 227316 249300 227322
rect 249248 227258 249300 227264
rect 249064 218204 249116 218210
rect 249064 218146 249116 218152
rect 249260 218074 249288 227258
rect 249432 223576 249484 223582
rect 249432 223518 249484 223524
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248328 218068 248380 218074
rect 248328 218010 248380 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 249248 218068 249300 218074
rect 249248 218010 249300 218016
rect 246086 217110 246160 217138
rect 246914 217246 246988 217274
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217274 249472 223518
rect 249996 222630 250024 231676
rect 250640 224126 250668 231676
rect 251284 228002 251312 231676
rect 251272 227996 251324 228002
rect 251272 227938 251324 227944
rect 251928 227458 251956 231676
rect 252586 231662 252784 231690
rect 251916 227452 251968 227458
rect 251916 227394 251968 227400
rect 252468 226024 252520 226030
rect 252468 225966 252520 225972
rect 251088 225752 251140 225758
rect 251088 225694 251140 225700
rect 250628 224120 250680 224126
rect 250628 224062 250680 224068
rect 250904 223304 250956 223310
rect 250904 223246 250956 223252
rect 249984 222624 250036 222630
rect 249984 222566 250036 222572
rect 250916 218074 250944 223246
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250904 218068 250956 218074
rect 250904 218010 250956 218016
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217246 249472 217274
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217246
rect 250272 217138 250300 218010
rect 251100 217274 251128 225694
rect 252480 218074 252508 225966
rect 252756 219842 252784 231662
rect 252940 231662 253230 231690
rect 252940 222154 252968 231662
rect 253860 227866 253888 231676
rect 253848 227860 253900 227866
rect 253848 227802 253900 227808
rect 254504 226302 254532 231676
rect 254952 228268 255004 228274
rect 254952 228210 255004 228216
rect 254492 226296 254544 226302
rect 254492 226238 254544 226244
rect 252928 222148 252980 222154
rect 252928 222090 252980 222096
rect 253848 220924 253900 220930
rect 253848 220866 253900 220872
rect 253572 219972 253624 219978
rect 253572 219914 253624 219920
rect 252744 219836 252796 219842
rect 252744 219778 252796 219784
rect 252744 218748 252796 218754
rect 252744 218690 252796 218696
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 250226 217110 250300 217138
rect 251054 217246 251128 217274
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218690
rect 253584 217274 253612 219914
rect 253860 219026 253888 220866
rect 254400 220788 254452 220794
rect 254400 220730 254452 220736
rect 253848 219020 253900 219026
rect 253848 218962 253900 218968
rect 254412 217274 254440 220730
rect 254964 219434 254992 228210
rect 255148 225078 255176 231676
rect 255136 225072 255188 225078
rect 255136 225014 255188 225020
rect 255792 223990 255820 231676
rect 256436 230450 256464 231676
rect 256424 230444 256476 230450
rect 256424 230386 256476 230392
rect 256516 229764 256568 229770
rect 256516 229706 256568 229712
rect 255780 223984 255832 223990
rect 255780 223926 255832 223932
rect 254964 219406 255176 219434
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 254366 217246 254440 217274
rect 255148 217274 255176 219406
rect 256528 218074 256556 229706
rect 257080 229090 257108 231676
rect 257264 231662 257738 231690
rect 257068 229084 257120 229090
rect 257068 229026 257120 229032
rect 257264 219706 257292 231662
rect 257528 229084 257580 229090
rect 257528 229026 257580 229032
rect 257252 219700 257304 219706
rect 257252 219642 257304 219648
rect 257540 218074 257568 229026
rect 257712 228948 257764 228954
rect 257712 228890 257764 228896
rect 256056 218068 256108 218074
rect 256056 218010 256108 218016
rect 256516 218068 256568 218074
rect 256516 218010 256568 218016
rect 256884 218068 256936 218074
rect 256884 218010 256936 218016
rect 257528 218068 257580 218074
rect 257528 218010 257580 218016
rect 255148 217246 255222 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254366 216988 254394 217246
rect 255194 216988 255222 217246
rect 256068 217138 256096 218010
rect 256896 217138 256924 218010
rect 257724 217274 257752 228890
rect 258368 222494 258396 231676
rect 258644 231662 259026 231690
rect 258356 222488 258408 222494
rect 258356 222430 258408 222436
rect 258080 222148 258132 222154
rect 258080 222090 258132 222096
rect 258092 219434 258120 222090
rect 258644 220930 258672 231662
rect 259368 226636 259420 226642
rect 259368 226578 259420 226584
rect 258632 220924 258684 220930
rect 258632 220866 258684 220872
rect 258080 219428 258132 219434
rect 258080 219370 258132 219376
rect 259184 219020 259236 219026
rect 259184 218962 259236 218968
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 256022 217110 256096 217138
rect 256850 217110 256924 217138
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217110
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259196 217274 259224 218962
rect 259380 218074 259408 226578
rect 259656 225486 259684 231676
rect 260300 228546 260328 231676
rect 260944 229094 260972 231676
rect 261588 230314 261616 231676
rect 261576 230308 261628 230314
rect 261576 230250 261628 230256
rect 260852 229066 260972 229094
rect 260288 228540 260340 228546
rect 260288 228482 260340 228488
rect 260656 226296 260708 226302
rect 260656 226238 260708 226244
rect 259644 225480 259696 225486
rect 259644 225422 259696 225428
rect 260668 219434 260696 226238
rect 260852 221202 260880 229066
rect 262232 227594 262260 231676
rect 262416 231662 262890 231690
rect 263152 231662 263534 231690
rect 263888 231662 264178 231690
rect 262220 227588 262272 227594
rect 262220 227530 262272 227536
rect 261852 225888 261904 225894
rect 261852 225830 261904 225836
rect 261024 222012 261076 222018
rect 261024 221954 261076 221960
rect 260840 221196 260892 221202
rect 260840 221138 260892 221144
rect 260668 219406 260788 219434
rect 260760 218074 260788 219406
rect 259368 218068 259420 218074
rect 259368 218010 259420 218016
rect 260196 218068 260248 218074
rect 260196 218010 260248 218016
rect 260748 218068 260800 218074
rect 260748 218010 260800 218016
rect 259196 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260208 217138 260236 218010
rect 261036 217274 261064 221954
rect 261864 217274 261892 225830
rect 262416 220386 262444 231662
rect 263152 221746 263180 231662
rect 263888 222154 263916 231662
rect 264244 230172 264296 230178
rect 264244 230114 264296 230120
rect 263876 222148 263928 222154
rect 263876 222090 263928 222096
rect 263140 221740 263192 221746
rect 263140 221682 263192 221688
rect 263508 221740 263560 221746
rect 263508 221682 263560 221688
rect 262404 220380 262456 220386
rect 262404 220322 262456 220328
rect 262680 220380 262732 220386
rect 262680 220322 262732 220328
rect 262692 217274 262720 220322
rect 263520 217274 263548 221682
rect 264256 220386 264284 230114
rect 264808 228682 264836 231676
rect 265176 231662 265466 231690
rect 264796 228676 264848 228682
rect 264796 228618 264848 228624
rect 264796 227452 264848 227458
rect 264796 227394 264848 227400
rect 264244 220380 264296 220386
rect 264244 220322 264296 220328
rect 264612 220380 264664 220386
rect 264612 220322 264664 220328
rect 264624 218618 264652 220322
rect 264612 218612 264664 218618
rect 264612 218554 264664 218560
rect 264808 218074 264836 227394
rect 265176 220250 265204 231662
rect 266096 225622 266124 231676
rect 266740 229634 266768 231676
rect 266728 229628 266780 229634
rect 266728 229570 266780 229576
rect 267384 226914 267412 231676
rect 268028 227730 268056 231676
rect 268212 231662 268686 231690
rect 268016 227724 268068 227730
rect 268016 227666 268068 227672
rect 267372 226908 267424 226914
rect 267372 226850 267424 226856
rect 266084 225616 266136 225622
rect 266084 225558 266136 225564
rect 267004 225616 267056 225622
rect 267004 225558 267056 225564
rect 266268 224120 266320 224126
rect 266268 224062 266320 224068
rect 265164 220244 265216 220250
rect 265164 220186 265216 220192
rect 265992 218612 266044 218618
rect 265992 218554 266044 218560
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 260162 217110 260236 217138
rect 260990 217246 261064 217274
rect 261818 217246 261892 217274
rect 262646 217246 262720 217274
rect 263474 217246 263548 217274
rect 260162 216988 260190 217110
rect 260990 216988 261018 217246
rect 261818 216988 261846 217246
rect 262646 216988 262674 217246
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217138 266032 218554
rect 266280 218074 266308 224062
rect 266820 221332 266872 221338
rect 266820 221274 266872 221280
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266832 217274 266860 221274
rect 267016 218482 267044 225558
rect 268212 221066 268240 231662
rect 268936 228540 268988 228546
rect 268936 228482 268988 228488
rect 268200 221060 268252 221066
rect 268200 221002 268252 221008
rect 267648 220244 267700 220250
rect 267648 220186 267700 220192
rect 267004 218476 267056 218482
rect 267004 218418 267056 218424
rect 267660 217274 267688 220186
rect 268948 218074 268976 228482
rect 269316 220386 269344 231676
rect 269960 226166 269988 231676
rect 269948 226160 270000 226166
rect 269948 226102 270000 226108
rect 270224 226160 270276 226166
rect 270224 226102 270276 226108
rect 270040 222148 270092 222154
rect 270040 222090 270092 222096
rect 269304 220380 269356 220386
rect 269304 220322 269356 220328
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 268936 218068 268988 218074
rect 268936 218010 268988 218016
rect 269304 218068 269356 218074
rect 269304 218010 269356 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217110 266032 217138
rect 266786 217246 266860 217274
rect 267614 217246 267688 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217110
rect 266786 216988 266814 217246
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218010
rect 270052 217274 270080 222090
rect 270236 218074 270264 226102
rect 270604 220522 270632 231676
rect 271248 227050 271276 231676
rect 271892 229498 271920 231676
rect 271880 229492 271932 229498
rect 271880 229434 271932 229440
rect 272536 228138 272564 231676
rect 272524 228132 272576 228138
rect 272524 228074 272576 228080
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 270592 220516 270644 220522
rect 270592 220458 270644 220464
rect 270776 219836 270828 219842
rect 270776 219778 270828 219784
rect 270788 218346 270816 219778
rect 270776 218340 270828 218346
rect 270776 218282 270828 218288
rect 270224 218068 270276 218074
rect 270224 218010 270276 218016
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 270052 217246 270126 217274
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272524 224936 272576 224942
rect 272524 224878 272576 224884
rect 272340 219156 272392 219162
rect 272340 219098 272392 219104
rect 272352 218618 272380 219098
rect 272340 218612 272392 218618
rect 272340 218554 272392 218560
rect 272536 218074 272564 224878
rect 273180 223854 273208 231676
rect 273824 228410 273852 231676
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274272 228404 274324 228410
rect 274272 228346 274324 228352
rect 273168 223848 273220 223854
rect 273168 223790 273220 223796
rect 273444 220380 273496 220386
rect 273444 220322 273496 220328
rect 272892 219428 272944 219434
rect 272892 219370 272944 219376
rect 272708 219292 272760 219298
rect 272708 219234 272760 219240
rect 272720 218618 272748 219234
rect 272708 218612 272760 218618
rect 272708 218554 272760 218560
rect 272524 218068 272576 218074
rect 272524 218010 272576 218016
rect 272904 217274 272932 219370
rect 273456 217274 273484 220322
rect 274284 217274 274312 228346
rect 274468 225622 274496 231676
rect 275112 229094 275140 231676
rect 274928 229066 275140 229094
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 274456 225616 274508 225622
rect 274456 225558 274508 225564
rect 274928 224670 274956 229066
rect 274916 224664 274968 224670
rect 274916 224606 274968 224612
rect 275100 224664 275152 224670
rect 275100 224606 275152 224612
rect 275112 217274 275140 224606
rect 275296 220114 275324 231662
rect 275652 230308 275704 230314
rect 275652 230250 275704 230256
rect 275664 229094 275692 230250
rect 275664 229066 275876 229094
rect 275284 220108 275336 220114
rect 275284 220050 275336 220056
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 272582 217246 272932 217274
rect 273410 217246 273484 217274
rect 274238 217246 274312 217274
rect 275066 217246 275140 217274
rect 275848 217274 275876 229066
rect 276124 221474 276152 231662
rect 276296 230444 276348 230450
rect 276296 230386 276348 230392
rect 276308 223582 276336 230386
rect 277044 229906 277072 231676
rect 277032 229900 277084 229906
rect 277032 229842 277084 229848
rect 277688 224398 277716 231676
rect 277964 231662 278346 231690
rect 277676 224392 277728 224398
rect 277676 224334 277728 224340
rect 276296 223576 276348 223582
rect 276296 223518 276348 223524
rect 277964 221882 277992 231662
rect 278412 225616 278464 225622
rect 278412 225558 278464 225564
rect 277952 221876 278004 221882
rect 277952 221818 278004 221824
rect 276112 221468 276164 221474
rect 276112 221410 276164 221416
rect 276756 220516 276808 220522
rect 276756 220458 276808 220464
rect 276768 217274 276796 220458
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272582 216988 272610 217246
rect 273410 216988 273438 217246
rect 274238 216988 274266 217246
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276722 217246 276796 217274
rect 276722 216988 276750 217246
rect 277596 217138 277624 218010
rect 278424 217274 278452 225558
rect 278976 224262 279004 231676
rect 279160 231662 279634 231690
rect 278964 224256 279016 224262
rect 278964 224198 279016 224204
rect 278596 223576 278648 223582
rect 278596 223518 278648 223524
rect 278608 218074 278636 223518
rect 279160 219842 279188 231662
rect 280264 226778 280292 231676
rect 280252 226772 280304 226778
rect 280252 226714 280304 226720
rect 279424 223916 279476 223922
rect 279424 223858 279476 223864
rect 279148 219836 279200 219842
rect 279148 219778 279200 219784
rect 279056 219156 279108 219162
rect 279056 219098 279108 219104
rect 279068 218890 279096 219098
rect 279056 218884 279108 218890
rect 279056 218826 279108 218832
rect 279240 218884 279292 218890
rect 279240 218826 279292 218832
rect 278596 218068 278648 218074
rect 278596 218010 278648 218016
rect 277550 217110 277624 217138
rect 278378 217246 278452 217274
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218826
rect 279436 218618 279464 223858
rect 280908 222358 280936 231676
rect 281356 227588 281408 227594
rect 281356 227530 281408 227536
rect 280896 222352 280948 222358
rect 280896 222294 280948 222300
rect 280068 221876 280120 221882
rect 280068 221818 280120 221824
rect 279424 218612 279476 218618
rect 279424 218554 279476 218560
rect 280080 217274 280108 221818
rect 281368 219434 281396 227530
rect 281552 222902 281580 231676
rect 282196 229362 282224 231676
rect 282552 229900 282604 229906
rect 282552 229842 282604 229848
rect 282184 229356 282236 229362
rect 282184 229298 282236 229304
rect 281540 222896 281592 222902
rect 281540 222838 281592 222844
rect 281368 219406 281488 219434
rect 281460 218074 281488 219406
rect 280896 218068 280948 218074
rect 280896 218010 280948 218016
rect 281448 218068 281500 218074
rect 281448 218010 281500 218016
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280908 217138 280936 218010
rect 281736 217138 281764 218010
rect 282564 217274 282592 229842
rect 282840 228818 282868 231676
rect 282828 228812 282880 228818
rect 282828 228754 282880 228760
rect 283484 223174 283512 231676
rect 283760 231662 284142 231690
rect 283472 223168 283524 223174
rect 283472 223110 283524 223116
rect 282736 222896 282788 222902
rect 282736 222838 282788 222844
rect 282748 218074 282776 222838
rect 283760 221610 283788 231662
rect 284772 223922 284800 231676
rect 285048 231662 285430 231690
rect 285048 225350 285076 231662
rect 285496 228676 285548 228682
rect 285496 228618 285548 228624
rect 285036 225344 285088 225350
rect 285036 225286 285088 225292
rect 284760 223916 284812 223922
rect 284760 223858 284812 223864
rect 284208 222760 284260 222766
rect 284208 222702 284260 222708
rect 283748 221604 283800 221610
rect 283748 221546 283800 221552
rect 284024 221468 284076 221474
rect 284024 221410 284076 221416
rect 284036 219434 284064 221410
rect 284036 219406 284156 219434
rect 282736 218068 282788 218074
rect 282736 218010 282788 218016
rect 283380 218068 283432 218074
rect 283380 218010 283432 218016
rect 280862 217110 280936 217138
rect 281690 217110 281764 217138
rect 282518 217246 282592 217274
rect 280862 216988 280890 217110
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283392 217138 283420 218010
rect 284128 217274 284156 219406
rect 284220 218090 284248 222702
rect 284220 218074 284340 218090
rect 285508 218074 285536 228618
rect 286060 223446 286088 231676
rect 286704 227186 286732 231676
rect 287348 230042 287376 231676
rect 287716 231662 288006 231690
rect 287336 230036 287388 230042
rect 287336 229978 287388 229984
rect 287520 230036 287572 230042
rect 287520 229978 287572 229984
rect 286692 227180 286744 227186
rect 286692 227122 286744 227128
rect 287532 226166 287560 229978
rect 287520 226160 287572 226166
rect 287520 226102 287572 226108
rect 287716 224806 287744 231662
rect 288072 226160 288124 226166
rect 288072 226102 288124 226108
rect 287704 224800 287756 224806
rect 287704 224742 287756 224748
rect 286324 224256 286376 224262
rect 286324 224198 286376 224204
rect 286048 223440 286100 223446
rect 286048 223382 286100 223388
rect 286336 219162 286364 224198
rect 286692 219836 286744 219842
rect 286692 219778 286744 219784
rect 286324 219156 286376 219162
rect 286324 219098 286376 219104
rect 285864 218884 285916 218890
rect 285864 218826 285916 218832
rect 284220 218068 284352 218074
rect 284220 218062 284300 218068
rect 284300 218010 284352 218016
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 283346 217110 283420 217138
rect 283346 216988 283374 217110
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 218826
rect 286704 217274 286732 219778
rect 288084 218074 288112 226102
rect 288256 223168 288308 223174
rect 288256 223110 288308 223116
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 288072 218068 288124 218074
rect 288072 218010 288124 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 223110
rect 288636 220658 288664 231676
rect 288992 223304 289044 223310
rect 288992 223246 289044 223252
rect 288624 220652 288676 220658
rect 288624 220594 288676 220600
rect 289004 218482 289032 223246
rect 289280 223038 289308 231676
rect 289636 224392 289688 224398
rect 289636 224334 289688 224340
rect 289268 223032 289320 223038
rect 289268 222974 289320 222980
rect 288992 218476 289044 218482
rect 288992 218418 289044 218424
rect 289648 218074 289676 224334
rect 289924 224262 289952 231676
rect 290568 227322 290596 231676
rect 291016 227724 291068 227730
rect 291016 227666 291068 227672
rect 290556 227316 290608 227322
rect 290556 227258 290608 227264
rect 289912 224256 289964 224262
rect 289912 224198 289964 224204
rect 290832 224256 290884 224262
rect 290832 224198 290884 224204
rect 289820 219564 289872 219570
rect 289820 219506 289872 219512
rect 289832 219298 289860 219506
rect 289820 219292 289872 219298
rect 289820 219234 289872 219240
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289636 218068 289688 218074
rect 289636 218010 289688 218016
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217138 290044 218010
rect 290844 217274 290872 224198
rect 291028 219434 291056 227666
rect 291212 223446 291240 231676
rect 291856 224534 291884 231676
rect 292500 230450 292528 231676
rect 292488 230444 292540 230450
rect 292488 230386 292540 230392
rect 293144 226030 293172 231676
rect 293328 231662 293802 231690
rect 293132 226024 293184 226030
rect 293132 225966 293184 225972
rect 291844 224528 291896 224534
rect 291844 224470 291896 224476
rect 291200 223440 291252 223446
rect 291200 223382 291252 223388
rect 291660 223032 291712 223038
rect 291660 222974 291712 222980
rect 291028 219406 291148 219434
rect 291120 218074 291148 219406
rect 291672 219026 291700 222974
rect 292488 220108 292540 220114
rect 292488 220050 292540 220056
rect 292028 219292 292080 219298
rect 292028 219234 292080 219240
rect 291660 219020 291712 219026
rect 291660 218962 291712 218968
rect 292040 218890 292068 219234
rect 292028 218884 292080 218890
rect 292028 218826 292080 218832
rect 291660 218748 291712 218754
rect 291660 218690 291712 218696
rect 291108 218068 291160 218074
rect 291108 218010 291160 218016
rect 291672 217274 291700 218690
rect 292500 217274 292528 220050
rect 293328 219978 293356 231662
rect 293776 227316 293828 227322
rect 293776 227258 293828 227264
rect 293316 219972 293368 219978
rect 293316 219914 293368 219920
rect 293788 218074 293816 227258
rect 294432 225758 294460 231676
rect 294420 225752 294472 225758
rect 294420 225694 294472 225700
rect 294880 224528 294932 224534
rect 294880 224470 294932 224476
rect 294892 219434 294920 224470
rect 295076 223310 295104 231676
rect 295720 228274 295748 231676
rect 296364 229090 296392 231676
rect 296824 231662 297022 231690
rect 296352 229084 296404 229090
rect 296352 229026 296404 229032
rect 296628 228812 296680 228818
rect 296628 228754 296680 228760
rect 295708 228268 295760 228274
rect 295708 228210 295760 228216
rect 296444 225752 296496 225758
rect 296444 225694 296496 225700
rect 295064 223304 295116 223310
rect 295064 223246 295116 223252
rect 296456 219434 296484 225694
rect 294892 219406 295012 219434
rect 296456 219406 296576 219434
rect 294144 218476 294196 218482
rect 294144 218418 294196 218424
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217246 290872 217274
rect 291626 217246 291700 217274
rect 292454 217246 292528 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217246
rect 291626 216988 291654 217246
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218418
rect 294984 217274 295012 219406
rect 295800 219156 295852 219162
rect 295800 219098 295852 219104
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 219098
rect 296548 217274 296576 219406
rect 296640 219178 296668 228754
rect 296824 220794 296852 231662
rect 297652 229770 297680 231676
rect 297640 229764 297692 229770
rect 297640 229706 297692 229712
rect 296996 229628 297048 229634
rect 296996 229570 297048 229576
rect 297008 224398 297036 229570
rect 298296 226642 298324 231676
rect 298284 226636 298336 226642
rect 298284 226578 298336 226584
rect 298940 226302 298968 231676
rect 299584 228954 299612 231676
rect 299572 228948 299624 228954
rect 299572 228890 299624 228896
rect 298928 226296 298980 226302
rect 298928 226238 298980 226244
rect 299388 226024 299440 226030
rect 299388 225966 299440 225972
rect 297364 225480 297416 225486
rect 297364 225422 297416 225428
rect 296996 224392 297048 224398
rect 296996 224334 297048 224340
rect 296812 220788 296864 220794
rect 296812 220730 296864 220736
rect 296640 219162 296760 219178
rect 296640 219156 296772 219162
rect 296640 219150 296720 219156
rect 296720 219098 296772 219104
rect 297376 219026 297404 225422
rect 299112 224392 299164 224398
rect 299112 224334 299164 224340
rect 297548 223372 297600 223378
rect 297548 223314 297600 223320
rect 297560 219434 297588 223314
rect 297548 219428 297600 219434
rect 297548 219370 297600 219376
rect 297364 219020 297416 219026
rect 297364 218962 297416 218968
rect 297456 218204 297508 218210
rect 297456 218146 297508 218152
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218146
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 298296 217138 298324 218010
rect 299124 217274 299152 224334
rect 299400 218074 299428 225966
rect 300228 223038 300256 231676
rect 300676 228948 300728 228954
rect 300676 228890 300728 228896
rect 300216 223032 300268 223038
rect 300216 222974 300268 222980
rect 300492 219156 300544 219162
rect 300492 219098 300544 219104
rect 299388 218068 299440 218074
rect 299388 218010 299440 218016
rect 299940 218068 299992 218074
rect 299940 218010 299992 218016
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217246 299152 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217246
rect 299952 217138 299980 218010
rect 300504 217274 300532 219098
rect 300688 218074 300716 228890
rect 300872 225894 300900 231676
rect 301056 231662 301530 231690
rect 301700 231662 302174 231690
rect 300860 225888 300912 225894
rect 300860 225830 300912 225836
rect 301056 221746 301084 231662
rect 301700 222018 301728 231662
rect 302804 230178 302832 231676
rect 302792 230172 302844 230178
rect 302792 230114 302844 230120
rect 302976 230172 303028 230178
rect 302976 230114 303028 230120
rect 302148 229084 302200 229090
rect 302148 229026 302200 229032
rect 301688 222012 301740 222018
rect 301688 221954 301740 221960
rect 301044 221740 301096 221746
rect 301044 221682 301096 221688
rect 302160 218074 302188 229026
rect 302424 221604 302476 221610
rect 302424 221546 302476 221552
rect 300676 218068 300728 218074
rect 300676 218010 300728 218016
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 300504 217246 300762 217274
rect 299906 217110 299980 217138
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218010
rect 302436 217274 302464 221546
rect 302988 219434 303016 230114
rect 303448 224126 303476 231676
rect 303816 231662 304106 231690
rect 303436 224120 303488 224126
rect 303436 224062 303488 224068
rect 303252 221740 303304 221746
rect 303252 221682 303304 221688
rect 302896 219406 303016 219434
rect 302896 218210 302924 219406
rect 302884 218204 302936 218210
rect 302884 218146 302936 218152
rect 303264 217274 303292 221682
rect 303816 221338 303844 231662
rect 304736 227458 304764 231676
rect 304724 227452 304776 227458
rect 304724 227394 304776 227400
rect 304264 224120 304316 224126
rect 304264 224062 304316 224068
rect 303804 221332 303856 221338
rect 303804 221274 303856 221280
rect 304080 219428 304132 219434
rect 304080 219370 304132 219376
rect 301562 217110 301636 217138
rect 302390 217246 302464 217274
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217246
rect 303218 216988 303246 217246
rect 304092 217138 304120 219370
rect 304276 218618 304304 224062
rect 305380 223378 305408 231676
rect 306024 228546 306052 231676
rect 306392 231662 306682 231690
rect 306852 231662 307326 231690
rect 306012 228540 306064 228546
rect 306012 228482 306064 228488
rect 306196 227180 306248 227186
rect 306196 227122 306248 227128
rect 305368 223372 305420 223378
rect 305368 223314 305420 223320
rect 304908 220652 304960 220658
rect 304908 220594 304960 220600
rect 304264 218612 304316 218618
rect 304264 218554 304316 218560
rect 304920 217274 304948 220594
rect 306208 218074 306236 227122
rect 306392 222154 306420 231662
rect 306380 222148 306432 222154
rect 306380 222090 306432 222096
rect 306852 220250 306880 231662
rect 307956 230042 307984 231676
rect 308404 230444 308456 230450
rect 308404 230386 308456 230392
rect 307944 230036 307996 230042
rect 307944 229978 307996 229984
rect 307668 223304 307720 223310
rect 307668 223246 307720 223252
rect 306840 220244 306892 220250
rect 306840 220186 306892 220192
rect 307392 219020 307444 219026
rect 307392 218962 307444 218968
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306196 218068 306248 218074
rect 306196 218010 306248 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217138 307432 218962
rect 307680 218074 307708 223246
rect 308416 219434 308444 230386
rect 308600 227050 308628 231676
rect 308588 227044 308640 227050
rect 308588 226986 308640 226992
rect 308864 226296 308916 226302
rect 308864 226238 308916 226244
rect 308404 219428 308456 219434
rect 308404 219370 308456 219376
rect 308876 218074 308904 226238
rect 309244 220386 309272 231676
rect 309888 224942 309916 231676
rect 310336 227044 310388 227050
rect 310336 226986 310388 226992
rect 309876 224936 309928 224942
rect 309876 224878 309928 224884
rect 309232 220380 309284 220386
rect 309232 220322 309284 220328
rect 309048 220244 309100 220250
rect 309048 220186 309100 220192
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308220 218068 308272 218074
rect 308220 218010 308272 218016
rect 308864 218068 308916 218074
rect 308864 218010 308916 218016
rect 308232 217138 308260 218010
rect 309060 217274 309088 220186
rect 310348 218074 310376 226986
rect 310532 225486 310560 231676
rect 310520 225480 310572 225486
rect 310520 225422 310572 225428
rect 311176 224670 311204 231676
rect 311360 231662 311834 231690
rect 311164 224664 311216 224670
rect 311164 224606 311216 224612
rect 310704 222148 310756 222154
rect 310704 222090 310756 222096
rect 309876 218068 309928 218074
rect 309876 218010 309928 218016
rect 310336 218068 310388 218074
rect 310336 218010 310388 218016
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217110 307432 217138
rect 308186 217110 308260 217138
rect 309014 217246 309088 217274
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217110
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309888 217138 309916 218010
rect 310716 217274 310744 222090
rect 311360 220522 311388 231662
rect 312464 228410 312492 231676
rect 313108 230314 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230308 313148 230314
rect 313096 230250 313148 230256
rect 312636 230036 312688 230042
rect 312636 229978 312688 229984
rect 312452 228404 312504 228410
rect 312452 228346 312504 228352
rect 311532 224800 311584 224806
rect 311532 224742 311584 224748
rect 311348 220516 311400 220522
rect 311348 220458 311400 220464
rect 311544 217274 311572 224742
rect 312648 222154 312676 229978
rect 312912 225888 312964 225894
rect 312912 225830 312964 225836
rect 312636 222148 312688 222154
rect 312636 222090 312688 222096
rect 312924 218074 312952 225830
rect 313292 225622 313320 231662
rect 313936 229094 313964 231662
rect 313752 229066 313964 229094
rect 313280 225616 313332 225622
rect 313280 225558 313332 225564
rect 313188 222012 313240 222018
rect 313188 221954 313240 221960
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 312912 218068 312964 218074
rect 312912 218010 312964 218016
rect 309842 217110 309916 217138
rect 310670 217246 310744 217274
rect 311498 217246 311572 217274
rect 309842 216988 309870 217110
rect 310670 216988 310698 217246
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313200 217274 313228 221954
rect 313752 221882 313780 229066
rect 313924 228540 313976 228546
rect 313924 228482 313976 228488
rect 313740 221876 313792 221882
rect 313740 221818 313792 221824
rect 313936 219298 313964 228482
rect 315040 223582 315068 231676
rect 315408 231662 315698 231690
rect 315408 229094 315436 231662
rect 315316 229066 315436 229094
rect 315316 224126 315344 229066
rect 315488 227452 315540 227458
rect 315488 227394 315540 227400
rect 315304 224120 315356 224126
rect 315304 224062 315356 224068
rect 315028 223576 315080 223582
rect 315028 223518 315080 223524
rect 313924 219292 313976 219298
rect 313924 219234 313976 219240
rect 314016 218884 314068 218890
rect 314016 218826 314068 218832
rect 312326 217110 312400 217138
rect 313154 217246 313228 217274
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218826
rect 315500 218074 315528 227394
rect 315672 223032 315724 223038
rect 315672 222974 315724 222980
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 315488 218068 315540 218074
rect 315488 218010 315540 218016
rect 314856 217138 314884 218010
rect 315684 217274 315712 222974
rect 316328 222902 316356 231676
rect 316684 223440 316736 223446
rect 316684 223382 316736 223388
rect 316316 222896 316368 222902
rect 316316 222838 316368 222844
rect 316500 220380 316552 220386
rect 316500 220322 316552 220328
rect 316512 217274 316540 220322
rect 316696 218482 316724 223382
rect 316972 222766 317000 231676
rect 317616 227594 317644 231676
rect 318260 229906 318288 231676
rect 318248 229900 318300 229906
rect 318248 229842 318300 229848
rect 318064 229764 318116 229770
rect 318064 229706 318116 229712
rect 317604 227588 317656 227594
rect 317604 227530 317656 227536
rect 316960 222760 317012 222766
rect 316960 222702 317012 222708
rect 318076 219434 318104 229706
rect 318904 228682 318932 231676
rect 319088 231662 319562 231690
rect 320206 231662 320404 231690
rect 318892 228676 318944 228682
rect 318892 228618 318944 228624
rect 318248 221876 318300 221882
rect 318248 221818 318300 221824
rect 318260 219434 318288 221818
rect 319088 219842 319116 231662
rect 320088 228404 320140 228410
rect 320088 228346 320140 228352
rect 319812 224936 319864 224942
rect 319812 224878 319864 224884
rect 319076 219836 319128 219842
rect 319076 219778 319128 219784
rect 317984 219406 318104 219434
rect 318168 219406 318288 219434
rect 316684 218476 316736 218482
rect 316684 218418 316736 218424
rect 317984 218074 318012 219406
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 317972 218068 318024 218074
rect 317972 218010 318024 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217246 315712 217274
rect 316466 217246 316540 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217246
rect 316466 216988 316494 217246
rect 317340 217138 317368 218010
rect 318168 217274 318196 219406
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 317294 217110 317368 217138
rect 318122 217246 318196 217274
rect 317294 216988 317322 217110
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 224878
rect 320100 218074 320128 228346
rect 320376 221474 320404 231662
rect 320836 228546 320864 231676
rect 320824 228540 320876 228546
rect 320824 228482 320876 228488
rect 321480 223174 321508 231676
rect 322124 227730 322152 231676
rect 322112 227724 322164 227730
rect 322112 227666 322164 227672
rect 322112 227588 322164 227594
rect 322112 227530 322164 227536
rect 321468 223168 321520 223174
rect 321468 223110 321520 223116
rect 321468 222896 321520 222902
rect 321468 222838 321520 222844
rect 320364 221468 320416 221474
rect 320364 221410 320416 221416
rect 320640 219428 320692 219434
rect 320640 219370 320692 219376
rect 320088 218068 320140 218074
rect 320088 218010 320140 218016
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219370
rect 321480 217274 321508 222838
rect 322124 219162 322152 227530
rect 322768 226166 322796 231676
rect 323412 229634 323440 231676
rect 323400 229628 323452 229634
rect 323400 229570 323452 229576
rect 322756 226160 322808 226166
rect 322756 226102 322808 226108
rect 322848 224664 322900 224670
rect 322848 224606 322900 224612
rect 322112 219156 322164 219162
rect 322112 219098 322164 219104
rect 322860 218074 322888 224606
rect 324056 224262 324084 231676
rect 324228 229900 324280 229906
rect 324228 229842 324280 229848
rect 324044 224256 324096 224262
rect 324044 224198 324096 224204
rect 323952 223168 324004 223174
rect 323952 223110 324004 223116
rect 323964 218074 323992 223110
rect 324240 219434 324268 229842
rect 324700 219434 324728 231676
rect 325344 227322 325372 231676
rect 325516 228676 325568 228682
rect 325516 228618 325568 228624
rect 325332 227316 325384 227322
rect 325332 227258 325384 227264
rect 324148 219406 324268 219434
rect 324608 219406 324728 219434
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 323124 218068 323176 218074
rect 323124 218010 323176 218016
rect 323952 218068 324004 218074
rect 323952 218010 324004 218016
rect 320606 217110 320680 217138
rect 321434 217246 321508 217274
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217138 323164 218010
rect 324148 217274 324176 219406
rect 324608 218754 324636 219406
rect 325332 219156 325384 219162
rect 325332 219098 325384 219104
rect 324596 218748 324648 218754
rect 324596 218690 324648 218696
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 322262 217110 322336 217138
rect 323090 217110 323164 217138
rect 323918 217246 324176 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217110
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325344 217274 325372 219098
rect 325528 218074 325556 228618
rect 325988 224534 326016 231676
rect 326172 231662 326646 231690
rect 325976 224528 326028 224534
rect 325976 224470 326028 224476
rect 326172 220114 326200 231662
rect 326896 228540 326948 228546
rect 326896 228482 326948 228488
rect 326160 220108 326212 220114
rect 326160 220050 326212 220056
rect 326908 218074 326936 228482
rect 327276 223446 327304 231676
rect 327920 225758 327948 231676
rect 328564 226030 328592 231676
rect 329208 228818 329236 231676
rect 329852 230178 329880 231676
rect 329840 230172 329892 230178
rect 329840 230114 329892 230120
rect 330496 228954 330524 231676
rect 331140 229090 331168 231676
rect 331416 231662 331798 231690
rect 331128 229084 331180 229090
rect 331128 229026 331180 229032
rect 330484 228948 330536 228954
rect 330484 228890 330536 228896
rect 329196 228812 329248 228818
rect 329196 228754 329248 228760
rect 331036 227792 331088 227798
rect 331036 227734 331088 227740
rect 328552 226024 328604 226030
rect 328552 225966 328604 225972
rect 327908 225752 327960 225758
rect 327908 225694 327960 225700
rect 329748 225752 329800 225758
rect 329748 225694 329800 225700
rect 327724 225616 327776 225622
rect 327724 225558 327776 225564
rect 327264 223440 327316 223446
rect 327264 223382 327316 223388
rect 327736 219162 327764 225558
rect 328092 220516 328144 220522
rect 328092 220458 328144 220464
rect 327724 219156 327776 219162
rect 327724 219098 327776 219104
rect 327264 218748 327316 218754
rect 327264 218690 327316 218696
rect 325516 218068 325568 218074
rect 325516 218010 325568 218016
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 325344 217246 325602 217274
rect 324746 217110 324820 217138
rect 324746 216988 324774 217110
rect 325574 216988 325602 217246
rect 326448 217138 326476 218010
rect 327276 217138 327304 218690
rect 328104 217274 328132 220458
rect 328920 220108 328972 220114
rect 328920 220050 328972 220056
rect 328932 217274 328960 220050
rect 329760 217274 329788 225694
rect 331048 218074 331076 227734
rect 331416 224398 331444 231662
rect 332428 227594 332456 231676
rect 332612 231662 333086 231690
rect 333256 231662 333730 231690
rect 334084 231662 334374 231690
rect 332416 227588 332468 227594
rect 332416 227530 332468 227536
rect 331864 224528 331916 224534
rect 331864 224470 331916 224476
rect 331404 224392 331456 224398
rect 331404 224334 331456 224340
rect 331404 222148 331456 222154
rect 331404 222090 331456 222096
rect 330576 218068 330628 218074
rect 330576 218010 330628 218016
rect 331036 218068 331088 218074
rect 331036 218010 331088 218016
rect 326402 217110 326476 217138
rect 327230 217110 327304 217138
rect 328058 217246 328132 217274
rect 328886 217246 328960 217274
rect 329714 217246 329788 217274
rect 326402 216988 326430 217110
rect 327230 216988 327258 217110
rect 328058 216988 328086 217246
rect 328886 216988 328914 217246
rect 329714 216988 329742 217246
rect 330588 217138 330616 218010
rect 331416 217274 331444 222090
rect 331876 219026 331904 224470
rect 332612 221746 332640 231662
rect 332600 221740 332652 221746
rect 332600 221682 332652 221688
rect 332600 221468 332652 221474
rect 332600 221410 332652 221416
rect 332612 219434 332640 221410
rect 333256 220658 333284 231662
rect 333888 227316 333940 227322
rect 333888 227258 333940 227264
rect 333244 220652 333296 220658
rect 333244 220594 333296 220600
rect 332244 219406 332640 219434
rect 331864 219020 331916 219026
rect 331864 218962 331916 218968
rect 332244 217274 332272 219406
rect 333704 219020 333756 219026
rect 333704 218962 333756 218968
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 332198 217246 332272 217274
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332198 216988 332226 217246
rect 333072 217138 333100 218010
rect 333716 217274 333744 218962
rect 333900 218074 333928 227258
rect 334084 221610 334112 231662
rect 335004 230450 335032 231676
rect 334992 230444 335044 230450
rect 334992 230386 335044 230392
rect 334256 230172 334308 230178
rect 334256 230114 334308 230120
rect 334268 227798 334296 230114
rect 334256 227792 334308 227798
rect 334256 227734 334308 227740
rect 335176 226024 335228 226030
rect 335176 225966 335228 225972
rect 334072 221604 334124 221610
rect 334072 221546 334124 221552
rect 335188 218074 335216 225966
rect 335648 223310 335676 231676
rect 336292 226302 336320 231676
rect 336464 228812 336516 228818
rect 336464 228754 336516 228760
rect 336280 226296 336332 226302
rect 336280 226238 336332 226244
rect 335636 223304 335688 223310
rect 335636 223246 335688 223252
rect 336476 219434 336504 228754
rect 336936 227186 336964 231676
rect 336924 227180 336976 227186
rect 336924 227122 336976 227128
rect 337580 224534 337608 231676
rect 337752 227588 337804 227594
rect 337752 227530 337804 227536
rect 337568 224528 337620 224534
rect 337568 224470 337620 224476
rect 336384 219406 336504 219434
rect 335544 218204 335596 218210
rect 335544 218146 335596 218152
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335176 218068 335228 218074
rect 335176 218010 335228 218016
rect 333716 217246 333882 217274
rect 333026 217110 333100 217138
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218146
rect 336384 217274 336412 219406
rect 337764 218074 337792 227530
rect 338224 227050 338252 231676
rect 338212 227044 338264 227050
rect 338212 226986 338264 226992
rect 338672 227044 338724 227050
rect 338672 226986 338724 226992
rect 337936 223304 337988 223310
rect 337936 223246 337988 223252
rect 337200 218068 337252 218074
rect 337200 218010 337252 218016
rect 337752 218068 337804 218074
rect 337752 218010 337804 218016
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336412 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218010
rect 337948 217274 337976 223246
rect 338684 218210 338712 226986
rect 338868 224806 338896 231676
rect 339526 231662 339724 231690
rect 338856 224800 338908 224806
rect 338856 224742 338908 224748
rect 339408 224256 339460 224262
rect 339408 224198 339460 224204
rect 338672 218204 338724 218210
rect 338672 218146 338724 218152
rect 339420 218074 339448 224198
rect 339696 220250 339724 231662
rect 340156 230042 340184 231676
rect 340432 231662 340814 231690
rect 340144 230036 340196 230042
rect 340144 229978 340196 229984
rect 340432 222018 340460 231662
rect 341444 227458 341472 231676
rect 341720 231662 342102 231690
rect 342364 231662 342746 231690
rect 342916 231662 343390 231690
rect 343836 231662 344034 231690
rect 341432 227452 341484 227458
rect 341432 227394 341484 227400
rect 340696 227180 340748 227186
rect 340696 227122 340748 227128
rect 340420 222012 340472 222018
rect 340420 221954 340472 221960
rect 340052 220788 340104 220794
rect 340052 220730 340104 220736
rect 339684 220244 339736 220250
rect 339684 220186 339736 220192
rect 340064 218890 340092 220730
rect 340512 219156 340564 219162
rect 340512 219098 340564 219104
rect 340052 218884 340104 218890
rect 340052 218826 340104 218832
rect 338856 218068 338908 218074
rect 338856 218010 338908 218016
rect 339408 218068 339460 218074
rect 339408 218010 339460 218016
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337948 217246 338022 217274
rect 337166 217110 337240 217138
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338868 217138 338896 218010
rect 339696 217138 339724 218010
rect 340524 217138 340552 219098
rect 340708 218074 340736 227122
rect 341720 225894 341748 231662
rect 341708 225888 341760 225894
rect 341708 225830 341760 225836
rect 341984 225888 342036 225894
rect 341984 225830 342036 225836
rect 341996 219434 342024 225830
rect 342168 224392 342220 224398
rect 342168 224334 342220 224340
rect 342180 219434 342208 224334
rect 342364 220794 342392 231662
rect 342352 220788 342404 220794
rect 342352 220730 342404 220736
rect 342916 220386 342944 231662
rect 343836 221882 343864 231662
rect 344664 223038 344692 231676
rect 345020 229764 345072 229770
rect 345020 229706 345072 229712
rect 345032 227594 345060 229706
rect 345308 229634 345336 231676
rect 345296 229628 345348 229634
rect 345296 229570 345348 229576
rect 345020 227588 345072 227594
rect 345020 227530 345072 227536
rect 345952 224942 345980 231676
rect 345940 224936 345992 224942
rect 345940 224878 345992 224884
rect 346308 224528 346360 224534
rect 346308 224470 346360 224476
rect 344652 223032 344704 223038
rect 344652 222974 344704 222980
rect 345296 222896 345348 222902
rect 345296 222838 345348 222844
rect 343824 221876 343876 221882
rect 343824 221818 343876 221824
rect 344652 221740 344704 221746
rect 344652 221682 344704 221688
rect 342904 220380 342956 220386
rect 342904 220322 342956 220328
rect 342996 220244 343048 220250
rect 342996 220186 343048 220192
rect 341340 219428 341392 219434
rect 341996 219406 342116 219434
rect 342180 219428 342312 219434
rect 342180 219406 342260 219428
rect 341340 219370 341392 219376
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217138 341380 219370
rect 342088 217274 342116 219406
rect 342260 219370 342312 219376
rect 343008 217274 343036 220186
rect 343824 219428 343876 219434
rect 343824 219370 343876 219376
rect 342088 217246 342162 217274
rect 338822 217110 338896 217138
rect 339650 217110 339724 217138
rect 340478 217110 340552 217138
rect 341306 217110 341380 217138
rect 338822 216988 338850 217110
rect 339650 216988 339678 217110
rect 340478 216988 340506 217110
rect 341306 216988 341334 217110
rect 342134 216988 342162 217246
rect 342962 217246 343036 217274
rect 342962 216988 342990 217246
rect 343836 217138 343864 219370
rect 344664 217274 344692 221682
rect 345308 219298 345336 222838
rect 345296 219292 345348 219298
rect 345296 219234 345348 219240
rect 345480 218068 345532 218074
rect 345480 218010 345532 218016
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345492 217138 345520 218010
rect 346320 217274 346348 224470
rect 346596 223038 346624 231676
rect 346872 231662 347254 231690
rect 346872 228410 346900 231662
rect 346860 228404 346912 228410
rect 346860 228346 346912 228352
rect 347044 228404 347096 228410
rect 347044 228346 347096 228352
rect 346584 223032 346636 223038
rect 346584 222974 346636 222980
rect 347056 219434 347084 228346
rect 347884 222902 347912 231676
rect 348528 223174 348556 231676
rect 349172 228682 349200 231676
rect 349160 228676 349212 228682
rect 349160 228618 349212 228624
rect 349816 224670 349844 231676
rect 350460 229906 350488 231676
rect 350448 229900 350500 229906
rect 350448 229842 350500 229848
rect 350172 228676 350224 228682
rect 350172 228618 350224 228624
rect 349804 224664 349856 224670
rect 349804 224606 349856 224612
rect 348516 223168 348568 223174
rect 348516 223110 348568 223116
rect 349068 223032 349120 223038
rect 349068 222974 349120 222980
rect 347872 222896 347924 222902
rect 347872 222838 347924 222844
rect 347228 222760 347280 222766
rect 347228 222702 347280 222708
rect 347044 219428 347096 219434
rect 347044 219370 347096 219376
rect 347044 218884 347096 218890
rect 347044 218826 347096 218832
rect 345446 217110 345520 217138
rect 346274 217246 346348 217274
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347056 217138 347084 218826
rect 347240 218074 347268 222702
rect 348792 221604 348844 221610
rect 348792 221546 348844 221552
rect 347228 218068 347280 218074
rect 347228 218010 347280 218016
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 347976 217138 348004 218010
rect 348804 217274 348832 221546
rect 349080 218074 349108 222974
rect 350184 218074 350212 228618
rect 351104 228546 351132 231676
rect 351288 231662 351762 231690
rect 351092 228540 351144 228546
rect 351092 228482 351144 228488
rect 351092 227792 351144 227798
rect 351092 227734 351144 227740
rect 350356 224732 350408 224738
rect 350356 224674 350408 224680
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 349620 218068 349672 218074
rect 349620 218010 349672 218016
rect 350172 218068 350224 218074
rect 350172 218010 350224 218016
rect 347056 217110 347130 217138
rect 347102 216988 347130 217110
rect 347930 217110 348004 217138
rect 348758 217246 348832 217274
rect 347930 216988 347958 217110
rect 348758 216988 348786 217246
rect 349632 217138 349660 218010
rect 350368 217274 350396 224674
rect 351104 218754 351132 227734
rect 351288 220522 351316 231662
rect 352392 225622 352420 231676
rect 353036 227798 353064 231676
rect 353024 227792 353076 227798
rect 353024 227734 353076 227740
rect 352564 227452 352616 227458
rect 352564 227394 352616 227400
rect 352380 225616 352432 225622
rect 352380 225558 352432 225564
rect 351276 220516 351328 220522
rect 351276 220458 351328 220464
rect 351276 220380 351328 220386
rect 351276 220322 351328 220328
rect 351092 218748 351144 218754
rect 351092 218690 351144 218696
rect 351288 217274 351316 220322
rect 352576 219162 352604 227394
rect 353680 225758 353708 231676
rect 353956 231662 354338 231690
rect 354784 231662 354982 231690
rect 353668 225752 353720 225758
rect 353668 225694 353720 225700
rect 352932 225616 352984 225622
rect 352932 225558 352984 225564
rect 352564 219156 352616 219162
rect 352564 219098 352616 219104
rect 352104 218068 352156 218074
rect 352104 218010 352156 218016
rect 350368 217246 350442 217274
rect 349586 217110 349660 217138
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351316 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 218010
rect 352944 217274 352972 225558
rect 353956 222154 353984 231662
rect 354588 228540 354640 228546
rect 354588 228482 354640 228488
rect 353944 222148 353996 222154
rect 353944 222090 353996 222096
rect 353300 221876 353352 221882
rect 353300 221818 353352 221824
rect 353312 218074 353340 221818
rect 353760 218748 353812 218754
rect 353760 218690 353812 218696
rect 353300 218068 353352 218074
rect 353300 218010 353352 218016
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218690
rect 354600 217274 354628 228482
rect 354784 220114 354812 231662
rect 355612 230178 355640 231676
rect 355600 230172 355652 230178
rect 355600 230114 355652 230120
rect 354956 230036 355008 230042
rect 354956 229978 355008 229984
rect 354968 224738 354996 229978
rect 356256 227322 356284 231676
rect 356244 227316 356296 227322
rect 356244 227258 356296 227264
rect 356900 226030 356928 231676
rect 357256 227316 357308 227322
rect 357256 227258 357308 227264
rect 356888 226024 356940 226030
rect 356888 225966 356940 225972
rect 355232 225004 355284 225010
rect 355232 224946 355284 224952
rect 354956 224732 355008 224738
rect 354956 224674 355008 224680
rect 354772 220108 354824 220114
rect 354772 220050 354824 220056
rect 355244 219026 355272 224946
rect 355416 220108 355468 220114
rect 355416 220050 355468 220056
rect 355232 219020 355284 219026
rect 355232 218962 355284 218968
rect 355428 217274 355456 220050
rect 357072 219020 357124 219026
rect 357072 218962 357124 218968
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 353726 217110 353800 217138
rect 354554 217246 354628 217274
rect 355382 217246 355456 217274
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355382 216988 355410 217246
rect 356256 217138 356284 218010
rect 357084 217138 357112 218962
rect 357268 218074 357296 227258
rect 357544 221474 357572 231676
rect 358188 225010 358216 231676
rect 358832 228818 358860 231676
rect 359200 231662 359490 231690
rect 358820 228812 358872 228818
rect 358820 228754 358872 228760
rect 358176 225004 358228 225010
rect 358176 224946 358228 224952
rect 359200 223310 359228 231662
rect 359924 228812 359976 228818
rect 359924 228754 359976 228760
rect 359464 224664 359516 224670
rect 359464 224606 359516 224612
rect 359188 223304 359240 223310
rect 359188 223246 359240 223252
rect 358544 223168 358596 223174
rect 358544 223110 358596 223116
rect 357532 221468 357584 221474
rect 357532 221410 357584 221416
rect 358556 218074 358584 223110
rect 359476 218210 359504 224606
rect 359936 219434 359964 228754
rect 360120 227050 360148 231676
rect 360764 229770 360792 231676
rect 360752 229764 360804 229770
rect 360752 229706 360804 229712
rect 361212 229764 361264 229770
rect 361212 229706 361264 229712
rect 361224 229094 361252 229706
rect 361040 229066 361252 229094
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359936 219406 360148 219434
rect 358728 218204 358780 218210
rect 358728 218146 358780 218152
rect 359464 218204 359516 218210
rect 359464 218146 359516 218152
rect 357256 218068 357308 218074
rect 357256 218010 357308 218016
rect 357900 218068 357952 218074
rect 357900 218010 357952 218016
rect 358544 218068 358596 218074
rect 358544 218010 358596 218016
rect 357912 217138 357940 218010
rect 358740 217138 358768 218146
rect 360120 218074 360148 219406
rect 361040 218074 361068 229066
rect 361408 227186 361436 231676
rect 361396 227180 361448 227186
rect 361396 227122 361448 227128
rect 361212 226024 361264 226030
rect 361212 225966 361264 225972
rect 359556 218068 359608 218074
rect 359556 218010 359608 218016
rect 360108 218068 360160 218074
rect 360108 218010 360160 218016
rect 360384 218068 360436 218074
rect 360384 218010 360436 218016
rect 361028 218068 361080 218074
rect 361028 218010 361080 218016
rect 359568 217138 359596 218010
rect 360396 217138 360424 218010
rect 361224 217274 361252 225966
rect 362052 224398 362080 231676
rect 362328 231662 362710 231690
rect 362040 224392 362092 224398
rect 362040 224334 362092 224340
rect 362328 224262 362356 231662
rect 363340 227458 363368 231676
rect 363524 231662 363998 231690
rect 364536 231662 364642 231690
rect 363328 227452 363380 227458
rect 363328 227394 363380 227400
rect 363524 227338 363552 231662
rect 363340 227310 363552 227338
rect 362776 227044 362828 227050
rect 362776 226986 362828 226992
rect 362316 224256 362368 224262
rect 362316 224198 362368 224204
rect 362040 219156 362092 219162
rect 362040 219098 362092 219104
rect 362052 217274 362080 219098
rect 356210 217110 356284 217138
rect 357038 217110 357112 217138
rect 357866 217110 357940 217138
rect 358694 217110 358768 217138
rect 359522 217110 359596 217138
rect 360350 217110 360424 217138
rect 361178 217246 361252 217274
rect 362006 217246 362080 217274
rect 362788 217274 362816 226986
rect 363340 220250 363368 227310
rect 363512 227180 363564 227186
rect 363512 227122 363564 227128
rect 363328 220244 363380 220250
rect 363328 220186 363380 220192
rect 363524 218890 363552 227122
rect 364536 221746 364564 231662
rect 365272 225894 365300 231676
rect 365916 228410 365944 231676
rect 365904 228404 365956 228410
rect 365904 228346 365956 228352
rect 365260 225888 365312 225894
rect 365260 225830 365312 225836
rect 365352 225752 365404 225758
rect 365352 225694 365404 225700
rect 364524 221740 364576 221746
rect 364524 221682 364576 221688
rect 364524 220516 364576 220522
rect 364524 220458 364576 220464
rect 363696 220244 363748 220250
rect 363696 220186 363748 220192
rect 363512 218884 363564 218890
rect 363512 218826 363564 218832
rect 363708 217274 363736 220186
rect 364536 217274 364564 220458
rect 365364 217274 365392 225694
rect 366560 224534 366588 231676
rect 366732 229900 366784 229906
rect 366732 229842 366784 229848
rect 366744 229094 366772 229842
rect 366744 229066 366956 229094
rect 366548 224528 366600 224534
rect 366548 224470 366600 224476
rect 366732 224392 366784 224398
rect 366732 224334 366784 224340
rect 366744 219570 366772 224334
rect 366732 219564 366784 219570
rect 366732 219506 366784 219512
rect 366180 219428 366232 219434
rect 366180 219370 366232 219376
rect 362788 217246 362862 217274
rect 356210 216988 356238 217110
rect 357038 216988 357066 217110
rect 357866 216988 357894 217110
rect 358694 216988 358722 217110
rect 359522 216988 359550 217110
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 362006 216988 362034 217246
rect 362834 216988 362862 217246
rect 363662 217246 363736 217274
rect 364490 217246 364564 217274
rect 365318 217246 365392 217274
rect 363662 216988 363690 217246
rect 364490 216988 364518 217246
rect 365318 216988 365346 217246
rect 366192 217138 366220 219370
rect 366928 217274 366956 229066
rect 367204 223038 367232 231676
rect 367192 223032 367244 223038
rect 367192 222974 367244 222980
rect 367848 222902 367876 231676
rect 368492 227186 368520 231676
rect 369136 228682 369164 231676
rect 369320 231662 369794 231690
rect 370056 231662 370438 231690
rect 369124 228676 369176 228682
rect 369124 228618 369176 228624
rect 368480 227180 368532 227186
rect 368480 227122 368532 227128
rect 369124 226500 369176 226506
rect 369124 226442 369176 226448
rect 368388 223032 368440 223038
rect 368388 222974 368440 222980
rect 367836 222896 367888 222902
rect 367836 222838 367888 222844
rect 368400 218074 368428 222974
rect 369136 219026 369164 226442
rect 369320 220386 369348 231662
rect 370056 221610 370084 231662
rect 371068 230042 371096 231676
rect 371056 230036 371108 230042
rect 371056 229978 371108 229984
rect 371712 229094 371740 231676
rect 371620 229066 371740 229094
rect 371148 228404 371200 228410
rect 371148 228346 371200 228352
rect 370964 221740 371016 221746
rect 370964 221682 371016 221688
rect 370044 221604 370096 221610
rect 370044 221546 370096 221552
rect 369492 221468 369544 221474
rect 369492 221410 369544 221416
rect 369308 220380 369360 220386
rect 369308 220322 369360 220328
rect 369124 219020 369176 219026
rect 369124 218962 369176 218968
rect 368664 218884 368716 218890
rect 368664 218826 368716 218832
rect 367836 218068 367888 218074
rect 367836 218010 367888 218016
rect 368388 218068 368440 218074
rect 368388 218010 368440 218016
rect 366928 217246 367002 217274
rect 366146 217110 366220 217138
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367848 217138 367876 218010
rect 368676 217138 368704 218826
rect 369504 217274 369532 221410
rect 370976 219162 371004 221682
rect 370964 219156 371016 219162
rect 370964 219098 371016 219104
rect 370320 219020 370372 219026
rect 370320 218962 370372 218968
rect 367802 217110 367876 217138
rect 368630 217110 368704 217138
rect 369458 217246 369532 217274
rect 367802 216988 367830 217110
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370332 217138 370360 218962
rect 371160 217274 371188 228346
rect 371620 225622 371648 229066
rect 372356 228546 372384 231676
rect 372724 231662 373014 231690
rect 372344 228540 372396 228546
rect 372344 228482 372396 228488
rect 371792 227792 371844 227798
rect 371792 227734 371844 227740
rect 371608 225616 371660 225622
rect 371608 225558 371660 225564
rect 371804 218754 371832 227734
rect 372528 224256 372580 224262
rect 372528 224198 372580 224204
rect 371792 218748 371844 218754
rect 371792 218690 371844 218696
rect 372540 218074 372568 224198
rect 372724 221882 372752 231662
rect 373448 228540 373500 228546
rect 373448 228482 373500 228488
rect 372712 221876 372764 221882
rect 372712 221818 372764 221824
rect 373460 219434 373488 228482
rect 373644 227798 373672 231676
rect 373632 227792 373684 227798
rect 373632 227734 373684 227740
rect 374288 227322 374316 231676
rect 374656 231662 374946 231690
rect 374276 227316 374328 227322
rect 374276 227258 374328 227264
rect 374656 223174 374684 231662
rect 375012 225888 375064 225894
rect 375012 225830 375064 225836
rect 374644 223168 374696 223174
rect 374644 223110 374696 223116
rect 373724 221604 373776 221610
rect 373724 221546 373776 221552
rect 373460 219406 373580 219434
rect 373552 218074 373580 219406
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 373540 218068 373592 218074
rect 373540 218010 373592 218016
rect 370286 217110 370360 217138
rect 371114 217246 371188 217274
rect 370286 216988 370314 217110
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373736 217274 373764 221546
rect 375024 218074 375052 225830
rect 375196 222896 375248 222902
rect 375196 222838 375248 222844
rect 374460 218068 374512 218074
rect 374460 218010 374512 218016
rect 375012 218068 375064 218074
rect 375012 218010 375064 218016
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217246 373764 217274
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217246
rect 374472 217138 374500 218010
rect 375208 217274 375236 222838
rect 375576 220114 375604 231676
rect 376220 226506 376248 231676
rect 376864 228818 376892 231676
rect 376852 228812 376904 228818
rect 376852 228754 376904 228760
rect 376668 227180 376720 227186
rect 376668 227122 376720 227128
rect 376208 226500 376260 226506
rect 376208 226442 376260 226448
rect 375564 220108 375616 220114
rect 375564 220050 375616 220056
rect 376680 218074 376708 227122
rect 377508 226030 377536 231676
rect 377772 228676 377824 228682
rect 377772 228618 377824 228624
rect 377496 226024 377548 226030
rect 377496 225966 377548 225972
rect 376944 220380 376996 220386
rect 376944 220322 376996 220328
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376668 218068 376720 218074
rect 376668 218010 376720 218016
rect 375208 217246 375282 217274
rect 374426 217110 374500 217138
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217274 376984 220322
rect 377784 217274 377812 228618
rect 378152 224670 378180 231676
rect 378796 229770 378824 231676
rect 379072 231662 379454 231690
rect 379716 231662 380098 231690
rect 380360 231662 380742 231690
rect 381096 231662 381386 231690
rect 381648 231662 382030 231690
rect 378784 229764 378836 229770
rect 378784 229706 378836 229712
rect 379072 227050 379100 231662
rect 379060 227044 379112 227050
rect 379060 226986 379112 226992
rect 378784 226840 378836 226846
rect 378784 226782 378836 226788
rect 378140 224664 378192 224670
rect 378140 224606 378192 224612
rect 378796 218890 378824 226782
rect 379244 224528 379296 224534
rect 379244 224470 379296 224476
rect 378784 218884 378836 218890
rect 378784 218826 378836 218832
rect 379256 218074 379284 224470
rect 379716 220522 379744 231662
rect 380360 221882 380388 231662
rect 380348 221876 380400 221882
rect 380348 221818 380400 221824
rect 380072 221740 380124 221746
rect 380072 221682 380124 221688
rect 379704 220516 379756 220522
rect 379704 220458 379756 220464
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 379244 218068 379296 218074
rect 379244 218010 379296 218016
rect 376082 217110 376156 217138
rect 376910 217246 376984 217274
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217246
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379440 217274 379468 220050
rect 380084 219026 380112 221682
rect 381096 220250 381124 231662
rect 381648 224398 381676 231662
rect 382096 227316 382148 227322
rect 382096 227258 382148 227264
rect 381636 224392 381688 224398
rect 381636 224334 381688 224340
rect 381084 220244 381136 220250
rect 381084 220186 381136 220192
rect 380072 219020 380124 219026
rect 380072 218962 380124 218968
rect 380256 219020 380308 219026
rect 380256 218962 380308 218968
rect 378566 217110 378640 217138
rect 379394 217246 379468 217274
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 218962
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381096 217138 381124 218010
rect 381924 217138 381952 218146
rect 382108 218074 382136 227258
rect 382660 223038 382688 231676
rect 383304 225758 383332 231676
rect 383948 229906 383976 231676
rect 384132 231662 384606 231690
rect 383936 229900 383988 229906
rect 383936 229842 383988 229848
rect 383292 225752 383344 225758
rect 383292 225694 383344 225700
rect 382924 225616 382976 225622
rect 382924 225558 382976 225564
rect 382648 223032 382700 223038
rect 382648 222974 382700 222980
rect 382740 218884 382792 218890
rect 382740 218826 382792 218832
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217138 382780 218826
rect 382936 218210 382964 225558
rect 383568 223032 383620 223038
rect 383568 222974 383620 222980
rect 383580 218890 383608 222974
rect 384132 221474 384160 231662
rect 384304 229560 384356 229566
rect 384304 229502 384356 229508
rect 384316 221610 384344 229502
rect 385236 228410 385264 231676
rect 385224 228404 385276 228410
rect 385224 228346 385276 228352
rect 385880 226846 385908 231676
rect 386236 228404 386288 228410
rect 386236 228346 386288 228352
rect 385868 226840 385920 226846
rect 385868 226782 385920 226788
rect 386052 226432 386104 226438
rect 386052 226374 386104 226380
rect 384304 221604 384356 221610
rect 384304 221546 384356 221552
rect 384120 221468 384172 221474
rect 384120 221410 384172 221416
rect 384396 221468 384448 221474
rect 384396 221410 384448 221416
rect 383568 218884 383620 218890
rect 383568 218826 383620 218832
rect 383568 218748 383620 218754
rect 383568 218690 383620 218696
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 383580 217138 383608 218690
rect 384408 217274 384436 221410
rect 386064 218074 386092 226374
rect 385224 218068 385276 218074
rect 385224 218010 385276 218016
rect 386052 218068 386104 218074
rect 386052 218010 386104 218016
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217110 381952 217138
rect 382706 217110 382780 217138
rect 383534 217110 383608 217138
rect 384362 217246 384436 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217110
rect 382706 216988 382734 217110
rect 383534 216988 383562 217110
rect 384362 216988 384390 217246
rect 385236 217138 385264 218010
rect 386248 217274 386276 228346
rect 386524 221746 386552 231676
rect 387168 228546 387196 231676
rect 387432 230376 387484 230382
rect 387432 230318 387484 230324
rect 387156 228540 387208 228546
rect 387156 228482 387208 228488
rect 387444 224262 387472 230318
rect 387812 225894 387840 231676
rect 388456 230382 388484 231676
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 388444 230240 388496 230246
rect 388444 230182 388496 230188
rect 387800 225888 387852 225894
rect 387800 225830 387852 225836
rect 387708 225752 387760 225758
rect 387708 225694 387760 225700
rect 387432 224256 387484 224262
rect 387432 224198 387484 224204
rect 386512 221740 386564 221746
rect 386512 221682 386564 221688
rect 386880 218884 386932 218890
rect 386880 218826 386932 218832
rect 385190 217110 385264 217138
rect 386018 217246 386276 217274
rect 385190 216988 385218 217110
rect 386018 216988 386046 217246
rect 386892 217138 386920 218826
rect 387720 217274 387748 225694
rect 388456 220386 388484 230182
rect 389100 229566 389128 231676
rect 389088 229560 389140 229566
rect 389088 229502 389140 229508
rect 389744 227186 389772 231676
rect 390388 228682 390416 231676
rect 390376 228676 390428 228682
rect 390376 228618 390428 228624
rect 390468 228540 390520 228546
rect 390468 228482 390520 228488
rect 389732 227180 389784 227186
rect 389732 227122 389784 227128
rect 388628 226296 388680 226302
rect 388628 226238 388680 226244
rect 388444 220380 388496 220386
rect 388444 220322 388496 220328
rect 388444 220244 388496 220250
rect 388444 220186 388496 220192
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 388456 217274 388484 220186
rect 388640 219026 388668 226238
rect 390192 224256 390244 224262
rect 390192 224198 390244 224204
rect 388628 219020 388680 219026
rect 388628 218962 388680 218968
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 388456 217246 388530 217274
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388502 216988 388530 217246
rect 389376 217138 389404 218010
rect 390204 217274 390232 224198
rect 390480 218074 390508 228482
rect 391032 222902 391060 231676
rect 391676 230246 391704 231676
rect 392136 231662 392334 231690
rect 391664 230240 391716 230246
rect 391664 230182 391716 230188
rect 391204 229764 391256 229770
rect 391204 229706 391256 229712
rect 391216 226438 391244 229706
rect 391756 227044 391808 227050
rect 391756 226986 391808 226992
rect 391204 226432 391256 226438
rect 391204 226374 391256 226380
rect 391020 222896 391072 222902
rect 391020 222838 391072 222844
rect 391020 221604 391072 221610
rect 391020 221546 391072 221552
rect 390468 218068 390520 218074
rect 390468 218010 390520 218016
rect 391032 217274 391060 221546
rect 389330 217110 389404 217138
rect 390158 217246 390232 217274
rect 390986 217246 391060 217274
rect 391768 217274 391796 226986
rect 392136 220114 392164 231662
rect 392964 227322 392992 231676
rect 392952 227316 393004 227322
rect 392952 227258 393004 227264
rect 393136 227180 393188 227186
rect 393136 227122 393188 227128
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 393148 218074 393176 227122
rect 393608 224534 393636 231676
rect 394252 226302 394280 231676
rect 394240 226296 394292 226302
rect 394240 226238 394292 226244
rect 394332 225888 394384 225894
rect 394332 225830 394384 225836
rect 393596 224528 393648 224534
rect 393596 224470 393648 224476
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393136 218068 393188 218074
rect 393136 218010 393188 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 391768 217246 391842 217274
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217274 394372 225830
rect 394516 224392 394568 224398
rect 394516 224334 394568 224340
rect 394528 218074 394556 224334
rect 394896 223038 394924 231676
rect 395172 231662 395554 231690
rect 394884 223032 394936 223038
rect 394884 222974 394936 222980
rect 395172 221474 395200 231662
rect 396184 225622 396212 231676
rect 396368 231662 396842 231690
rect 396172 225616 396224 225622
rect 396172 225558 396224 225564
rect 395804 222896 395856 222902
rect 395804 222838 395856 222844
rect 395160 221468 395212 221474
rect 395160 221410 395212 221416
rect 395816 218074 395844 222838
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395804 218068 395856 218074
rect 395804 218010 395856 218016
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217246 394372 217274
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217246
rect 395172 217138 395200 218010
rect 396000 217274 396028 220050
rect 396368 219434 396396 231662
rect 397472 228410 397500 231676
rect 397840 231662 398130 231690
rect 397460 228404 397512 228410
rect 397460 228346 397512 228352
rect 397840 225758 397868 231662
rect 398104 230376 398156 230382
rect 398104 230318 398156 230324
rect 397828 225752 397880 225758
rect 397828 225694 397880 225700
rect 396816 221468 396868 221474
rect 396816 221410 396868 221416
rect 396276 219406 396396 219434
rect 396276 218754 396304 219406
rect 396264 218748 396316 218754
rect 396264 218690 396316 218696
rect 396828 217274 396856 221410
rect 398116 218890 398144 230318
rect 398760 229770 398788 231676
rect 399404 230382 399432 231676
rect 399392 230376 399444 230382
rect 399392 230318 399444 230324
rect 398748 229764 398800 229770
rect 398748 229706 398800 229712
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 399864 219434 399892 229706
rect 400048 228546 400076 231676
rect 400416 231662 400706 231690
rect 400968 231662 401350 231690
rect 400036 228540 400088 228546
rect 400036 228482 400088 228488
rect 400128 228132 400180 228138
rect 400128 228074 400180 228080
rect 400140 219434 400168 228074
rect 400416 221610 400444 231662
rect 400404 221604 400456 221610
rect 400404 221546 400456 221552
rect 400968 220250 400996 231662
rect 401980 224262 402008 231676
rect 402624 227322 402652 231676
rect 402796 228404 402848 228410
rect 402796 228346 402848 228352
rect 402612 227316 402664 227322
rect 402612 227258 402664 227264
rect 402244 227180 402296 227186
rect 402244 227122 402296 227128
rect 401968 224256 402020 224262
rect 401968 224198 402020 224204
rect 401324 221604 401376 221610
rect 401324 221546 401376 221552
rect 400956 220244 401008 220250
rect 400956 220186 401008 220192
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 398104 218884 398156 218890
rect 398104 218826 398156 218832
rect 398472 218612 398524 218618
rect 398472 218554 398524 218560
rect 397644 218068 397696 218074
rect 397644 218010 397696 218016
rect 397656 217274 397684 218010
rect 395126 217110 395200 217138
rect 395954 217246 396028 217274
rect 396782 217246 396856 217274
rect 397610 217246 397684 217274
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397610 216988 397638 217246
rect 398484 217138 398512 218554
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 400956 218204 401008 218210
rect 400956 218146 401008 218152
rect 400048 217246 400122 217274
rect 398438 217110 398512 217138
rect 399266 217110 399340 217138
rect 398438 216988 398466 217110
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218146
rect 401336 218074 401364 221546
rect 402256 218210 402284 227122
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 401324 218068 401376 218074
rect 401324 218010 401376 218016
rect 401784 218068 401836 218074
rect 401784 218010 401836 218016
rect 401796 217138 401824 218010
rect 402624 217138 402652 218826
rect 402808 218074 402836 228346
rect 403268 225894 403296 231676
rect 403544 231662 403926 231690
rect 403544 227050 403572 231662
rect 403532 227044 403584 227050
rect 403532 226986 403584 226992
rect 403992 226500 404044 226506
rect 403992 226442 404044 226448
rect 403256 225888 403308 225894
rect 403256 225830 403308 225836
rect 404004 218074 404032 226442
rect 404176 225004 404228 225010
rect 404176 224946 404228 224952
rect 402796 218068 402848 218074
rect 402796 218010 402848 218016
rect 403440 218068 403492 218074
rect 403440 218010 403492 218016
rect 403992 218068 404044 218074
rect 403992 218010 404044 218016
rect 403452 217138 403480 218010
rect 404188 217274 404216 224946
rect 404556 224398 404584 231676
rect 404740 231662 405214 231690
rect 404544 224392 404596 224398
rect 404544 224334 404596 224340
rect 404740 220114 404768 231662
rect 405556 224256 405608 224262
rect 405556 224198 405608 224204
rect 404728 220108 404780 220114
rect 404728 220050 404780 220056
rect 405568 218074 405596 224198
rect 405844 221610 405872 231676
rect 406488 222902 406516 231676
rect 407146 231662 407344 231690
rect 406752 223576 406804 223582
rect 406752 223518 406804 223524
rect 406476 222896 406528 222902
rect 406476 222838 406528 222844
rect 405832 221604 405884 221610
rect 405832 221546 405884 221552
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405096 218068 405148 218074
rect 405096 218010 405148 218016
rect 405556 218068 405608 218074
rect 405556 218010 405608 218016
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405108 217138 405136 218010
rect 405936 217274 405964 219438
rect 406764 217274 406792 223518
rect 407316 221474 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 408696 231662 409078 231690
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 408696 226370 408724 231662
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228540 409840 228546
rect 409788 228482 409840 228488
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 408684 226364 408736 226370
rect 408684 226306 408736 226312
rect 407304 221468 407356 221474
rect 407304 221410 407356 221416
rect 407776 218618 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218612 407816 218618
rect 407764 218554 407816 218560
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 405062 217110 405136 217138
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217110
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 221410
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228482
rect 410352 227798 410380 231676
rect 410720 231662 411010 231690
rect 410720 229094 410748 231662
rect 410892 229764 410944 229770
rect 410892 229706 410944 229712
rect 410904 229094 410932 229706
rect 410628 229066 410748 229094
rect 410812 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410628 225010 410656 229066
rect 410616 225004 410668 225010
rect 410616 224946 410668 224952
rect 410812 219434 410840 229066
rect 411640 228410 411668 231676
rect 411628 228404 411680 228410
rect 411628 228346 411680 228352
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 410984 225616 411036 225622
rect 410984 225558 411036 225564
rect 410996 219434 411024 225558
rect 410720 219406 410840 219434
rect 410904 219406 411024 219434
rect 410720 218074 410748 219406
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 219406
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412284 226506 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 226500 412324 226506
rect 412272 226442 412324 226448
rect 412560 218890 412588 226986
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229356 413888 229362
rect 413836 229298 413888 229304
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229298
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223582 414888 231676
rect 415504 228546 415532 231676
rect 415492 228540 415544 228546
rect 415492 228482 415544 228488
rect 415032 228064 415084 228070
rect 415032 228006 415084 228012
rect 414848 223576 414900 223582
rect 414848 223518 414900 223524
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 228006
rect 416148 225622 416176 231676
rect 416792 229094 416820 231676
rect 417436 229770 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229764 417476 229770
rect 417424 229706 417476 229712
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416688 227928 416740 227934
rect 416688 227870 416740 227876
rect 416136 225616 416188 225622
rect 416136 225558 416188 225564
rect 416504 225004 416556 225010
rect 416504 224946 416556 224952
rect 416516 219434 416544 224946
rect 416700 219434 416728 227870
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418356 224954 418384 231662
rect 419368 227050 419396 231676
rect 420012 229362 420040 231676
rect 420000 229356 420052 229362
rect 420000 229298 420052 229304
rect 420656 227934 420684 231676
rect 421024 231662 421314 231690
rect 420644 227928 420696 227934
rect 420644 227870 420696 227876
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 418172 224926 418384 224954
rect 418172 220794 418200 224926
rect 418344 220856 418396 220862
rect 418344 220798 418396 220804
rect 418160 220788 418212 220794
rect 418160 220730 418212 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 418356 217274 418384 220798
rect 420656 219434 420684 227734
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420656 219406 420776 219434
rect 419172 219292 419224 219298
rect 419172 219234 419224 219240
rect 419184 217274 419212 219234
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 417482 217110 417556 217138
rect 418310 217246 418384 217274
rect 419138 217246 419212 217274
rect 417482 216988 417510 217110
rect 418310 216988 418338 217246
rect 419138 216988 419166 217246
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 228070 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 421932 228064 421984 228070
rect 421932 228006 421984 228012
rect 422220 225010 422248 229066
rect 422208 225004 422260 225010
rect 422208 224946 422260 224952
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 423508 219434 423536 229094
rect 423876 227798 423904 231676
rect 424060 231662 424534 231690
rect 423864 227792 423916 227798
rect 423864 227734 423916 227740
rect 424060 220862 424088 231662
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 221944 425020 221950
rect 424968 221886 425020 221892
rect 424048 220856 424100 220862
rect 424048 220798 424100 220804
rect 422680 219406 422892 219434
rect 423324 219406 423536 219434
rect 422680 219298 422708 219406
rect 422668 219292 422720 219298
rect 422668 219234 422720 219240
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 419966 217110 420040 217138
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 219406
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 221886
rect 425440 218210 425468 231662
rect 426452 225214 426480 231676
rect 426728 231662 427110 231690
rect 426440 225208 426492 225214
rect 426440 225150 426492 225156
rect 426728 220114 426756 231662
rect 427740 229158 427768 231676
rect 427924 231662 428398 231690
rect 428752 231662 429042 231690
rect 429212 231662 429686 231690
rect 429856 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432156 231662 432262 231690
rect 432616 231662 432906 231690
rect 433550 231662 433748 231690
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 426992 225208 427044 225214
rect 426992 225150 427044 225156
rect 426716 220108 426768 220114
rect 426716 220050 426768 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 225150
rect 427924 218210 427952 231662
rect 428752 219434 428780 231662
rect 429212 221950 429240 231662
rect 429200 221944 429252 221950
rect 429200 221886 429252 221892
rect 429856 219434 429884 231662
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 431960 220788 432012 220794
rect 431960 220730 432012 220736
rect 428280 219428 428332 219434
rect 428280 219370 428332 219376
rect 428476 219406 428780 219434
rect 429396 219406 429884 219434
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 427912 218204 427964 218210
rect 427912 218146 427964 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 219370
rect 428476 218074 428504 219406
rect 429396 218346 429424 219406
rect 429936 218612 429988 218618
rect 429936 218554 429988 218560
rect 429384 218340 429436 218346
rect 429384 218282 429436 218288
rect 428464 218068 428516 218074
rect 428464 218010 428516 218016
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217274 429148 218010
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217246 429148 217274
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217246
rect 429948 217138 429976 218554
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 220730
rect 432156 219570 432184 231662
rect 432144 219564 432196 219570
rect 432144 219506 432196 219512
rect 432616 219434 432644 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432156 219406 432644 219434
rect 432156 218618 432184 219406
rect 432144 218612 432196 218618
rect 432144 218554 432196 218560
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220794 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436324 231690
rect 434812 220788 434864 220794
rect 434812 220730 434864 220736
rect 434904 218340 434956 218346
rect 434904 218282 434956 218288
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218282
rect 435284 218210 435312 231662
rect 436100 230376 436152 230382
rect 436100 230318 436152 230324
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435732 218068 435784 218074
rect 435732 218010 435784 218016
rect 435744 217138 435772 218010
rect 436112 217258 436140 230318
rect 436296 218074 436324 231662
rect 436756 230382 436784 231676
rect 436940 231662 437414 231690
rect 437584 231662 438058 231690
rect 436744 230376 436796 230382
rect 436744 230318 436796 230324
rect 436940 219434 436968 231662
rect 437584 219434 437612 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 219434 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 219434 439360 230318
rect 436664 219406 436968 219434
rect 437492 219406 437612 219434
rect 438872 219406 438992 219434
rect 439056 219406 439360 219434
rect 436664 218346 436692 219406
rect 436652 218340 436704 218346
rect 436652 218282 436704 218288
rect 437492 218074 437520 219406
rect 438872 218074 438900 219406
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436560 218068 436612 218074
rect 436560 218010 436612 218016
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438216 218068 438268 218074
rect 438216 218010 438268 218016
rect 438860 218068 438912 218074
rect 438860 218010 438912 218016
rect 436100 217252 436152 217258
rect 436100 217194 436152 217200
rect 436572 217138 436600 218010
rect 437342 217252 437394 217258
rect 437342 217194 437394 217200
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436526 217110 436600 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217194
rect 438228 217138 438256 218010
rect 439056 217274 439084 219406
rect 440344 218074 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 218068 439924 218074
rect 439872 218010 439924 218016
rect 440332 218068 440384 218074
rect 440332 218010 440384 218016
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 218010
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441540 218062 441660 218090
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441540 217138 441568 218062
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230382 443868 231676
rect 443828 230376 443880 230382
rect 443828 230318 443880 230324
rect 444484 230246 444512 231676
rect 444668 231662 445142 231690
rect 444472 230240 444524 230246
rect 444472 230182 444524 230188
rect 444668 229094 444696 231662
rect 444840 230376 444892 230382
rect 444840 230318 444892 230324
rect 444852 229094 444880 230318
rect 445772 229094 445800 231676
rect 446416 230382 446444 231676
rect 446404 230376 446456 230382
rect 446404 230318 446456 230324
rect 443472 229066 443960 229094
rect 444668 229066 444788 229094
rect 444852 229066 445616 229094
rect 445772 229066 446444 229094
rect 443932 217274 443960 229066
rect 444760 217274 444788 229066
rect 445588 217274 445616 229066
rect 446416 217274 446444 229066
rect 447060 227934 447088 231676
rect 447520 231662 447718 231690
rect 447048 227928 447100 227934
rect 447048 227870 447100 227876
rect 447520 224534 447548 231662
rect 447692 230240 447744 230246
rect 447692 230182 447744 230188
rect 447508 224528 447560 224534
rect 447508 224470 447560 224476
rect 447704 219434 447732 230182
rect 448348 229094 448376 231676
rect 448704 230376 448756 230382
rect 448704 230318 448756 230324
rect 448716 229094 448744 230318
rect 448992 229566 449020 231676
rect 449636 230382 449664 231676
rect 449624 230376 449676 230382
rect 449624 230318 449676 230324
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 450280 229294 450308 231676
rect 450544 230376 450596 230382
rect 450544 230318 450596 230324
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 230318
rect 450924 229430 450952 231676
rect 451568 230246 451596 231676
rect 452226 231662 452608 231690
rect 451556 230240 451608 230246
rect 451556 230182 451608 230188
rect 451924 229560 451976 229566
rect 451924 229502 451976 229508
rect 450912 229424 450964 229430
rect 450912 229366 450964 229372
rect 451740 229288 451792 229294
rect 451740 229230 451792 229236
rect 448348 229066 448560 229094
rect 448716 229066 448928 229094
rect 450556 229066 450768 229094
rect 448060 224528 448112 224534
rect 448060 224470 448112 224476
rect 447336 219406 447732 219434
rect 447336 217274 447364 219406
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444760 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 441494 217110 441568 217138
rect 441494 216988 441522 217110
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447290 217246 447364 217274
rect 448072 217274 448100 224470
rect 448072 217246 448146 217274
rect 448532 217258 448560 229066
rect 448900 217274 448928 229066
rect 450544 227928 450596 227934
rect 450544 227870 450596 227876
rect 450556 217274 450584 227870
rect 450740 218346 450768 229066
rect 451752 219434 451780 229230
rect 451936 229094 451964 229502
rect 451936 229066 452240 229094
rect 451476 219406 451780 219434
rect 450728 218340 450780 218346
rect 450728 218282 450780 218288
rect 451476 217274 451504 219406
rect 447290 216988 447318 217246
rect 448118 216988 448146 217246
rect 448520 217252 448572 217258
rect 448900 217246 448974 217274
rect 448520 217194 448572 217200
rect 448946 216988 448974 217246
rect 449762 217252 449814 217258
rect 450556 217246 450630 217274
rect 449762 217194 449814 217200
rect 449774 216988 449802 217194
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 229066
rect 452580 222154 452608 231662
rect 452856 230382 452884 231676
rect 452844 230376 452896 230382
rect 452844 230318 452896 230324
rect 453500 230246 453528 231676
rect 453304 230240 453356 230246
rect 453304 230182 453356 230188
rect 453488 230240 453540 230246
rect 453488 230182 453540 230188
rect 453028 229424 453080 229430
rect 453028 229366 453080 229372
rect 452568 222148 452620 222154
rect 452568 222090 452620 222096
rect 453040 217274 453068 229366
rect 453316 218074 453344 230182
rect 454144 230110 454172 231676
rect 454316 230376 454368 230382
rect 454316 230318 454368 230324
rect 454132 230104 454184 230110
rect 454132 230046 454184 230052
rect 454328 229094 454356 230318
rect 454788 229094 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455788 230240 455840 230246
rect 455788 230182 455840 230188
rect 455328 230104 455380 230110
rect 455328 230046 455380 230052
rect 454328 229066 454724 229094
rect 454788 229066 454908 229094
rect 453856 218340 453908 218346
rect 453856 218282 453908 218288
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 218282
rect 454696 217274 454724 229066
rect 454880 223582 454908 229066
rect 454868 223576 454920 223582
rect 454868 223518 454920 223524
rect 455340 220726 455368 230046
rect 455604 222148 455656 222154
rect 455604 222090 455656 222096
rect 455328 220720 455380 220726
rect 455328 220662 455380 220668
rect 455616 218074 455644 222090
rect 455800 219434 455828 230182
rect 456076 224534 456104 231676
rect 456064 224528 456116 224534
rect 456064 224470 456116 224476
rect 456720 220862 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 220856 456760 220862
rect 456708 220798 456760 220804
rect 457180 219434 457208 230318
rect 457364 229906 457392 231676
rect 457352 229900 457404 229906
rect 457352 229842 457404 229848
rect 458008 229094 458036 231676
rect 458008 229066 458128 229094
rect 455800 219406 456380 219434
rect 457180 219406 458036 219434
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455604 218068 455656 218074
rect 455604 218010 455656 218016
rect 455432 217274 455460 218010
rect 456352 217274 456380 219406
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 454696 217246 454770 217274
rect 455432 217246 455598 217274
rect 456352 217246 456426 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458100 218498 458128 229066
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 458824 220720 458876 220726
rect 458824 220662 458876 220668
rect 458100 218470 458220 218498
rect 458192 218414 458220 218470
rect 458180 218408 458232 218414
rect 458180 218350 458232 218356
rect 458836 217274 458864 220662
rect 459480 220250 459508 231662
rect 459744 224528 459796 224534
rect 459744 224470 459796 224476
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217274 459784 224470
rect 459940 222902 459968 231676
rect 460584 223718 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 223712 460624 223718
rect 460572 223654 460624 223660
rect 460480 223576 460532 223582
rect 460480 223518 460532 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 217246 459784 217274
rect 460492 217274 460520 223518
rect 461308 218340 461360 218346
rect 461308 218282 461360 218288
rect 460492 217246 460566 217274
rect 459710 216988 459738 217246
rect 460538 216988 460566 217246
rect 461320 217138 461348 218282
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224806 462544 231676
rect 462964 225820 463016 225826
rect 462964 225762 463016 225768
rect 462504 224800 462556 224806
rect 462504 224742 462556 224748
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 220856 462188 220862
rect 462136 220798 462188 220804
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 220798
rect 462976 217274 463004 225762
rect 463160 225418 463188 231676
rect 463804 229634 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 464068 229900 464120 229906
rect 464068 229842 464120 229848
rect 463792 229628 463844 229634
rect 463792 229570 463844 229576
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 223712 463200 223718
rect 463148 223654 463200 223660
rect 463160 218074 463188 223654
rect 464080 219434 464108 229842
rect 465000 219638 465028 231662
rect 465460 229498 465488 231662
rect 465724 229628 465776 229634
rect 465724 229570 465776 229576
rect 465448 229492 465500 229498
rect 465448 229434 465500 229440
rect 465736 220726 465764 229570
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220862 466132 231662
rect 467024 229770 467052 231676
rect 467012 229764 467064 229770
rect 467012 229706 467064 229712
rect 467472 229492 467524 229498
rect 467472 229434 467524 229440
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 463896 219406 464108 219434
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 219406
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 461320 217110 461394 217138
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229434
rect 467668 225622 467696 231676
rect 468312 230246 468340 231676
rect 468300 230240 468352 230246
rect 468300 230182 468352 230188
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 468956 221474 468984 231676
rect 469128 230240 469180 230246
rect 469128 230182 469180 230188
rect 468944 221468 468996 221474
rect 468944 221410 468996 221416
rect 469140 220522 469168 230182
rect 469600 229906 469628 231676
rect 469588 229900 469640 229906
rect 469588 229842 469640 229848
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224800 469364 224806
rect 469312 224742 469364 224748
rect 469128 220516 469180 220522
rect 469128 220458 469180 220464
rect 468772 217246 468846 217274
rect 469324 217258 469352 224742
rect 469588 220720 469640 220726
rect 469588 220662 469640 220668
rect 469600 217274 469628 220662
rect 469876 218618 469904 227598
rect 470244 224262 470272 231676
rect 470888 230382 470916 231676
rect 470876 230376 470928 230382
rect 470876 230318 470928 230324
rect 471532 227798 471560 231676
rect 472176 230382 472204 231676
rect 472834 231662 473032 231690
rect 471888 230376 471940 230382
rect 471888 230318 471940 230324
rect 472164 230376 472216 230382
rect 472164 230318 472216 230324
rect 471520 227792 471572 227798
rect 471520 227734 471572 227740
rect 470232 224256 470284 224262
rect 470232 224198 470284 224204
rect 471900 222154 471928 230318
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471336 220856 471388 220862
rect 471336 220798 471388 220804
rect 471348 218754 471376 220798
rect 473004 220250 473032 231662
rect 473176 230376 473228 230382
rect 473176 230318 473228 230324
rect 473188 220386 473216 230318
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474004 229764 474056 229770
rect 474004 229706 474056 229712
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 473176 220380 473228 220386
rect 473176 220322 473228 220328
rect 472992 220244 473044 220250
rect 472992 220186 473044 220192
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471336 218748 471388 218754
rect 471336 218690 471388 218696
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 472084 217274 472112 219574
rect 472900 218748 472952 218754
rect 472900 218690 472952 218696
rect 472912 217274 472940 218690
rect 473740 217274 473768 222838
rect 474016 220794 474044 229706
rect 474476 228410 474504 231662
rect 474464 228404 474516 228410
rect 474464 228346 474516 228352
rect 474752 226506 474780 231676
rect 475410 231662 475884 231690
rect 474740 226500 474792 226506
rect 474740 226442 474792 226448
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 474004 220788 474056 220794
rect 474004 220730 474056 220736
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474556 220516 474608 220522
rect 474556 220458 474608 220464
rect 474568 217274 474596 220458
rect 475396 217274 475424 220730
rect 475580 218618 475608 223518
rect 475856 221610 475884 231662
rect 476040 229838 476068 231676
rect 476684 230042 476712 231676
rect 476672 230036 476724 230042
rect 476672 229978 476724 229984
rect 476028 229832 476080 229838
rect 476028 229774 476080 229780
rect 476764 229696 476816 229702
rect 476764 229638 476816 229644
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475844 221604 475896 221610
rect 475844 221546 475896 221552
rect 476212 221468 476264 221474
rect 476212 221410 476264 221416
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 221410
rect 476592 217274 476620 225558
rect 476776 220794 476804 229638
rect 477328 225622 477356 231676
rect 477986 231662 478368 231690
rect 478630 231662 478828 231690
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478340 220114 478368 231662
rect 478604 229832 478656 229838
rect 478604 229774 478656 229780
rect 478616 227186 478644 229774
rect 478800 229094 478828 231662
rect 479260 229770 479288 231676
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 478800 229066 478920 229094
rect 478892 228818 478920 229066
rect 478880 228812 478932 228818
rect 478880 228754 478932 228760
rect 479524 227792 479576 227798
rect 479524 227734 479576 227740
rect 478604 227180 478656 227186
rect 478604 227122 478656 227128
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478328 220108 478380 220114
rect 478328 220050 478380 220056
rect 478708 217274 478736 220730
rect 479536 217274 479564 227734
rect 479904 222902 479932 231676
rect 480548 224398 480576 231676
rect 481192 225758 481220 231676
rect 481640 230036 481692 230042
rect 481640 229978 481692 229984
rect 481652 226370 481680 229978
rect 481836 229906 481864 231676
rect 482494 231662 482968 231690
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 482744 226500 482796 226506
rect 482744 226442 482796 226448
rect 481640 226364 481692 226370
rect 481640 226306 481692 226312
rect 481180 225752 481232 225758
rect 481180 225694 481232 225700
rect 480536 224392 480588 224398
rect 480536 224334 480588 224340
rect 480352 224256 480404 224262
rect 480352 224198 480404 224204
rect 479892 222896 479944 222902
rect 479892 222838 479944 222844
rect 480364 217274 480392 224198
rect 482756 222630 482784 226442
rect 482744 222624 482796 222630
rect 482744 222566 482796 222572
rect 481180 220380 481232 220386
rect 481180 220322 481232 220328
rect 481192 217274 481220 220322
rect 482008 220244 482060 220250
rect 482008 220186 482060 220192
rect 482020 217274 482048 220186
rect 482756 218754 482784 222566
rect 482940 220250 482968 231662
rect 483124 223174 483152 231676
rect 483768 224262 483796 231676
rect 484426 231662 484808 231690
rect 484584 228404 484636 228410
rect 484584 228346 484636 228352
rect 483756 224256 483808 224262
rect 483756 224198 483808 224204
rect 483112 223168 483164 223174
rect 483112 223110 483164 223116
rect 484596 222358 484624 228346
rect 484584 222352 484636 222358
rect 484584 222294 484636 222300
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 482928 220244 482980 220250
rect 482928 220186 482980 220192
rect 482744 218748 482796 218754
rect 482744 218690 482796 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 472084 217246 472158 217274
rect 472912 217246 472986 217274
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 480364 217246 480438 217274
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472958 216988 472986 217246
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480410 216988 480438 217246
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 484596 217274 484624 222294
rect 484780 221746 484808 231662
rect 485056 228410 485084 231676
rect 485700 228546 485728 231676
rect 486358 231662 486648 231690
rect 485688 228540 485740 228546
rect 485688 228482 485740 228488
rect 485044 228404 485096 228410
rect 485044 228346 485096 228352
rect 486620 223038 486648 231662
rect 486792 227180 486844 227186
rect 486792 227122 486844 227128
rect 486608 223032 486660 223038
rect 486608 222974 486660 222980
rect 484768 221740 484820 221746
rect 484768 221682 484820 221688
rect 486148 221604 486200 221610
rect 486148 221546 486200 221552
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 483722 217246 483796 217274
rect 484550 217246 484624 217274
rect 485332 217274 485360 218690
rect 486160 217274 486188 221546
rect 486804 219434 486832 227122
rect 486988 227050 487016 231676
rect 487632 230382 487660 231676
rect 487620 230376 487672 230382
rect 487620 230318 487672 230324
rect 488080 229764 488132 229770
rect 488080 229706 488132 229712
rect 486976 227044 487028 227050
rect 486976 226986 487028 226992
rect 488092 226370 488120 229706
rect 488276 229498 488304 231676
rect 488934 231662 489408 231690
rect 488448 230376 488500 230382
rect 488448 230318 488500 230324
rect 488264 229492 488316 229498
rect 488264 229434 488316 229440
rect 487804 226364 487856 226370
rect 487804 226306 487856 226312
rect 488080 226364 488132 226370
rect 488080 226306 488132 226312
rect 486974 219464 487030 219473
rect 486804 219408 486974 219434
rect 486804 219406 487030 219408
rect 486974 219399 487030 219406
rect 486988 217274 487016 219399
rect 487816 218113 487844 226306
rect 488460 220522 488488 230318
rect 489380 225622 489408 231662
rect 489564 229094 489592 231676
rect 490208 230246 490236 231676
rect 490866 231662 491248 231690
rect 490196 230240 490248 230246
rect 490196 230182 490248 230188
rect 489920 229900 489972 229906
rect 489920 229842 489972 229848
rect 489564 229066 489684 229094
rect 488724 225616 488776 225622
rect 488724 225558 488776 225564
rect 489368 225616 489420 225622
rect 489368 225558 489420 225564
rect 488448 220516 488500 220522
rect 488448 220458 488500 220464
rect 487802 218104 487858 218113
rect 487802 218039 487858 218048
rect 487816 217274 487844 218039
rect 488736 217274 488764 225558
rect 489656 220114 489684 229066
rect 489932 227798 489960 229842
rect 490380 229492 490432 229498
rect 490380 229434 490432 229440
rect 490196 228812 490248 228818
rect 490196 228754 490248 228760
rect 489920 227792 489972 227798
rect 489920 227734 489972 227740
rect 490012 226364 490064 226370
rect 490012 226306 490064 226312
rect 490024 222426 490052 226306
rect 490012 222420 490064 222426
rect 490012 222362 490064 222368
rect 489460 220108 489512 220114
rect 489460 220050 489512 220056
rect 489644 220108 489696 220114
rect 489644 220050 489696 220056
rect 485332 217246 485406 217274
rect 486160 217246 486234 217274
rect 486988 217246 487062 217274
rect 487816 217246 487890 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485378 216988 485406 217246
rect 486206 216988 486234 217246
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488690 217246 488764 217274
rect 489472 217274 489500 220050
rect 490024 219434 490052 222362
rect 489932 219406 490052 219434
rect 490208 219434 490236 228754
rect 490392 227186 490420 229434
rect 491220 229094 491248 231662
rect 491496 230110 491524 231676
rect 491484 230104 491536 230110
rect 491484 230046 491536 230052
rect 492140 229770 492168 231676
rect 492798 231662 493088 231690
rect 492496 230104 492548 230110
rect 492496 230046 492548 230052
rect 492128 229764 492180 229770
rect 492128 229706 492180 229712
rect 491220 229066 491340 229094
rect 490380 227180 490432 227186
rect 490380 227122 490432 227128
rect 491312 224534 491340 229066
rect 491300 224528 491352 224534
rect 491300 224470 491352 224476
rect 492036 222896 492088 222902
rect 492036 222838 492088 222844
rect 490208 219406 490420 219434
rect 489472 217246 489546 217274
rect 489932 217258 489960 219406
rect 490392 218657 490420 219406
rect 490378 218648 490434 218657
rect 490378 218583 490434 218592
rect 490392 217274 490420 218583
rect 492048 218074 492076 222838
rect 492508 221882 492536 230046
rect 492680 225752 492732 225758
rect 492680 225694 492732 225700
rect 492496 221876 492548 221882
rect 492496 221818 492548 221824
rect 492692 218929 492720 225694
rect 492864 224392 492916 224398
rect 492864 224334 492916 224340
rect 492678 218920 492734 218929
rect 492678 218855 492734 218864
rect 492036 218068 492088 218074
rect 492036 218010 492088 218016
rect 488690 217161 488718 217246
rect 488676 217152 488732 217161
rect 488676 217087 488732 217096
rect 488690 216988 488718 217087
rect 489518 216988 489546 217246
rect 489920 217252 489972 217258
rect 489920 217194 489972 217200
rect 490346 217246 490420 217274
rect 491162 217252 491214 217258
rect 490346 216988 490374 217246
rect 491162 217194 491214 217200
rect 491174 216988 491202 217194
rect 492048 217138 492076 218010
rect 492876 217274 492904 224334
rect 493060 223310 493088 231662
rect 493428 230382 493456 231676
rect 493416 230376 493468 230382
rect 493416 230318 493468 230324
rect 493692 230240 493744 230246
rect 493692 230182 493744 230188
rect 493704 225758 493732 230182
rect 493692 225752 493744 225758
rect 493692 225694 493744 225700
rect 494072 224670 494100 231676
rect 494520 227792 494572 227798
rect 494520 227734 494572 227740
rect 494060 224664 494112 224670
rect 494060 224606 494112 224612
rect 493048 223304 493100 223310
rect 493048 223246 493100 223252
rect 494532 219434 494560 227734
rect 494716 227458 494744 231676
rect 495360 229294 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 229288 495400 229294
rect 495348 229230 495400 229236
rect 496188 229094 496216 231662
rect 497292 230382 497320 231676
rect 497476 231662 497950 231690
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 497280 230376 497332 230382
rect 497280 230318 497332 230324
rect 496372 229094 496400 230318
rect 497476 229094 497504 231662
rect 498108 230376 498160 230382
rect 498108 230318 498160 230324
rect 496188 229066 496308 229094
rect 496372 229066 496492 229094
rect 497476 229066 497688 229094
rect 494704 227452 494756 227458
rect 494704 227394 494756 227400
rect 496084 223168 496136 223174
rect 496084 223110 496136 223116
rect 495348 220244 495400 220250
rect 495348 220186 495400 220192
rect 494532 219406 494744 219434
rect 494716 218929 494744 219406
rect 493782 218920 493838 218929
rect 494702 218920 494758 218929
rect 493782 218855 493838 218864
rect 494532 218878 494702 218906
rect 493796 217297 493824 218855
rect 492002 217110 492076 217138
rect 492830 217246 492904 217274
rect 493782 217288 493838 217297
rect 492002 216988 492030 217110
rect 492830 216988 492858 217246
rect 494532 217274 494560 218878
rect 494702 218855 494758 218864
rect 495360 217297 495388 220186
rect 493782 217223 493838 217232
rect 494486 217246 494560 217274
rect 495346 217288 495402 217297
rect 493796 217138 493824 217223
rect 493658 217110 493824 217138
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 496096 217274 496124 223110
rect 496280 221610 496308 229066
rect 496268 221604 496320 221610
rect 496268 221546 496320 221552
rect 496464 220386 496492 229066
rect 497464 224256 497516 224262
rect 497464 224198 497516 224204
rect 496452 220380 496504 220386
rect 496452 220322 496504 220328
rect 497476 218657 497504 224198
rect 497660 220250 497688 229066
rect 498120 226030 498148 230318
rect 498580 228682 498608 231676
rect 498568 228676 498620 228682
rect 498568 228618 498620 228624
rect 498292 228540 498344 228546
rect 498292 228482 498344 228488
rect 498108 226024 498160 226030
rect 498108 225966 498160 225972
rect 497832 221740 497884 221746
rect 497832 221682 497884 221688
rect 497844 220969 497872 221682
rect 497830 220960 497886 220969
rect 497830 220895 497886 220904
rect 497648 220244 497700 220250
rect 497648 220186 497700 220192
rect 497844 219434 497872 220895
rect 498304 219434 498332 228482
rect 498568 228404 498620 228410
rect 498568 228346 498620 228352
rect 497752 219406 497872 219434
rect 498212 219406 498332 219434
rect 497462 218648 497518 218657
rect 497462 218583 497518 218592
rect 497476 217274 497504 218583
rect 496096 217246 496170 217274
rect 495346 217223 495402 217232
rect 495360 217138 495388 217223
rect 495314 217110 495388 217138
rect 495314 216988 495342 217110
rect 496142 216988 496170 217246
rect 496970 217246 497504 217274
rect 497752 217274 497780 219406
rect 497752 217246 497826 217274
rect 498212 217258 498240 219406
rect 498580 217297 498608 228346
rect 499224 224398 499252 231676
rect 499868 228546 499896 231676
rect 500526 231662 500816 231690
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 499856 228540 499908 228546
rect 499856 228482 499908 228488
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 500236 220794 500264 229230
rect 500408 223032 500460 223038
rect 500408 222974 500460 222980
rect 500224 220788 500276 220794
rect 500224 220730 500276 220736
rect 500420 218346 500448 222974
rect 500788 222902 500816 231662
rect 500960 227044 501012 227050
rect 500960 226986 501012 226992
rect 500776 222896 500828 222902
rect 500776 222838 500828 222844
rect 500972 220368 501000 226986
rect 501156 225894 501184 231676
rect 501340 231662 501814 231690
rect 501144 225888 501196 225894
rect 501144 225830 501196 225836
rect 501340 221746 501368 231662
rect 502444 228954 502472 231676
rect 503102 231662 503392 231690
rect 502432 228948 502484 228954
rect 502432 228890 502484 228896
rect 502984 227180 503036 227186
rect 502984 227122 503036 227128
rect 502432 222488 502484 222494
rect 502432 222430 502484 222436
rect 502444 222222 502472 222430
rect 502432 222216 502484 222222
rect 502432 222158 502484 222164
rect 501328 221740 501380 221746
rect 501328 221682 501380 221688
rect 501880 220516 501932 220522
rect 501880 220458 501932 220464
rect 500972 220340 501184 220368
rect 501156 219570 501184 220340
rect 501144 219564 501196 219570
rect 501144 219506 501196 219512
rect 500408 218340 500460 218346
rect 500408 218282 500460 218288
rect 498566 217288 498622 217297
rect 496970 216988 496998 217246
rect 497798 216988 497826 217246
rect 498200 217252 498252 217258
rect 500420 217274 500448 218282
rect 501156 217274 501184 219506
rect 498566 217223 498622 217232
rect 499442 217252 499494 217258
rect 498200 217194 498252 217200
rect 498580 217138 498608 217223
rect 499442 217194 499494 217200
rect 500282 217246 500448 217274
rect 501110 217246 501184 217274
rect 501892 217274 501920 220458
rect 502996 218210 503024 227122
rect 503168 225616 503220 225622
rect 503168 225558 503220 225564
rect 502984 218204 503036 218210
rect 502984 218146 503036 218152
rect 502996 217274 503024 218146
rect 501892 217246 501966 217274
rect 498580 217110 498654 217138
rect 498626 216988 498654 217110
rect 499454 216988 499482 217194
rect 500282 216988 500310 217246
rect 501110 216988 501138 217246
rect 501938 216988 501966 217246
rect 502766 217246 503024 217274
rect 502766 216988 502794 217246
rect 503180 217122 503208 225558
rect 503364 223174 503392 231662
rect 503732 229158 503760 231676
rect 503720 229152 503772 229158
rect 503720 229094 503772 229100
rect 504376 224126 504404 231676
rect 505020 227186 505048 231676
rect 505192 229764 505244 229770
rect 505192 229706 505244 229712
rect 505008 227180 505060 227186
rect 505008 227122 505060 227128
rect 504364 224120 504416 224126
rect 504364 224062 504416 224068
rect 505204 223786 505232 229706
rect 505664 229294 505692 231676
rect 505652 229288 505704 229294
rect 505652 229230 505704 229236
rect 506308 227050 506336 231676
rect 506572 229900 506624 229906
rect 506572 229842 506624 229848
rect 506584 228410 506612 229842
rect 506572 228404 506624 228410
rect 506572 228346 506624 228352
rect 506296 227044 506348 227050
rect 506296 226986 506348 226992
rect 505376 225752 505428 225758
rect 505376 225694 505428 225700
rect 505192 223780 505244 223786
rect 505192 223722 505244 223728
rect 505388 223650 505416 225694
rect 506952 224806 506980 231676
rect 507596 229770 507624 231676
rect 507584 229764 507636 229770
rect 507584 229706 507636 229712
rect 506940 224800 506992 224806
rect 506940 224742 506992 224748
rect 506020 224528 506072 224534
rect 506020 224470 506072 224476
rect 505376 223644 505428 223650
rect 505376 223586 505428 223592
rect 503352 223168 503404 223174
rect 503352 223110 503404 223116
rect 504364 220108 504416 220114
rect 504364 220050 504416 220056
rect 504376 217274 504404 220050
rect 505388 217274 505416 223586
rect 506032 219774 506060 224470
rect 507676 223780 507728 223786
rect 507676 223722 507728 223728
rect 506848 221876 506900 221882
rect 506848 221818 506900 221824
rect 506020 219768 506072 219774
rect 506020 219710 506072 219716
rect 505652 218068 505704 218074
rect 505652 218010 505704 218016
rect 505664 217569 505692 218010
rect 505650 217560 505706 217569
rect 505650 217495 505706 217504
rect 504376 217246 504450 217274
rect 503168 217116 503220 217122
rect 503168 217058 503220 217064
rect 503582 217116 503634 217122
rect 503582 217058 503634 217064
rect 503594 216988 503622 217058
rect 504422 216988 504450 217246
rect 505250 217246 505416 217274
rect 505250 216988 505278 217246
rect 506032 217138 506060 219710
rect 506860 217138 506888 221818
rect 507688 218074 507716 223722
rect 508240 223038 508268 231676
rect 508884 225758 508912 231676
rect 509528 229634 509556 231676
rect 509516 229628 509568 229634
rect 509516 229570 509568 229576
rect 509884 229152 509936 229158
rect 509884 229094 509936 229100
rect 508872 225752 508924 225758
rect 508872 225694 508924 225700
rect 508504 223304 508556 223310
rect 508504 223246 508556 223252
rect 508228 223032 508280 223038
rect 508228 222974 508280 222980
rect 507676 218068 507728 218074
rect 507676 218010 507728 218016
rect 507688 217138 507716 218010
rect 508516 217841 508544 223246
rect 509896 220658 509924 229094
rect 510172 225622 510200 231676
rect 510816 229906 510844 231676
rect 511460 230382 511488 231676
rect 511448 230376 511500 230382
rect 511448 230318 511500 230324
rect 510804 229900 510856 229906
rect 510804 229842 510856 229848
rect 511908 229900 511960 229906
rect 511908 229842 511960 229848
rect 510620 229288 510672 229294
rect 510620 229230 510672 229236
rect 510632 227322 510660 229230
rect 511920 229094 511948 229842
rect 511644 229066 511948 229094
rect 511080 227452 511132 227458
rect 511080 227394 511132 227400
rect 510620 227316 510672 227322
rect 510620 227258 510672 227264
rect 510160 225616 510212 225622
rect 510160 225558 510212 225564
rect 510160 224664 510212 224670
rect 510160 224606 510212 224612
rect 509884 220652 509936 220658
rect 509884 220594 509936 220600
rect 509332 220380 509384 220386
rect 509332 220322 509384 220328
rect 508502 217832 508558 217841
rect 508502 217767 508558 217776
rect 508516 217138 508544 217767
rect 509344 217274 509372 220322
rect 510172 217841 510200 224606
rect 510158 217832 510214 217841
rect 510158 217767 510214 217776
rect 509344 217246 509418 217274
rect 506032 217110 506106 217138
rect 506860 217110 506934 217138
rect 507688 217110 507762 217138
rect 508516 217110 508590 217138
rect 506078 216988 506106 217110
rect 506906 216988 506934 217110
rect 507734 216988 507762 217110
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510172 217138 510200 217767
rect 511092 217274 511120 227394
rect 511644 220522 511672 229066
rect 512104 228410 512132 231676
rect 512762 231662 513144 231690
rect 512092 228404 512144 228410
rect 512092 228346 512144 228352
rect 512736 228268 512788 228274
rect 512736 228210 512788 228216
rect 511816 220788 511868 220794
rect 511816 220730 511868 220736
rect 511632 220516 511684 220522
rect 511632 220458 511684 220464
rect 511046 217246 511120 217274
rect 511046 217190 511074 217246
rect 511034 217184 511086 217190
rect 510172 217110 510246 217138
rect 511034 217126 511086 217132
rect 511828 217138 511856 220730
rect 512748 218482 512776 228210
rect 513116 220114 513144 231662
rect 513392 229294 513420 231676
rect 513380 229288 513432 229294
rect 513380 229230 513432 229236
rect 514036 227458 514064 231676
rect 514024 227452 514076 227458
rect 514024 227394 514076 227400
rect 514300 226024 514352 226030
rect 514300 225966 514352 225972
rect 513378 221640 513434 221649
rect 513378 221575 513380 221584
rect 513432 221575 513434 221584
rect 513380 221546 513432 221552
rect 513104 220108 513156 220114
rect 513104 220050 513156 220056
rect 512736 218476 512788 218482
rect 512736 218418 512788 218424
rect 512748 217274 512776 218418
rect 512702 217246 512776 217274
rect 513392 217274 513420 221546
rect 514312 217274 514340 225966
rect 514680 223310 514708 231676
rect 515324 230042 515352 231676
rect 515312 230036 515364 230042
rect 515312 229978 515364 229984
rect 515404 229628 515456 229634
rect 515404 229570 515456 229576
rect 514668 223304 514720 223310
rect 514668 223246 514720 223252
rect 515416 220386 515444 229570
rect 515772 228676 515824 228682
rect 515772 228618 515824 228624
rect 515784 220862 515812 228618
rect 515968 224534 515996 231676
rect 516612 226030 516640 231676
rect 517256 229906 517284 231676
rect 517520 230376 517572 230382
rect 517520 230318 517572 230324
rect 517244 229900 517296 229906
rect 517244 229842 517296 229848
rect 516784 229764 516836 229770
rect 516784 229706 516836 229712
rect 516796 229094 516824 229706
rect 516796 229066 517008 229094
rect 516600 226024 516652 226030
rect 516600 225966 516652 225972
rect 515956 224528 516008 224534
rect 515956 224470 516008 224476
rect 516784 224392 516836 224398
rect 516784 224334 516836 224340
rect 515772 220856 515824 220862
rect 515772 220798 515824 220804
rect 515404 220380 515456 220386
rect 515404 220322 515456 220328
rect 515220 220244 515272 220250
rect 515220 220186 515272 220192
rect 515232 219745 515260 220186
rect 515218 219736 515274 219745
rect 515218 219671 515274 219680
rect 515232 217274 515260 219671
rect 515784 219434 515812 220798
rect 515784 219406 515996 219434
rect 513392 217246 513558 217274
rect 514312 217246 514386 217274
rect 510218 216988 510246 217110
rect 511046 216988 511074 217126
rect 511828 217110 511902 217138
rect 511874 216988 511902 217110
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515186 217246 515260 217274
rect 515968 217274 515996 219406
rect 516796 217274 516824 224334
rect 516980 221610 517008 229066
rect 517532 223446 517560 230318
rect 517900 228682 517928 231676
rect 518544 228818 518572 231676
rect 519188 229158 519216 231676
rect 519360 229288 519412 229294
rect 519360 229230 519412 229236
rect 519176 229152 519228 229158
rect 519176 229094 519228 229100
rect 518532 228812 518584 228818
rect 518532 228754 518584 228760
rect 517888 228676 517940 228682
rect 517888 228618 517940 228624
rect 517704 228540 517756 228546
rect 517704 228482 517756 228488
rect 517716 223786 517744 228482
rect 519176 225888 519228 225894
rect 519176 225830 519228 225836
rect 517704 223780 517756 223786
rect 517704 223722 517756 223728
rect 517520 223440 517572 223446
rect 517520 223382 517572 223388
rect 517520 222896 517572 222902
rect 517520 222838 517572 222844
rect 516968 221604 517020 221610
rect 516968 221546 517020 221552
rect 517532 221134 517560 222838
rect 517520 221128 517572 221134
rect 517520 221070 517572 221076
rect 517716 219434 517744 223722
rect 518440 221128 518492 221134
rect 518440 221070 518492 221076
rect 517624 219406 517744 219434
rect 517624 217274 517652 219406
rect 518452 217274 518480 221070
rect 519188 219434 519216 225830
rect 519372 224942 519400 229230
rect 519360 224936 519412 224942
rect 519360 224878 519412 224884
rect 519832 222902 519860 231676
rect 520476 224670 520504 231676
rect 521120 230178 521148 231676
rect 521108 230172 521160 230178
rect 521108 230114 521160 230120
rect 521016 228948 521068 228954
rect 521016 228890 521068 228896
rect 520464 224664 520516 224670
rect 520464 224606 520516 224612
rect 519820 222896 519872 222902
rect 519820 222838 519872 222844
rect 520188 221808 520240 221814
rect 520188 221750 520240 221756
rect 520200 221241 520228 221750
rect 520186 221232 520242 221241
rect 520186 221167 520242 221176
rect 519188 219406 519308 219434
rect 519280 217274 519308 219406
rect 520200 217274 520228 221167
rect 521028 220998 521056 228890
rect 521764 225894 521792 231676
rect 522422 231662 522712 231690
rect 521752 225888 521804 225894
rect 521752 225830 521804 225836
rect 521752 223168 521804 223174
rect 521752 223110 521804 223116
rect 521016 220992 521068 220998
rect 521016 220934 521068 220940
rect 521028 217274 521056 220934
rect 515968 217246 516042 217274
rect 516796 217246 516870 217274
rect 517624 217246 517698 217274
rect 518452 217246 518526 217274
rect 519280 217246 519354 217274
rect 515186 216988 515214 217246
rect 516014 216988 516042 217246
rect 516842 216988 516870 217246
rect 517670 216988 517698 217246
rect 518498 216988 518526 217246
rect 519326 216988 519354 217246
rect 520154 217246 520228 217274
rect 520982 217246 521056 217274
rect 521764 217274 521792 223110
rect 522684 221882 522712 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523696 227186 523724 231676
rect 524248 231662 524354 231690
rect 523040 227180 523092 227186
rect 523040 227122 523092 227128
rect 523684 227180 523736 227186
rect 523684 227122 523736 227128
rect 522672 221876 522724 221882
rect 522672 221818 522724 221824
rect 522580 220652 522632 220658
rect 522580 220594 522632 220600
rect 522592 217841 522620 220594
rect 523052 217870 523080 227122
rect 523500 224256 523552 224262
rect 523500 224198 523552 224204
rect 523512 221270 523540 224198
rect 524248 221746 524276 231662
rect 524604 230036 524656 230042
rect 524604 229978 524656 229984
rect 524616 227594 524644 229978
rect 524984 229158 525012 231676
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524604 227588 524656 227594
rect 524604 227530 524656 227536
rect 524420 227316 524472 227322
rect 524420 227258 524472 227264
rect 524432 223922 524460 227258
rect 525628 224398 525656 231676
rect 525984 229900 526036 229906
rect 525984 229842 526036 229848
rect 525996 226166 526024 229842
rect 526272 227322 526300 231676
rect 526916 230450 526944 231676
rect 526904 230444 526956 230450
rect 526904 230386 526956 230392
rect 527560 228546 527588 231676
rect 528218 231662 528416 231690
rect 527548 228540 527600 228546
rect 527548 228482 527600 228488
rect 526260 227316 526312 227322
rect 526260 227258 526312 227264
rect 526536 227044 526588 227050
rect 526536 226986 526588 226992
rect 525984 226160 526036 226166
rect 525984 226102 526036 226108
rect 526352 224800 526404 224806
rect 526352 224742 526404 224748
rect 525616 224392 525668 224398
rect 525616 224334 525668 224340
rect 524420 223916 524472 223922
rect 524420 223858 524472 223864
rect 525064 223916 525116 223922
rect 525064 223858 525116 223864
rect 524236 221740 524288 221746
rect 524236 221682 524288 221688
rect 523500 221264 523552 221270
rect 523500 221206 523552 221212
rect 523040 217864 523092 217870
rect 522578 217832 522634 217841
rect 523040 217806 523092 217812
rect 522578 217767 522634 217776
rect 521764 217246 521838 217274
rect 520154 216988 520182 217246
rect 520982 216988 521010 217246
rect 521810 216988 521838 217246
rect 522592 217138 522620 217767
rect 523512 217274 523540 221206
rect 524236 217864 524288 217870
rect 524236 217806 524288 217812
rect 523466 217246 523540 217274
rect 522592 217110 522666 217138
rect 522638 216988 522666 217110
rect 523466 216988 523494 217246
rect 524248 217138 524276 217806
rect 525076 217274 525104 223858
rect 525984 217728 526036 217734
rect 525984 217670 526036 217676
rect 525996 217274 526024 217670
rect 525076 217246 525150 217274
rect 524248 217110 524322 217138
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 217246 526024 217274
rect 526364 217274 526392 224742
rect 526548 217734 526576 226986
rect 527180 223032 527232 223038
rect 527180 222974 527232 222980
rect 527192 222086 527220 222974
rect 527180 222080 527232 222086
rect 527180 222022 527232 222028
rect 528192 222080 528244 222086
rect 528192 222022 528244 222028
rect 527548 221604 527600 221610
rect 527548 221546 527600 221552
rect 527560 219638 527588 221546
rect 527548 219632 527600 219638
rect 527548 219574 527600 219580
rect 526536 217728 526588 217734
rect 526536 217670 526588 217676
rect 526548 217462 526576 217670
rect 526536 217456 526588 217462
rect 526536 217398 526588 217404
rect 527560 217274 527588 219574
rect 528204 219434 528232 222022
rect 528388 220250 528416 231662
rect 528848 230314 528876 231676
rect 528836 230308 528888 230314
rect 528836 230250 528888 230256
rect 529204 230172 529256 230178
rect 529204 230114 529256 230120
rect 529216 229094 529244 230114
rect 529032 229066 529244 229094
rect 529032 220658 529060 229066
rect 529204 225752 529256 225758
rect 529204 225694 529256 225700
rect 529020 220652 529072 220658
rect 529020 220594 529072 220600
rect 528376 220244 528428 220250
rect 528376 220186 528428 220192
rect 528204 219406 528416 219434
rect 528388 217274 528416 219406
rect 529216 217274 529244 225694
rect 529492 223174 529520 231676
rect 530136 229634 530164 231676
rect 530124 229628 530176 229634
rect 530124 229570 530176 229576
rect 530780 229498 530808 231676
rect 531136 229628 531188 229634
rect 531136 229570 531188 229576
rect 530768 229492 530820 229498
rect 530768 229434 530820 229440
rect 529940 229152 529992 229158
rect 529940 229094 529992 229100
rect 529952 224806 529980 229094
rect 530584 225616 530636 225622
rect 530584 225558 530636 225564
rect 529940 224800 529992 224806
rect 529940 224742 529992 224748
rect 529480 223168 529532 223174
rect 529480 223110 529532 223116
rect 530032 220380 530084 220386
rect 530032 220322 530084 220328
rect 530044 219910 530072 220322
rect 530032 219904 530084 219910
rect 530032 219846 530084 219852
rect 530044 217274 530072 219846
rect 530596 217598 530624 225558
rect 531148 220386 531176 229570
rect 531424 225622 531452 231676
rect 531412 225616 531464 225622
rect 531412 225558 531464 225564
rect 532068 223038 532096 231676
rect 532712 230178 532740 231676
rect 532700 230172 532752 230178
rect 532700 230114 532752 230120
rect 533356 227050 533384 231676
rect 533528 228404 533580 228410
rect 533528 228346 533580 228352
rect 533344 227044 533396 227050
rect 533344 226986 533396 226992
rect 532516 223440 532568 223446
rect 532516 223382 532568 223388
rect 532056 223032 532108 223038
rect 532056 222974 532108 222980
rect 532528 222222 532556 223382
rect 532516 222216 532568 222222
rect 532516 222158 532568 222164
rect 531688 220516 531740 220522
rect 531688 220458 531740 220464
rect 531136 220380 531188 220386
rect 531136 220322 531188 220328
rect 530584 217592 530636 217598
rect 530584 217534 530636 217540
rect 530952 217592 531004 217598
rect 530952 217534 531004 217540
rect 526364 217246 526806 217274
rect 527560 217246 527634 217274
rect 528388 217246 528462 217274
rect 529216 217246 529290 217274
rect 530044 217246 530118 217274
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527606 216988 527634 217246
rect 528434 216988 528462 217246
rect 529262 216988 529290 217246
rect 530090 216988 530118 217246
rect 530964 217138 530992 217534
rect 531700 217274 531728 220458
rect 532528 217274 532556 222158
rect 533540 219434 533568 228346
rect 534000 221610 534028 231676
rect 534644 230042 534672 231676
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534816 229764 534868 229770
rect 534816 229706 534868 229712
rect 534828 223446 534856 229706
rect 535000 224936 535052 224942
rect 535000 224878 535052 224884
rect 534816 223440 534868 223446
rect 534816 223382 534868 223388
rect 533988 221604 534040 221610
rect 533988 221546 534040 221552
rect 534172 220108 534224 220114
rect 534172 220050 534224 220056
rect 533448 219406 533568 219434
rect 533448 217326 533476 219406
rect 533436 217320 533488 217326
rect 531700 217246 531774 217274
rect 532528 217246 532602 217274
rect 533436 217262 533488 217268
rect 534184 217274 534212 220050
rect 535012 217274 535040 224878
rect 535288 224262 535316 231676
rect 535736 227452 535788 227458
rect 535736 227394 535788 227400
rect 535276 224256 535328 224262
rect 535276 224198 535328 224204
rect 535460 223304 535512 223310
rect 535460 223246 535512 223252
rect 535472 217870 535500 223246
rect 535748 219434 535776 227394
rect 535932 225758 535960 231676
rect 536104 230444 536156 230450
rect 536104 230386 536156 230392
rect 536116 227458 536144 230386
rect 536576 229906 536604 231676
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 537220 228410 537248 231676
rect 537878 231662 538168 231690
rect 537208 228404 537260 228410
rect 537208 228346 537260 228352
rect 537484 227588 537536 227594
rect 537484 227530 537536 227536
rect 536104 227452 536156 227458
rect 536104 227394 536156 227400
rect 535920 225752 535972 225758
rect 535920 225694 535972 225700
rect 535748 219406 535960 219434
rect 535460 217864 535512 217870
rect 535460 217806 535512 217812
rect 535932 217734 535960 219406
rect 537496 218618 537524 227530
rect 538140 220114 538168 231662
rect 538508 229770 538536 231676
rect 538784 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 538312 229628 538364 229634
rect 538312 229570 538364 229576
rect 538324 226030 538352 229570
rect 538496 226160 538548 226166
rect 538496 226102 538548 226108
rect 538312 226024 538364 226030
rect 538312 225966 538364 225972
rect 538508 225842 538536 226102
rect 538324 225814 538536 225842
rect 538128 220108 538180 220114
rect 538128 220050 538180 220056
rect 538324 219434 538352 225814
rect 538784 221474 538812 231662
rect 539600 230308 539652 230314
rect 539600 230250 539652 230256
rect 539612 228682 539640 230250
rect 547144 230172 547196 230178
rect 547144 230114 547196 230120
rect 542820 228948 542872 228954
rect 542820 228890 542872 228896
rect 541624 228812 541676 228818
rect 541624 228754 541676 228760
rect 539416 228676 539468 228682
rect 539416 228618 539468 228624
rect 539600 228676 539652 228682
rect 539600 228618 539652 228624
rect 539428 228274 539456 228618
rect 539416 228268 539468 228274
rect 539416 228210 539468 228216
rect 540888 228268 540940 228274
rect 540888 228210 540940 228216
rect 539968 226296 540020 226302
rect 539968 226238 540020 226244
rect 538956 224528 539008 224534
rect 538956 224470 539008 224476
rect 538968 221474 538996 224470
rect 539980 224058 540008 226238
rect 539968 224052 540020 224058
rect 539968 223994 540020 224000
rect 538772 221468 538824 221474
rect 538772 221410 538824 221416
rect 538956 221468 539008 221474
rect 538956 221410 539008 221416
rect 538968 219434 538996 221410
rect 538232 219406 538352 219434
rect 538416 219406 538996 219434
rect 537484 218612 537536 218618
rect 537484 218554 537536 218560
rect 536656 217864 536708 217870
rect 536656 217806 536708 217812
rect 536840 217864 536892 217870
rect 536840 217806 536892 217812
rect 535920 217728 535972 217734
rect 535920 217670 535972 217676
rect 535932 217274 535960 217670
rect 530918 217110 530992 217138
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532574 216988 532602 217246
rect 533448 217138 533476 217262
rect 534184 217246 534258 217274
rect 535012 217246 535086 217274
rect 533402 217110 533476 217138
rect 533402 216988 533430 217110
rect 534230 216988 534258 217246
rect 535058 216988 535086 217246
rect 535886 217246 535960 217274
rect 535886 216988 535914 217246
rect 536668 217138 536696 217806
rect 536852 217598 536880 217806
rect 536840 217592 536892 217598
rect 536840 217534 536892 217540
rect 537496 217274 537524 218554
rect 538232 217598 538260 219406
rect 538220 217592 538272 217598
rect 538220 217534 538272 217540
rect 538416 217274 538444 219406
rect 539140 217592 539192 217598
rect 539140 217534 539192 217540
rect 537496 217246 537570 217274
rect 536668 217110 536742 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217246
rect 538370 217246 538444 217274
rect 538370 216988 538398 217246
rect 539152 217138 539180 217534
rect 539980 217274 540008 223994
rect 540900 222057 540928 228210
rect 540886 222048 540942 222057
rect 540886 221983 540942 221992
rect 540900 217274 540928 221983
rect 539980 217246 540054 217274
rect 539152 217110 539226 217138
rect 539198 216988 539226 217110
rect 540026 216988 540054 217246
rect 540854 217246 540928 217274
rect 541636 217274 541664 228754
rect 542832 224534 542860 228890
rect 545764 225888 545816 225894
rect 545764 225830 545816 225836
rect 544384 224664 544436 224670
rect 544384 224606 544436 224612
rect 542452 224528 542504 224534
rect 542452 224470 542504 224476
rect 542820 224528 542872 224534
rect 542820 224470 542872 224476
rect 542464 217274 542492 224470
rect 543280 222896 543332 222902
rect 543280 222838 543332 222844
rect 543094 221776 543150 221785
rect 543094 221711 543150 221720
rect 543108 221474 543136 221711
rect 543096 221468 543148 221474
rect 543096 221410 543148 221416
rect 543292 221406 543320 222838
rect 543830 222048 543886 222057
rect 544198 222048 544254 222057
rect 543830 221983 543886 221992
rect 544028 222006 544198 222034
rect 543844 221746 543872 221983
rect 544028 221950 544056 222006
rect 544198 221983 544254 221992
rect 544016 221944 544068 221950
rect 544016 221886 544068 221892
rect 544200 221876 544252 221882
rect 544200 221818 544252 221824
rect 544014 221776 544070 221785
rect 543694 221740 543746 221746
rect 543694 221682 543746 221688
rect 543832 221740 543884 221746
rect 544014 221711 544070 221720
rect 543832 221682 543884 221688
rect 543280 221400 543332 221406
rect 543280 221342 543332 221348
rect 542820 218748 542872 218754
rect 542820 218690 542872 218696
rect 542832 218482 542860 218690
rect 542820 218476 542872 218482
rect 542820 218418 542872 218424
rect 543292 217274 543320 221342
rect 543706 221218 543734 221682
rect 544028 221474 544056 221711
rect 544016 221468 544068 221474
rect 544016 221410 544068 221416
rect 543832 221400 543884 221406
rect 544212 221354 544240 221818
rect 543884 221348 544240 221354
rect 543832 221342 544240 221348
rect 543844 221326 544240 221342
rect 543706 221190 543872 221218
rect 543844 220726 543872 221190
rect 543832 220720 543884 220726
rect 543832 220662 543884 220668
rect 544396 217274 544424 224606
rect 545028 220584 545080 220590
rect 545028 220526 545080 220532
rect 545040 218618 545068 220526
rect 545028 218612 545080 218618
rect 545028 218554 545080 218560
rect 541636 217246 541710 217274
rect 542464 217246 542538 217274
rect 543292 217246 543366 217274
rect 540854 216988 540882 217246
rect 541682 216988 541710 217246
rect 542510 216988 542538 217246
rect 543338 216988 543366 217246
rect 544166 217246 544424 217274
rect 544166 216988 544194 217246
rect 545040 217138 545068 218554
rect 545776 217598 545804 225830
rect 546590 222048 546646 222057
rect 546590 221983 546646 221992
rect 545764 217592 545816 217598
rect 545764 217534 545816 217540
rect 545776 217274 545804 217534
rect 545776 217246 545850 217274
rect 544994 217110 545068 217138
rect 544994 216988 545022 217110
rect 545822 216988 545850 217246
rect 546604 217138 546632 221983
rect 547156 221921 547184 230114
rect 549260 230036 549312 230042
rect 549260 229978 549312 229984
rect 548340 227180 548392 227186
rect 548340 227122 548392 227128
rect 547420 223440 547472 223446
rect 547420 223382 547472 223388
rect 547142 221912 547198 221921
rect 547142 221847 547198 221856
rect 547432 219026 547460 223382
rect 548352 220522 548380 227122
rect 549272 224806 549300 229978
rect 553308 228540 553360 228546
rect 553308 228482 553360 228488
rect 552664 227452 552716 227458
rect 552664 227394 552716 227400
rect 551560 227316 551612 227322
rect 551560 227258 551612 227264
rect 549260 224800 549312 224806
rect 549260 224742 549312 224748
rect 549996 224664 550048 224670
rect 549996 224606 550048 224612
rect 549076 220720 549128 220726
rect 549076 220662 549128 220668
rect 548340 220516 548392 220522
rect 548340 220458 548392 220464
rect 547420 219020 547472 219026
rect 547420 218962 547472 218968
rect 547432 217138 547460 218962
rect 548352 217274 548380 220458
rect 548524 218748 548576 218754
rect 548524 218690 548576 218696
rect 548536 218210 548564 218690
rect 548524 218204 548576 218210
rect 548524 218146 548576 218152
rect 548306 217246 548380 217274
rect 546604 217110 546678 217138
rect 547432 217110 547506 217138
rect 546650 216988 546678 217110
rect 547478 216988 547506 217110
rect 548306 216988 548334 217246
rect 549088 217138 549116 220662
rect 550008 217138 550036 224606
rect 550640 224392 550692 224398
rect 550640 224334 550692 224340
rect 550652 220726 550680 224334
rect 550640 220720 550692 220726
rect 550640 220662 550692 220668
rect 550824 220720 550876 220726
rect 550824 220662 550876 220668
rect 550836 217138 550864 220662
rect 551572 217274 551600 227258
rect 552676 219162 552704 227394
rect 553320 224954 553348 228482
rect 553136 224926 553348 224954
rect 553136 222194 553164 224926
rect 554056 222902 554084 249047
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244322 554544 244695
rect 554504 244316 554556 244322
rect 554504 244258 554556 244264
rect 554502 240408 554558 240417
rect 554502 240343 554558 240352
rect 554516 240174 554544 240343
rect 554504 240168 554556 240174
rect 554504 240110 554556 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 555436 228546 555464 255546
rect 556804 251252 556856 251258
rect 556804 251194 556856 251200
rect 555976 228676 556028 228682
rect 555976 228618 556028 228624
rect 555424 228540 555476 228546
rect 555424 228482 555476 228488
rect 555988 224954 556016 228618
rect 556816 227186 556844 251194
rect 558184 246356 558236 246362
rect 558184 246298 558236 246304
rect 558196 236094 558224 246298
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 559564 229900 559616 229906
rect 559564 229842 559616 229848
rect 556804 227180 556856 227186
rect 556804 227122 556856 227128
rect 557264 226024 557316 226030
rect 557264 225966 557316 225972
rect 555896 224926 556016 224954
rect 555896 224330 555924 224926
rect 557276 224806 557304 225966
rect 558184 225616 558236 225622
rect 558184 225558 558236 225564
rect 558196 224954 558224 225558
rect 557920 224926 558224 224954
rect 557080 224800 557132 224806
rect 557078 224768 557080 224777
rect 557264 224800 557316 224806
rect 557132 224768 557134 224777
rect 557264 224742 557316 224748
rect 557078 224703 557134 224712
rect 554964 224324 555016 224330
rect 554964 224266 555016 224272
rect 555884 224324 555936 224330
rect 555884 224266 555936 224272
rect 554044 222896 554096 222902
rect 554044 222838 554096 222844
rect 552938 222184 552994 222193
rect 553136 222166 553256 222194
rect 552938 222119 552994 222128
rect 552952 222018 552980 222119
rect 552940 222012 552992 222018
rect 552940 221954 552992 221960
rect 553228 220640 553256 222166
rect 553582 222184 553638 222193
rect 553638 222142 553992 222170
rect 553582 222119 553638 222128
rect 553964 222086 553992 222142
rect 553952 222080 554004 222086
rect 553952 222022 554004 222028
rect 553228 220612 553302 220640
rect 552848 220516 552900 220522
rect 553274 220504 553302 220612
rect 552848 220458 552900 220464
rect 553228 220476 553302 220504
rect 552860 220289 552888 220458
rect 552846 220280 552902 220289
rect 552846 220215 552902 220224
rect 553228 219201 553256 220476
rect 553950 220416 554006 220425
rect 553400 220380 553452 220386
rect 553950 220351 553952 220360
rect 553400 220322 553452 220328
rect 554004 220351 554006 220360
rect 553952 220322 554004 220328
rect 553214 219192 553270 219201
rect 552664 219156 552716 219162
rect 553214 219127 553270 219136
rect 552664 219098 552716 219104
rect 552676 217274 552704 219098
rect 551572 217246 551646 217274
rect 549088 217110 549162 217138
rect 549134 216988 549162 217110
rect 549962 217110 550036 217138
rect 550790 217110 550864 217138
rect 549962 216988 549990 217110
rect 550790 216988 550818 217110
rect 551618 216988 551646 217246
rect 552446 217246 552704 217274
rect 553228 217274 553256 219127
rect 553412 218210 553440 220322
rect 553584 220244 553636 220250
rect 553584 220186 553636 220192
rect 553596 218226 553624 220186
rect 553400 218204 553452 218210
rect 553596 218198 554084 218226
rect 553400 218146 553452 218152
rect 554056 217274 554084 218198
rect 554976 217274 555004 224266
rect 555700 223168 555752 223174
rect 555700 223110 555752 223116
rect 555712 217841 555740 223110
rect 556528 218204 556580 218210
rect 556528 218146 556580 218152
rect 555698 217832 555754 217841
rect 555698 217767 555754 217776
rect 553228 217246 553302 217274
rect 554056 217246 554130 217274
rect 552446 216988 552474 217246
rect 553274 216988 553302 217246
rect 554102 216988 554130 217246
rect 554930 217246 555004 217274
rect 554930 216988 554958 217246
rect 555712 217138 555740 217767
rect 556540 217138 556568 218146
rect 557276 217274 557304 224742
rect 557920 222329 557948 224926
rect 559012 223032 559064 223038
rect 559012 222974 559064 222980
rect 558184 222760 558236 222766
rect 558184 222702 558236 222708
rect 558196 222494 558224 222702
rect 558184 222488 558236 222494
rect 558184 222430 558236 222436
rect 558552 222488 558604 222494
rect 558552 222430 558604 222436
rect 557906 222320 557962 222329
rect 557906 222255 557962 222264
rect 557920 221490 557948 222255
rect 558564 221921 558592 222430
rect 558550 221912 558606 221921
rect 558550 221847 558606 221856
rect 558092 221740 558144 221746
rect 558092 221682 558144 221688
rect 558104 221626 558132 221682
rect 558104 221610 558684 221626
rect 558104 221604 558696 221610
rect 558104 221598 558644 221604
rect 558644 221546 558696 221552
rect 557920 221462 558224 221490
rect 557816 219292 557868 219298
rect 557816 219234 557868 219240
rect 557632 219020 557684 219026
rect 557632 218962 557684 218968
rect 557644 218210 557672 218962
rect 557828 218618 557856 219234
rect 558000 218884 558052 218890
rect 558000 218826 558052 218832
rect 558012 218618 558040 218826
rect 557816 218612 557868 218618
rect 557816 218554 557868 218560
rect 558000 218612 558052 218618
rect 558000 218554 558052 218560
rect 557632 218204 557684 218210
rect 557632 218146 557684 218152
rect 558196 217274 558224 221462
rect 557276 217246 557442 217274
rect 558196 217246 558270 217274
rect 555712 217110 555786 217138
rect 556540 217110 556614 217138
rect 555758 216988 555786 217110
rect 556586 216988 556614 217110
rect 557414 216988 557442 217246
rect 558242 216988 558270 217246
rect 559024 217138 559052 222974
rect 559576 222057 559604 229842
rect 560760 227044 560812 227050
rect 560760 226986 560812 226992
rect 560772 224954 560800 226986
rect 560588 224926 560800 224954
rect 559840 222488 559892 222494
rect 559840 222430 559892 222436
rect 559562 222048 559618 222057
rect 559562 221983 559618 221992
rect 559852 217274 559880 222430
rect 560588 220522 560616 224926
rect 560956 221814 560984 259422
rect 563704 256760 563756 256766
rect 563704 256702 563756 256708
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 561678 224768 561734 224777
rect 561678 224703 561734 224712
rect 560760 221808 560812 221814
rect 560760 221750 560812 221756
rect 560944 221808 560996 221814
rect 560944 221750 560996 221756
rect 560576 220516 560628 220522
rect 560576 220458 560628 220464
rect 560208 219904 560260 219910
rect 560208 219846 560260 219852
rect 560220 219201 560248 219846
rect 560206 219192 560262 219201
rect 560206 219127 560262 219136
rect 560208 218612 560260 218618
rect 560208 218554 560260 218560
rect 560220 218210 560248 218554
rect 560208 218204 560260 218210
rect 560208 218146 560260 218152
rect 559852 217246 559926 217274
rect 559024 217110 559098 217138
rect 559070 216988 559098 217110
rect 559898 216988 559926 217246
rect 560588 217138 560616 220458
rect 560772 217274 560800 221750
rect 561692 219366 561720 224703
rect 562336 224262 562364 252554
rect 563716 226302 563744 256702
rect 566464 229764 566516 229770
rect 566464 229706 566516 229712
rect 565636 228404 565688 228410
rect 565636 228346 565688 228352
rect 563704 226296 563756 226302
rect 563704 226238 563756 226244
rect 563060 225752 563112 225758
rect 563060 225694 563112 225700
rect 563072 224954 563100 225694
rect 563072 224926 564020 224954
rect 562324 224256 562376 224262
rect 562324 224198 562376 224204
rect 562140 224188 562192 224194
rect 562140 224130 562192 224136
rect 562152 223514 562180 224130
rect 562140 223508 562192 223514
rect 562140 223450 562192 223456
rect 563336 223508 563388 223514
rect 563336 223450 563388 223456
rect 563150 222320 563206 222329
rect 563150 222255 563206 222264
rect 562874 222048 562930 222057
rect 562874 221983 562930 221992
rect 562692 221808 562744 221814
rect 562690 221776 562692 221785
rect 562744 221776 562746 221785
rect 562888 221746 562916 221983
rect 563164 221746 563192 222255
rect 562690 221711 562746 221720
rect 562876 221740 562928 221746
rect 562876 221682 562928 221688
rect 563014 221740 563066 221746
rect 563014 221682 563066 221688
rect 563152 221740 563204 221746
rect 563152 221682 563204 221688
rect 563026 221626 563054 221682
rect 563026 221598 563192 221626
rect 563164 220697 563192 221598
rect 563150 220688 563206 220697
rect 563150 220623 563206 220632
rect 562876 220516 562928 220522
rect 562876 220458 562928 220464
rect 562888 220017 562916 220458
rect 563348 220425 563376 223450
rect 563334 220416 563390 220425
rect 563334 220351 563390 220360
rect 562874 220008 562930 220017
rect 562874 219943 562930 219952
rect 561680 219360 561732 219366
rect 561680 219302 561732 219308
rect 562324 219360 562376 219366
rect 562324 219302 562376 219308
rect 562140 218204 562192 218210
rect 562140 218146 562192 218152
rect 560772 217246 561582 217274
rect 560588 217110 560754 217138
rect 560726 216988 560754 217110
rect 561554 216988 561582 217246
rect 562152 217190 562180 218146
rect 562140 217184 562192 217190
rect 562140 217126 562192 217132
rect 562336 217138 562364 219302
rect 563060 218204 563112 218210
rect 563060 218146 563112 218152
rect 562690 217832 562746 217841
rect 562690 217767 562746 217776
rect 562874 217832 562930 217841
rect 562874 217767 562930 217776
rect 562704 217190 562732 217767
rect 562508 217184 562560 217190
rect 562336 217110 562410 217138
rect 562508 217126 562560 217132
rect 562692 217184 562744 217190
rect 562692 217126 562744 217132
rect 562382 216988 562410 217110
rect 562520 217036 562548 217126
rect 562888 217036 562916 217767
rect 563072 217190 563100 218146
rect 563348 217274 563376 220351
rect 563520 220244 563572 220250
rect 563520 220186 563572 220192
rect 563532 220017 563560 220186
rect 563518 220008 563574 220017
rect 563518 219943 563574 219952
rect 563520 218000 563572 218006
rect 563520 217942 563572 217948
rect 563532 217841 563560 217942
rect 563518 217832 563574 217841
rect 563518 217767 563574 217776
rect 563210 217246 563376 217274
rect 563992 217274 564020 224926
rect 564806 220688 564862 220697
rect 564806 220623 564862 220632
rect 564820 220017 564848 220623
rect 565648 220425 565676 228346
rect 566476 224954 566504 229706
rect 568120 226296 568172 226302
rect 568120 226238 568172 226244
rect 566476 224926 566688 224954
rect 565634 220416 565690 220425
rect 566660 220386 566688 224926
rect 565634 220351 565690 220360
rect 566464 220380 566516 220386
rect 564806 220008 564862 220017
rect 564806 219943 564862 219952
rect 563992 217246 564066 217274
rect 563060 217184 563112 217190
rect 563060 217126 563112 217132
rect 562520 217008 562916 217036
rect 563210 216988 563238 217246
rect 564038 216988 564066 217246
rect 564820 217138 564848 219943
rect 565648 217274 565676 220351
rect 566464 220322 566516 220328
rect 566648 220380 566700 220386
rect 566648 220322 566700 220328
rect 567292 220380 567344 220386
rect 567292 220322 567344 220328
rect 565648 217246 565722 217274
rect 564820 217110 564894 217138
rect 564866 216988 564894 217110
rect 565694 216988 565722 217246
rect 566476 217138 566504 220322
rect 566752 219422 567148 219450
rect 566752 218890 566780 219422
rect 567120 219366 567148 219422
rect 566924 219360 566976 219366
rect 566924 219302 566976 219308
rect 567108 219360 567160 219366
rect 567108 219302 567160 219308
rect 566740 218884 566792 218890
rect 566740 218826 566792 218832
rect 566936 217841 566964 219302
rect 567106 219192 567162 219201
rect 567106 219127 567162 219136
rect 567120 219026 567148 219127
rect 567108 219020 567160 219026
rect 567108 218962 567160 218968
rect 566922 217832 566978 217841
rect 566922 217767 566978 217776
rect 567304 217138 567332 220322
rect 567476 219156 567528 219162
rect 567476 219098 567528 219104
rect 567488 218618 567516 219098
rect 567660 219020 567712 219026
rect 567660 218962 567712 218968
rect 567476 218612 567528 218618
rect 567476 218554 567528 218560
rect 567672 218482 567700 218962
rect 567660 218476 567712 218482
rect 567660 218418 567712 218424
rect 568132 217274 568160 226238
rect 568592 220386 568620 260850
rect 570616 234598 570644 261462
rect 647252 246362 647280 278038
rect 647240 246356 647292 246362
rect 647240 246298 647292 246304
rect 596824 245676 596876 245682
rect 596824 245618 596876 245624
rect 573364 244316 573416 244322
rect 573364 244258 573416 244264
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 571340 228540 571392 228546
rect 571340 228482 571392 228488
rect 570604 227180 570656 227186
rect 570604 227122 570656 227128
rect 568946 221776 569002 221785
rect 568946 221711 569002 221720
rect 568396 220380 568448 220386
rect 568396 220322 568448 220328
rect 568580 220380 568632 220386
rect 568580 220322 568632 220328
rect 568408 219314 568436 220322
rect 568408 219286 568528 219314
rect 568302 219192 568358 219201
rect 568302 219127 568358 219136
rect 568316 218890 568344 219127
rect 568304 218884 568356 218890
rect 568304 218826 568356 218832
rect 568500 218754 568528 219286
rect 568488 218748 568540 218754
rect 568488 218690 568540 218696
rect 568132 217246 568206 217274
rect 566476 217110 566550 217138
rect 567304 217110 567378 217138
rect 566522 216988 566550 217110
rect 567350 216988 567378 217110
rect 568178 216988 568206 217246
rect 568960 217138 568988 221711
rect 569958 220416 570014 220425
rect 569776 220380 569828 220386
rect 569958 220351 569960 220360
rect 569776 220322 569828 220328
rect 570012 220351 570014 220360
rect 569960 220322 570012 220328
rect 569788 217138 569816 220322
rect 570616 217274 570644 227122
rect 571352 224954 571380 228482
rect 571352 224926 571748 224954
rect 571432 224256 571484 224262
rect 571432 224198 571484 224204
rect 571444 217274 571472 224198
rect 571720 217274 571748 224926
rect 572994 220552 573050 220561
rect 572456 220510 572994 220538
rect 572456 220386 572484 220510
rect 572994 220487 573050 220496
rect 572626 220416 572682 220425
rect 572444 220380 572496 220386
rect 572626 220351 572682 220360
rect 572810 220416 572866 220425
rect 572810 220351 572866 220360
rect 572996 220380 573048 220386
rect 572444 220322 572496 220328
rect 572640 220250 572668 220351
rect 572824 220250 572852 220351
rect 572996 220322 573048 220328
rect 572628 220244 572680 220250
rect 572628 220186 572680 220192
rect 572812 220244 572864 220250
rect 572812 220186 572864 220192
rect 573008 220153 573036 220322
rect 573376 220289 573404 244258
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 573362 220280 573418 220289
rect 573362 220215 573418 220224
rect 572994 220144 573050 220153
rect 572088 220102 572760 220130
rect 571892 219360 571944 219366
rect 571892 219302 571944 219308
rect 571904 218362 571932 219302
rect 572088 218890 572116 220102
rect 572534 220008 572590 220017
rect 572534 219943 572590 219952
rect 572260 219360 572312 219366
rect 572260 219302 572312 219308
rect 572076 218884 572128 218890
rect 572076 218826 572128 218832
rect 572272 218754 572300 219302
rect 572548 218890 572576 219943
rect 572732 218890 572760 220102
rect 572994 220079 573050 220088
rect 574284 219156 574336 219162
rect 574284 219098 574336 219104
rect 572536 218884 572588 218890
rect 572536 218826 572588 218832
rect 572720 218884 572772 218890
rect 572720 218826 572772 218832
rect 572260 218748 572312 218754
rect 572260 218690 572312 218696
rect 571904 218334 572484 218362
rect 572456 218210 572484 218334
rect 572444 218204 572496 218210
rect 572444 218146 572496 218152
rect 572076 218000 572128 218006
rect 572076 217942 572128 217948
rect 572088 217841 572116 217942
rect 572074 217832 572130 217841
rect 572074 217767 572130 217776
rect 574098 217832 574154 217841
rect 574098 217767 574154 217776
rect 570616 217246 570690 217274
rect 571444 217246 571518 217274
rect 571720 217246 572346 217274
rect 568960 217110 569034 217138
rect 569788 217110 569862 217138
rect 569006 216988 569034 217110
rect 569834 216988 569862 217110
rect 570662 216988 570690 217246
rect 571490 216988 571518 217246
rect 572318 216988 572346 217246
rect 574112 216918 574140 217767
rect 574100 216912 574152 216918
rect 574100 216854 574152 216860
rect 574098 216744 574154 216753
rect 574098 216679 574154 216688
rect 574112 213518 574140 216679
rect 574296 214742 574324 219098
rect 575480 219020 575532 219026
rect 575480 218962 575532 218968
rect 574468 218884 574520 218890
rect 574468 218826 574520 218832
rect 574284 214736 574336 214742
rect 574284 214678 574336 214684
rect 574480 214606 574508 218826
rect 574834 217832 574890 217841
rect 574834 217767 574890 217776
rect 574650 216744 574706 216753
rect 574650 216679 574706 216688
rect 574468 214600 574520 214606
rect 574468 214542 574520 214548
rect 574100 213512 574152 213518
rect 574100 213454 574152 213460
rect 574664 213382 574692 216679
rect 574652 213376 574704 213382
rect 574652 213318 574704 213324
rect 574848 213246 574876 217767
rect 575492 214878 575520 218962
rect 575480 214872 575532 214878
rect 575480 214814 575532 214820
rect 574836 213240 574888 213246
rect 574836 213182 574888 213188
rect 577516 99142 577544 240110
rect 596836 231130 596864 245618
rect 648632 242214 648660 278052
rect 651944 277394 651972 282095
rect 652128 277394 652156 282254
rect 651944 277366 652064 277394
rect 652128 277366 652248 277394
rect 650642 256728 650698 256737
rect 650642 256663 650698 256672
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 629944 241528 629996 241534
rect 629944 241470 629996 241476
rect 596824 231124 596876 231130
rect 596824 231066 596876 231072
rect 629956 229094 629984 241470
rect 639604 232552 639656 232558
rect 639604 232494 639656 232500
rect 633624 231124 633676 231130
rect 633624 231066 633676 231072
rect 636844 231124 636896 231130
rect 636844 231066 636896 231072
rect 629956 229066 630076 229094
rect 621020 224936 621072 224942
rect 621020 224878 621072 224884
rect 619640 223916 619692 223922
rect 619640 223858 619692 223864
rect 617064 223780 617116 223786
rect 617064 223722 617116 223728
rect 614948 223644 615000 223650
rect 614948 223586 615000 223592
rect 593972 222624 594024 222630
rect 593972 222566 594024 222572
rect 589646 220552 589702 220561
rect 589646 220487 589702 220496
rect 586334 220280 586390 220289
rect 586334 220215 586390 220224
rect 586348 220130 586376 220215
rect 586348 220114 586560 220130
rect 586348 220108 586572 220114
rect 586348 220102 586520 220108
rect 586520 220050 586572 220056
rect 586336 220040 586388 220046
rect 586334 220008 586336 220017
rect 586388 220008 586390 220017
rect 586334 219943 586390 219952
rect 589462 220008 589518 220017
rect 589462 219943 589518 219952
rect 589280 219768 589332 219774
rect 589280 219710 589332 219716
rect 589292 219230 589320 219710
rect 589476 219502 589504 219943
rect 589660 219774 589688 220487
rect 589648 219768 589700 219774
rect 589648 219710 589700 219716
rect 589464 219496 589516 219502
rect 589464 219438 589516 219444
rect 589280 219224 589332 219230
rect 589280 219166 589332 219172
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578570 211656
rect 578528 211206 578556 211647
rect 578516 211200 578568 211206
rect 578516 211142 578568 211148
rect 578896 208350 578924 213959
rect 580908 211200 580960 211206
rect 580908 211142 580960 211148
rect 579528 209840 579580 209846
rect 579526 209808 579528 209817
rect 579580 209808 579582 209817
rect 579526 209743 579582 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 580920 206922 580948 211142
rect 593984 210202 594012 222566
rect 596928 222142 597324 222170
rect 596928 222086 596956 222142
rect 596916 222080 596968 222086
rect 596916 222022 596968 222028
rect 597296 222034 597324 222142
rect 597100 222012 597152 222018
rect 597296 222006 597508 222034
rect 597100 221954 597152 221960
rect 597112 221474 597140 221954
rect 597480 221882 597508 222006
rect 605012 222012 605064 222018
rect 605012 221954 605064 221960
rect 597284 221876 597336 221882
rect 597284 221818 597336 221824
rect 597468 221876 597520 221882
rect 597468 221818 597520 221824
rect 603172 221876 603224 221882
rect 603172 221818 603224 221824
rect 597100 221468 597152 221474
rect 597100 221410 597152 221416
rect 597296 221406 597324 221818
rect 598938 221504 598994 221513
rect 598938 221439 598994 221448
rect 597284 221400 597336 221406
rect 597284 221342 597336 221348
rect 596824 219360 596876 219366
rect 596824 219302 596876 219308
rect 594798 218376 594854 218385
rect 594798 218311 594854 218320
rect 594812 216782 594840 218311
rect 595166 217560 595222 217569
rect 595166 217495 595222 217504
rect 594800 216776 594852 216782
rect 594800 216718 594852 216724
rect 594800 213512 594852 213518
rect 594800 213454 594852 213460
rect 594812 210202 594840 213454
rect 595180 210202 595208 217495
rect 596362 217288 596418 217297
rect 596362 217223 596418 217232
rect 595718 217016 595774 217025
rect 595718 216951 595774 216960
rect 595732 210202 595760 216951
rect 596376 210202 596404 217223
rect 596836 210202 596864 219302
rect 597928 219224 597980 219230
rect 597928 219166 597980 219172
rect 597560 216912 597612 216918
rect 597560 216854 597612 216860
rect 597572 210202 597600 216854
rect 597940 210202 597968 219166
rect 598756 218612 598808 218618
rect 598756 218554 598808 218560
rect 598572 217864 598624 217870
rect 598572 217806 598624 217812
rect 598204 217728 598256 217734
rect 598204 217670 598256 217676
rect 598216 216918 598244 217670
rect 598584 217326 598612 217806
rect 598768 217326 598796 218554
rect 598572 217320 598624 217326
rect 598572 217262 598624 217268
rect 598756 217320 598808 217326
rect 598756 217262 598808 217268
rect 598952 217274 598980 221439
rect 601700 221264 601752 221270
rect 601700 221206 601752 221212
rect 600596 221128 600648 221134
rect 600596 221070 600648 221076
rect 600320 220856 600372 220862
rect 600320 220798 600372 220804
rect 600136 217592 600188 217598
rect 600136 217534 600188 217540
rect 600148 217326 600176 217534
rect 600136 217320 600188 217326
rect 598952 217246 599532 217274
rect 600136 217262 600188 217268
rect 599124 217184 599176 217190
rect 599124 217126 599176 217132
rect 598204 216912 598256 216918
rect 598204 216854 598256 216860
rect 598478 215928 598534 215937
rect 598478 215863 598534 215872
rect 598492 210202 598520 215863
rect 599136 210202 599164 217126
rect 599504 210202 599532 217246
rect 600332 210202 600360 220798
rect 600608 210202 600636 221070
rect 601332 220992 601384 220998
rect 601332 220934 601384 220940
rect 601148 220516 601200 220522
rect 601148 220458 601200 220464
rect 601160 219858 601188 220458
rect 600792 219830 601188 219858
rect 600792 219774 600820 219830
rect 600780 219768 600832 219774
rect 600780 219710 600832 219716
rect 600964 219768 601016 219774
rect 600964 219710 601016 219716
rect 600976 219502 601004 219710
rect 600964 219496 601016 219502
rect 600964 219438 601016 219444
rect 601344 219434 601372 220934
rect 601516 220788 601568 220794
rect 601516 220730 601568 220736
rect 601528 219502 601556 220730
rect 601516 219496 601568 219502
rect 601516 219438 601568 219444
rect 601160 219406 601372 219434
rect 600778 217152 600834 217161
rect 600778 217087 600834 217096
rect 600792 216918 600820 217087
rect 600780 216912 600832 216918
rect 600780 216854 600832 216860
rect 601160 210202 601188 219406
rect 601516 217728 601568 217734
rect 601516 217670 601568 217676
rect 601528 217462 601556 217670
rect 601516 217456 601568 217462
rect 601516 217398 601568 217404
rect 601332 217184 601384 217190
rect 601516 217184 601568 217190
rect 601332 217126 601384 217132
rect 601514 217152 601516 217161
rect 601568 217152 601570 217161
rect 601344 216782 601372 217126
rect 601514 217087 601570 217096
rect 601332 216776 601384 216782
rect 601332 216718 601384 216724
rect 601712 210202 601740 221206
rect 601884 218748 601936 218754
rect 601884 218690 601936 218696
rect 601896 217462 601924 218690
rect 602344 217728 602396 217734
rect 602344 217670 602396 217676
rect 601884 217456 601936 217462
rect 601884 217398 601936 217404
rect 602356 210202 602384 217670
rect 603184 210202 603212 221818
rect 603354 218648 603410 218657
rect 603354 218583 603410 218592
rect 603368 217870 603396 218583
rect 604460 218476 604512 218482
rect 604460 218418 604512 218424
rect 603356 217864 603408 217870
rect 603356 217806 603408 217812
rect 604472 217734 604500 218418
rect 604000 217728 604052 217734
rect 604000 217670 604052 217676
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 603448 217592 603500 217598
rect 603448 217534 603500 217540
rect 603460 210202 603488 217534
rect 604012 210202 604040 217670
rect 604552 217184 604604 217190
rect 604552 217126 604604 217132
rect 604564 210202 604592 217126
rect 605024 210202 605052 221954
rect 609428 221740 609480 221746
rect 609428 221682 609480 221688
rect 605932 221604 605984 221610
rect 605932 221546 605984 221552
rect 605944 210202 605972 221546
rect 606116 221400 606168 221406
rect 606116 221342 606168 221348
rect 606128 210202 606156 221342
rect 607312 220652 607364 220658
rect 607312 220594 607364 220600
rect 606760 217320 606812 217326
rect 606760 217262 606812 217268
rect 606772 210202 606800 217262
rect 607324 210202 607352 220594
rect 608692 219904 608744 219910
rect 608692 219846 608744 219852
rect 607496 219496 607548 219502
rect 607496 219438 607548 219444
rect 607508 210338 607536 219438
rect 607508 210310 607812 210338
rect 607784 210202 607812 210310
rect 608704 210202 608732 219846
rect 608968 217048 609020 217054
rect 608968 216990 609020 216996
rect 608980 210202 609008 216990
rect 609440 210202 609468 221682
rect 611452 220516 611504 220522
rect 611452 220458 611504 220464
rect 610072 220380 610124 220386
rect 610072 220322 610124 220328
rect 609888 218340 609940 218346
rect 609888 218282 609940 218288
rect 609900 217054 609928 218282
rect 609888 217048 609940 217054
rect 609888 216990 609940 216996
rect 610084 214470 610112 220322
rect 610256 220244 610308 220250
rect 610256 220186 610308 220192
rect 610072 214464 610124 214470
rect 610072 214406 610124 214412
rect 610268 210202 610296 220186
rect 610624 214464 610676 214470
rect 610624 214406 610676 214412
rect 610636 210202 610664 214406
rect 611464 210202 611492 220458
rect 611634 219464 611690 219473
rect 611634 219399 611690 219408
rect 611648 210202 611676 219399
rect 614488 218204 614540 218210
rect 614488 218146 614540 218152
rect 613384 217864 613436 217870
rect 613384 217806 613436 217812
rect 612280 216912 612332 216918
rect 612280 216854 612332 216860
rect 612292 210202 612320 216854
rect 612832 213376 612884 213382
rect 612832 213318 612884 213324
rect 612844 210202 612872 213318
rect 613396 210202 613424 217806
rect 614120 217048 614172 217054
rect 614120 216990 614172 216996
rect 614132 210202 614160 216990
rect 614500 210202 614528 218146
rect 614960 210202 614988 223586
rect 615684 218068 615736 218074
rect 615684 218010 615736 218016
rect 615696 210202 615724 218010
rect 616880 217728 616932 217734
rect 616880 217670 616932 217676
rect 616696 214736 616748 214742
rect 616696 214678 616748 214684
rect 616708 214470 616736 214678
rect 616696 214464 616748 214470
rect 616696 214406 616748 214412
rect 616144 213240 616196 213246
rect 616144 213182 616196 213188
rect 616156 210202 616184 213182
rect 616892 210202 616920 217670
rect 617076 214742 617104 223722
rect 618258 221232 618314 221241
rect 618258 221167 618314 221176
rect 617246 219736 617302 219745
rect 617246 219671 617302 219680
rect 617064 214736 617116 214742
rect 617064 214678 617116 214684
rect 617260 210202 617288 219671
rect 617800 214736 617852 214742
rect 617800 214678 617852 214684
rect 617812 210202 617840 214678
rect 618272 210202 618300 221167
rect 618902 215384 618958 215393
rect 618902 215319 618958 215328
rect 618916 210202 618944 215319
rect 619652 210202 619680 223858
rect 620284 222760 620336 222766
rect 620284 222702 620336 222708
rect 620296 222494 620324 222702
rect 620284 222488 620336 222494
rect 620284 222430 620336 222436
rect 620468 219904 620520 219910
rect 620468 219846 620520 219852
rect 619916 219632 619968 219638
rect 619916 219574 619968 219580
rect 619928 210202 619956 219574
rect 620480 210202 620508 219846
rect 621032 214742 621060 224878
rect 626540 224800 626592 224806
rect 626540 224742 626592 224748
rect 625252 224664 625304 224670
rect 625252 224606 625304 224612
rect 623228 224528 623280 224534
rect 623228 224470 623280 224476
rect 622584 224052 622636 224058
rect 622584 223994 622636 224000
rect 621204 222216 621256 222222
rect 621204 222158 621256 222164
rect 621020 214736 621072 214742
rect 621020 214678 621072 214684
rect 621216 210202 621244 222158
rect 622400 214872 622452 214878
rect 622400 214814 622452 214820
rect 621664 214736 621716 214742
rect 621664 214678 621716 214684
rect 621676 210202 621704 214678
rect 622412 210202 622440 214814
rect 622596 210338 622624 223994
rect 622596 210310 622716 210338
rect 622688 210202 622716 210310
rect 623240 210202 623268 224470
rect 623872 216776 623924 216782
rect 623872 216718 623924 216724
rect 623884 210202 623912 216718
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 624436 210202 624464 214406
rect 625264 210202 625292 224606
rect 625988 224392 626040 224398
rect 625988 224334 626040 224340
rect 625528 214600 625580 214606
rect 625528 214542 625580 214548
rect 625540 210202 625568 214542
rect 626000 210202 626028 224334
rect 626356 218884 626408 218890
rect 626356 218826 626408 218832
rect 626368 214334 626396 218826
rect 626356 214328 626408 214334
rect 626356 214270 626408 214276
rect 626552 210202 626580 224742
rect 627092 222624 627144 222630
rect 627092 222566 627144 222572
rect 627104 210202 627132 222566
rect 629852 222352 629904 222358
rect 629852 222294 629904 222300
rect 627458 218104 627514 218113
rect 627458 218039 627514 218048
rect 627472 213994 627500 218039
rect 628288 217456 628340 217462
rect 628288 217398 628340 217404
rect 627918 216200 627974 216209
rect 627918 216135 627974 216144
rect 627460 213988 627512 213994
rect 627460 213930 627512 213936
rect 627932 210202 627960 216135
rect 628300 210202 628328 217398
rect 628840 214328 628892 214334
rect 628840 214270 628892 214276
rect 628852 210202 628880 214270
rect 629392 213988 629444 213994
rect 629392 213930 629444 213936
rect 629404 210202 629432 213930
rect 629864 210202 629892 222294
rect 630048 214742 630076 229066
rect 632704 222896 632756 222902
rect 632704 222838 632756 222844
rect 630680 222488 630732 222494
rect 630680 222430 630732 222436
rect 630036 214736 630088 214742
rect 630036 214678 630088 214684
rect 630692 212430 630720 222430
rect 631322 220960 631378 220969
rect 631322 220895 631378 220904
rect 631138 218648 631194 218657
rect 631138 218583 631194 218592
rect 630680 212424 630732 212430
rect 630680 212366 630732 212372
rect 631152 210202 631180 218583
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599136 210174 599380 210202
rect 599504 210174 599932 210202
rect 600332 210174 600484 210202
rect 600608 210174 601036 210202
rect 601160 210174 601588 210202
rect 601712 210174 602140 210202
rect 602356 210174 602692 210202
rect 603184 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604564 210174 604900 210202
rect 605024 210174 605452 210202
rect 605944 210174 606004 210202
rect 606128 210174 606556 210202
rect 606772 210174 607108 210202
rect 607324 210174 607660 210202
rect 607784 210174 608212 210202
rect 608704 210174 608764 210202
rect 608980 210174 609316 210202
rect 609440 210174 609868 210202
rect 610268 210174 610420 210202
rect 610636 210174 610972 210202
rect 611464 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 614960 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 616892 210174 617044 210202
rect 617260 210174 617596 210202
rect 617812 210174 618148 210202
rect 618272 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 619928 210174 620356 210202
rect 620480 210174 620908 210202
rect 621216 210174 621460 210202
rect 621676 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623240 210174 623668 210202
rect 623884 210174 624220 210202
rect 624436 210174 624772 210202
rect 625264 210174 625324 210202
rect 625540 210174 625876 210202
rect 626000 210174 626428 210202
rect 626552 210174 626980 210202
rect 627104 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630844 210174 631180 210202
rect 631336 210202 631364 220895
rect 632716 212566 632744 222838
rect 633440 220108 633492 220114
rect 633440 220050 633492 220056
rect 633452 219434 633480 220050
rect 633452 219406 633572 219434
rect 632888 214736 632940 214742
rect 632888 214678 632940 214684
rect 632704 212560 632756 212566
rect 632704 212502 632756 212508
rect 631600 212424 631652 212430
rect 631600 212366 631652 212372
rect 631612 210202 631640 212366
rect 632900 210202 632928 214678
rect 633544 212534 633572 219406
rect 633452 212506 633572 212534
rect 633452 211070 633480 212506
rect 633440 211064 633492 211070
rect 633440 211006 633492 211012
rect 633636 210746 633664 231066
rect 634360 212560 634412 212566
rect 634360 212502 634412 212508
rect 633808 211064 633860 211070
rect 633808 211006 633860 211012
rect 633636 210718 633756 210746
rect 633728 210202 633756 210718
rect 631336 210174 631396 210202
rect 631612 210174 631948 210202
rect 632900 210174 633052 210202
rect 633604 210174 633756 210202
rect 633820 210202 633848 211006
rect 634372 210202 634400 212502
rect 636856 210202 636884 231066
rect 639616 229094 639644 232494
rect 650656 231130 650684 256663
rect 650644 231124 650696 231130
rect 650644 231066 650696 231072
rect 639616 229066 639828 229094
rect 639800 210338 639828 229066
rect 651288 224256 651340 224262
rect 651288 224198 651340 224204
rect 650642 222864 650698 222873
rect 650642 222799 650698 222808
rect 649906 221504 649962 221513
rect 649906 221439 649962 221448
rect 644754 220416 644810 220425
rect 644754 220351 644810 220360
rect 642180 217320 642232 217326
rect 642180 217262 642232 217268
rect 638972 210310 639828 210338
rect 638972 210202 639000 210310
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210186 635596 210202
rect 636580 210186 636916 210202
rect 635260 210180 635608 210186
rect 635260 210174 635556 210180
rect 635556 210122 635608 210128
rect 636568 210180 636916 210186
rect 636620 210174 636916 210180
rect 638572 210174 639000 210202
rect 639800 210202 639828 210310
rect 642192 210202 642220 217262
rect 644572 214736 644624 214742
rect 644572 214678 644624 214684
rect 643836 213240 643888 213246
rect 643836 213182 643888 213188
rect 643848 210202 643876 213182
rect 639800 210174 640228 210202
rect 641884 210174 642220 210202
rect 643540 210174 643876 210202
rect 644584 210202 644612 214678
rect 644768 210202 644796 220351
rect 648526 218648 648582 218657
rect 648526 218583 648582 218592
rect 646596 218068 646648 218074
rect 646596 218010 646648 218016
rect 646608 210202 646636 218010
rect 648252 216640 648304 216646
rect 648252 216582 648304 216588
rect 647148 213512 647200 213518
rect 647148 213454 647200 213460
rect 647160 210202 647188 213454
rect 648264 210202 648292 216582
rect 648540 210202 648568 218583
rect 649724 214872 649776 214878
rect 649724 214814 649776 214820
rect 649736 210202 649764 214814
rect 649920 213518 649948 221439
rect 649908 213512 649960 213518
rect 649908 213454 649960 213460
rect 650656 213246 650684 222799
rect 651104 213376 651156 213382
rect 651104 213318 651156 213324
rect 650644 213240 650696 213246
rect 650644 213182 650696 213188
rect 650460 212764 650512 212770
rect 650460 212706 650512 212712
rect 650472 210202 650500 212706
rect 644584 210174 644644 210202
rect 644768 210174 645196 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647956 210174 648292 210202
rect 648508 210174 648568 210202
rect 649612 210174 649764 210202
rect 650164 210174 650500 210202
rect 651116 210202 651144 213318
rect 651300 212770 651328 224198
rect 651470 221776 651526 221785
rect 651470 221711 651526 221720
rect 651288 212764 651340 212770
rect 651288 212706 651340 212712
rect 651484 210202 651512 221711
rect 651116 210174 651268 210202
rect 651484 210174 651820 210202
rect 636568 210122 636620 210128
rect 582288 209840 582340 209846
rect 582288 209782 582340 209788
rect 581644 208616 581696 208622
rect 581644 208558 581696 208564
rect 580908 206916 580960 206922
rect 580908 206858 580960 206864
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579988 167068 580040 167074
rect 579988 167010 580040 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 165232 579396 165238
rect 579344 165174 579396 165180
rect 578240 163668 578292 163674
rect 578240 163610 578292 163616
rect 578252 159905 578280 163610
rect 579356 162761 579384 165174
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 580000 163674 580028 167010
rect 579988 163668 580040 163674
rect 579988 163610 580040 163616
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579342 162752 579398 162761
rect 578424 162716 578476 162722
rect 579342 162687 579398 162696
rect 578424 162658 578476 162664
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154698 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154692 578384 154698
rect 578332 154634 578384 154640
rect 580540 154692 580592 154698
rect 580540 154634 580592 154640
rect 578344 154057 578372 154634
rect 578330 154048 578386 154057
rect 578330 153983 578386 153992
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580264 151836 580316 151842
rect 580264 151778 580316 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 578884 146328 578936 146334
rect 578884 146270 578936 146276
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578896 136649 578924 146270
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580276 140758 580304 151778
rect 580448 140820 580500 140826
rect 580448 140762 580500 140768
rect 580264 140752 580316 140758
rect 580264 140694 580316 140700
rect 579528 138712 579580 138718
rect 579528 138654 579580 138660
rect 579068 137352 579120 137358
rect 579068 137294 579120 137300
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579080 132297 579108 137294
rect 579540 134473 579568 138654
rect 580264 134564 580316 134570
rect 580264 134506 580316 134512
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131164 578936 131170
rect 578884 131106 578936 131112
rect 578896 129713 578924 131106
rect 578882 129704 578938 129713
rect 578882 129639 578938 129648
rect 579528 129056 579580 129062
rect 579528 128998 579580 129004
rect 579540 127945 579568 128998
rect 579526 127936 579582 127945
rect 579526 127871 579582 127880
rect 578332 125656 578384 125662
rect 578332 125598 578384 125604
rect 578344 125361 578372 125598
rect 578330 125352 578386 125361
rect 578330 125287 578386 125296
rect 579068 124908 579120 124914
rect 579068 124850 579120 124856
rect 578700 124160 578752 124166
rect 578700 124102 578752 124108
rect 578712 123593 578740 124102
rect 578698 123584 578754 123593
rect 578698 123519 578754 123528
rect 578884 122188 578936 122194
rect 578884 122130 578936 122136
rect 578896 121417 578924 122130
rect 578882 121408 578938 121417
rect 578882 121343 578938 121352
rect 578516 118584 578568 118590
rect 578516 118526 578568 118532
rect 578528 118425 578556 118526
rect 578514 118416 578570 118425
rect 578514 118351 578570 118360
rect 578332 108996 578384 109002
rect 578332 108938 578384 108944
rect 578344 108361 578372 108938
rect 578330 108352 578386 108361
rect 578330 108287 578386 108296
rect 579080 105913 579108 124850
rect 580276 118590 580304 134506
rect 580460 125662 580488 140762
rect 580448 125656 580500 125662
rect 580448 125598 580500 125604
rect 580632 122052 580684 122058
rect 580632 121994 580684 122000
rect 580264 118584 580316 118590
rect 580264 118526 580316 118532
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 579528 112872 579580 112878
rect 579528 112814 579580 112820
rect 579540 112577 579568 112814
rect 579526 112568 579582 112577
rect 579526 112503 579582 112512
rect 579344 110288 579396 110294
rect 579344 110230 579396 110236
rect 579356 110129 579384 110230
rect 579342 110120 579398 110129
rect 579342 110055 579398 110064
rect 580448 109132 580500 109138
rect 580448 109074 580500 109080
rect 580264 106344 580316 106350
rect 580264 106286 580316 106292
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 579344 105664 579396 105670
rect 579344 105606 579396 105612
rect 578516 103420 578568 103426
rect 578516 103362 578568 103368
rect 578528 103193 578556 103362
rect 578514 103184 578570 103193
rect 578514 103119 578570 103128
rect 579160 102128 579212 102134
rect 579160 102070 579212 102076
rect 579172 101697 579200 102070
rect 579158 101688 579214 101697
rect 579158 101623 579214 101632
rect 578608 100020 578660 100026
rect 578608 99962 578660 99968
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578620 97481 578648 99962
rect 578606 97472 578662 97481
rect 578606 97407 578662 97416
rect 578332 95192 578384 95198
rect 578332 95134 578384 95140
rect 578344 95033 578372 95134
rect 578330 95024 578386 95033
rect 578330 94959 578386 94968
rect 579356 93854 579384 105606
rect 579528 99272 579580 99278
rect 579526 99240 579528 99249
rect 579580 99240 579582 99249
rect 579526 99175 579582 99184
rect 579356 93826 579476 93854
rect 579252 93424 579304 93430
rect 579252 93366 579304 93372
rect 579264 93129 579292 93366
rect 579250 93120 579306 93129
rect 579250 93055 579306 93064
rect 578608 91180 578660 91186
rect 578608 91122 578660 91128
rect 578620 90953 578648 91122
rect 578606 90944 578662 90953
rect 578606 90879 578662 90888
rect 579252 88324 579304 88330
rect 579252 88266 579304 88272
rect 579264 88097 579292 88266
rect 579250 88088 579306 88097
rect 579250 88023 579306 88032
rect 578332 86964 578384 86970
rect 578332 86906 578384 86912
rect 578344 86465 578372 86906
rect 578330 86456 578386 86465
rect 578330 86391 578386 86400
rect 579252 84040 579304 84046
rect 579250 84008 579252 84017
rect 579304 84008 579306 84017
rect 579250 83943 579306 83952
rect 578884 82816 578936 82822
rect 578884 82758 578936 82764
rect 578896 82249 578924 82758
rect 578882 82240 578938 82249
rect 578882 82175 578938 82184
rect 579252 82136 579304 82142
rect 579252 82078 579304 82084
rect 578240 78124 578292 78130
rect 578240 78066 578292 78072
rect 578252 77897 578280 78066
rect 578238 77888 578294 77897
rect 578238 77823 578294 77832
rect 579264 75721 579292 82078
rect 579448 80073 579476 93826
rect 579434 80064 579490 80073
rect 579434 79999 579490 80008
rect 580276 78130 580304 106286
rect 580460 86970 580488 109074
rect 580644 109002 580672 121994
rect 581656 114510 581684 208558
rect 582300 205562 582328 209782
rect 652036 209574 652064 277366
rect 652220 227050 652248 277366
rect 652404 233918 652432 291479
rect 652574 283248 652630 283257
rect 652574 283183 652630 283192
rect 652392 233912 652444 233918
rect 652392 233854 652444 233860
rect 652588 229809 652616 283183
rect 654796 232558 654824 300863
rect 656164 297084 656216 297090
rect 656164 297026 656216 297032
rect 656176 271153 656204 297026
rect 656162 271144 656218 271153
rect 656162 271079 656218 271088
rect 654784 232552 654836 232558
rect 654784 232494 654836 232500
rect 652574 229800 652630 229809
rect 652574 229735 652630 229744
rect 652208 227044 652260 227050
rect 652208 226986 652260 226992
rect 654782 226400 654838 226409
rect 654782 226335 654838 226344
rect 653402 225312 653458 225321
rect 653402 225247 653458 225256
rect 653034 220688 653090 220697
rect 653034 220623 653090 220632
rect 652850 215928 652906 215937
rect 652850 215863 652906 215872
rect 652864 210202 652892 215863
rect 653048 210202 653076 220623
rect 653416 218074 653444 225247
rect 653404 218068 653456 218074
rect 653404 218010 653456 218016
rect 654796 214742 654824 226335
rect 656162 225584 656218 225593
rect 656162 225519 656218 225528
rect 655426 218920 655482 218929
rect 655426 218855 655482 218864
rect 654784 214736 654836 214742
rect 654784 214678 654836 214684
rect 654876 214600 654928 214606
rect 654876 214542 654928 214548
rect 654888 210202 654916 214542
rect 655440 210202 655468 218855
rect 656176 216646 656204 225519
rect 657726 225040 657782 225049
rect 657726 224975 657782 224984
rect 657542 223952 657598 223961
rect 657542 223887 657598 223896
rect 656806 217288 656862 217297
rect 656806 217223 656862 217232
rect 656164 216640 656216 216646
rect 656164 216582 656216 216588
rect 656530 213208 656586 213217
rect 656530 213143 656586 213152
rect 656544 210202 656572 213143
rect 656820 210202 656848 217223
rect 657556 213382 657584 223887
rect 657740 214878 657768 224975
rect 658936 217326 658964 346423
rect 664442 311944 664498 311953
rect 664442 311879 664498 311888
rect 664456 300830 664484 311879
rect 664444 300824 664496 300830
rect 664444 300766 664496 300772
rect 662420 298172 662472 298178
rect 662420 298114 662472 298120
rect 662432 293865 662460 298114
rect 665824 295996 665876 296002
rect 665824 295938 665876 295944
rect 664444 294024 664496 294030
rect 664444 293966 664496 293972
rect 662418 293856 662474 293865
rect 662418 293791 662474 293800
rect 663064 292596 663116 292602
rect 663064 292538 663116 292544
rect 660304 289876 660356 289882
rect 660304 289818 660356 289824
rect 660316 232558 660344 289818
rect 661684 288448 661736 288454
rect 661684 288390 661736 288396
rect 661696 234666 661724 288390
rect 661684 234660 661736 234666
rect 661684 234602 661736 234608
rect 660304 232552 660356 232558
rect 660304 232494 660356 232500
rect 663076 231538 663104 292538
rect 664456 248033 664484 293966
rect 665836 268569 665864 295938
rect 668124 285728 668176 285734
rect 668124 285670 668176 285676
rect 668136 283937 668164 285670
rect 668122 283928 668178 283937
rect 668122 283863 668178 283872
rect 667204 280356 667256 280362
rect 667204 280298 667256 280304
rect 665822 268560 665878 268569
rect 665822 268495 665878 268504
rect 664442 248024 664498 248033
rect 664442 247959 664498 247968
rect 665456 231668 665508 231674
rect 665456 231610 665508 231616
rect 663064 231532 663116 231538
rect 663064 231474 663116 231480
rect 662328 231396 662380 231402
rect 662328 231338 662380 231344
rect 660948 229152 661000 229158
rect 660948 229094 661000 229100
rect 660488 227792 660540 227798
rect 660488 227734 660540 227740
rect 659106 222592 659162 222601
rect 659106 222527 659162 222536
rect 658924 217320 658976 217326
rect 658924 217262 658976 217268
rect 657728 214872 657780 214878
rect 657728 214814 657780 214820
rect 658738 214568 658794 214577
rect 658738 214503 658794 214512
rect 657544 213376 657596 213382
rect 657544 213318 657596 213324
rect 658188 212900 658240 212906
rect 658188 212842 658240 212848
rect 658200 210202 658228 212842
rect 658752 210202 658780 214503
rect 659120 212906 659148 222527
rect 659568 213648 659620 213654
rect 659568 213590 659620 213596
rect 659108 212900 659160 212906
rect 659108 212842 659160 212848
rect 659580 210202 659608 213590
rect 660500 210202 660528 227734
rect 660960 210202 660988 229094
rect 662050 217560 662106 217569
rect 662050 217495 662106 217504
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662064 210202 662092 217495
rect 662340 210202 662368 231338
rect 664996 231192 665048 231198
rect 664996 231134 665048 231140
rect 663706 229392 663762 229401
rect 663706 229327 663762 229336
rect 663524 228404 663576 228410
rect 663524 228346 663576 228352
rect 663156 213920 663208 213926
rect 663156 213862 663208 213868
rect 663168 210202 663196 213862
rect 663536 210202 663564 228346
rect 663720 213926 663748 229327
rect 664442 223816 664498 223825
rect 664442 223751 664498 223760
rect 664456 214606 664484 223751
rect 665008 219434 665036 231134
rect 665468 229158 665496 231610
rect 665822 230480 665878 230489
rect 665822 230415 665878 230424
rect 665456 229152 665508 229158
rect 665178 229120 665234 229129
rect 665456 229094 665508 229100
rect 665178 229055 665234 229064
rect 665192 227798 665220 229055
rect 665180 227792 665232 227798
rect 665180 227734 665232 227740
rect 665008 219406 665128 219434
rect 664444 214600 664496 214606
rect 664444 214542 664496 214548
rect 664812 214600 664864 214606
rect 664812 214542 664864 214548
rect 663708 213920 663760 213926
rect 663708 213862 663760 213868
rect 664260 212764 664312 212770
rect 664260 212706 664312 212712
rect 664272 210202 664300 212706
rect 664824 210202 664852 214542
rect 665100 212770 665128 219406
rect 665546 216200 665602 216209
rect 665546 216135 665602 216144
rect 665560 213654 665588 216135
rect 665836 214606 665864 230415
rect 666468 225208 666520 225214
rect 666468 225150 666520 225156
rect 666480 224262 666508 225150
rect 666468 224256 666520 224262
rect 666468 224198 666520 224204
rect 667018 221096 667074 221105
rect 667018 221031 667074 221040
rect 665824 214600 665876 214606
rect 665824 214542 665876 214548
rect 665548 213648 665600 213654
rect 665548 213590 665600 213596
rect 665088 212764 665140 212770
rect 665088 212706 665140 212712
rect 652864 210174 652924 210202
rect 653048 210174 653476 210202
rect 654580 210174 654916 210202
rect 655132 210174 655468 210202
rect 656236 210174 656572 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660528 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663564 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 632152 209568 632204 209574
rect 652024 209568 652076 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652024 209510 652076 209516
rect 632164 209494 632500 209510
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 206916 589516 206922
rect 589464 206858 589516 206864
rect 589476 206417 589504 206858
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 582288 205556 582340 205562
rect 582288 205498 582340 205504
rect 589464 205556 589516 205562
rect 589464 205498 589516 205504
rect 589476 204785 589504 205498
rect 589462 204776 589518 204785
rect 589462 204711 589518 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 667032 176497 667060 221031
rect 667018 176488 667074 176497
rect 667018 176423 667074 176432
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589646 170504 589702 170513
rect 589646 170439 589702 170448
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 582380 168428 582432 168434
rect 582380 168370 582432 168376
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 582392 165238 582420 168370
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 170439
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 582380 165232 582432 165238
rect 582380 165174 582432 165180
rect 589476 164286 589504 165543
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 582484 162722 582512 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158778 589504 159015
rect 585784 158772 585836 158778
rect 585784 158714 585836 158720
rect 589464 158772 589516 158778
rect 589464 158714 589516 158720
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 150618 585824 158714
rect 589278 157448 589334 157457
rect 587164 157412 587216 157418
rect 589278 157383 589280 157392
rect 587164 157354 587216 157360
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 585784 150612 585836 150618
rect 585784 150554 585836 150560
rect 585140 149116 585192 149122
rect 585140 149058 585192 149064
rect 585152 146334 585180 149058
rect 587176 148374 587204 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585140 146328 585192 146334
rect 585140 146270 585192 146276
rect 584772 144968 584824 144974
rect 584772 144910 584824 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 139460 583076 139466
rect 583024 139402 583076 139408
rect 581828 131300 581880 131306
rect 581828 131242 581880 131248
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 110492 581696 110498
rect 581644 110434 581696 110440
rect 580632 108996 580684 109002
rect 580632 108938 580684 108944
rect 580448 86964 580500 86970
rect 580448 86906 580500 86912
rect 581656 84046 581684 110434
rect 581840 110294 581868 131242
rect 583036 124166 583064 139402
rect 584784 137358 584812 144910
rect 585784 143608 585836 143614
rect 585784 143550 585836 143556
rect 584772 137352 584824 137358
rect 584772 137294 584824 137300
rect 584588 136672 584640 136678
rect 584588 136614 584640 136620
rect 583392 129192 583444 129198
rect 583392 129134 583444 129140
rect 583024 124160 583076 124166
rect 583024 124102 583076 124108
rect 583208 120760 583260 120766
rect 583208 120702 583260 120708
rect 583024 113212 583076 113218
rect 583024 113154 583076 113160
rect 581828 110288 581880 110294
rect 581828 110230 581880 110236
rect 582288 107704 582340 107710
rect 582288 107646 582340 107652
rect 582300 105670 582328 107646
rect 582288 105664 582340 105670
rect 582288 105606 582340 105612
rect 581644 84040 581696 84046
rect 581644 83982 581696 83988
rect 583036 82822 583064 113154
rect 583220 99278 583248 120702
rect 583404 116958 583432 129134
rect 584404 122868 584456 122874
rect 584404 122810 584456 122816
rect 583392 116952 583444 116958
rect 583392 116894 583444 116900
rect 584416 102134 584444 122810
rect 584600 122194 584628 136614
rect 585796 131170 585824 143550
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 132524 586020 132530
rect 585968 132466 586020 132472
rect 585784 131164 585836 131170
rect 585784 131106 585836 131112
rect 584588 122188 584640 122194
rect 584588 122130 584640 122136
rect 585784 116000 585836 116006
rect 585784 115942 585836 115948
rect 584588 115252 584640 115258
rect 584588 115194 584640 115200
rect 584404 102128 584456 102134
rect 584404 102070 584456 102076
rect 584404 100156 584456 100162
rect 584404 100098 584456 100104
rect 583208 99272 583260 99278
rect 583208 99214 583260 99220
rect 583024 82816 583076 82822
rect 583024 82758 583076 82764
rect 583024 79348 583076 79354
rect 583024 79290 583076 79296
rect 580264 78124 580316 78130
rect 580264 78066 580316 78072
rect 580446 77888 580502 77897
rect 580446 77823 580502 77832
rect 579250 75712 579306 75721
rect 579250 75647 579306 75656
rect 578884 75200 578936 75206
rect 578884 75142 578936 75148
rect 578516 71596 578568 71602
rect 578516 71538 578568 71544
rect 578528 71233 578556 71538
rect 578514 71224 578570 71233
rect 578514 71159 578570 71168
rect 578896 60489 578924 75142
rect 579528 73160 579580 73166
rect 579526 73128 579528 73137
rect 579580 73128 579582 73137
rect 579526 73063 579582 73072
rect 579528 66904 579580 66910
rect 579526 66872 579528 66881
rect 579580 66872 579582 66881
rect 579526 66807 579582 66816
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 579528 62076 579580 62082
rect 579528 62018 579580 62024
rect 579540 61849 579568 62018
rect 579526 61840 579582 61849
rect 579526 61775 579582 61784
rect 578882 60480 578938 60489
rect 578882 60415 578938 60424
rect 578332 60036 578384 60042
rect 578332 59978 578384 59984
rect 577504 58812 577556 58818
rect 577504 58754 577556 58760
rect 576124 58676 576176 58682
rect 576124 58618 576176 58624
rect 574928 57248 574980 57254
rect 574928 57190 574980 57196
rect 574744 56024 574796 56030
rect 574744 55966 574796 55972
rect 574468 55888 574520 55894
rect 574468 55830 574520 55836
rect 574480 54777 574508 55830
rect 574466 54768 574522 54777
rect 574466 54703 574522 54712
rect 574756 53990 574784 55966
rect 574744 53984 574796 53990
rect 574744 53926 574796 53932
rect 574940 53854 574968 57190
rect 576136 55049 576164 58618
rect 576122 55040 576178 55049
rect 576122 54975 576178 54984
rect 577516 54233 577544 58754
rect 578344 56137 578372 59978
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 578330 56128 578386 56137
rect 578330 56063 578386 56072
rect 577502 54224 577558 54233
rect 577502 54159 577558 54168
rect 580460 54126 580488 77823
rect 583036 54262 583064 79290
rect 584416 71602 584444 100098
rect 584600 95198 584628 115194
rect 584588 95192 584640 95198
rect 584588 95134 584640 95140
rect 585796 91186 585824 115942
rect 585980 112878 586008 132466
rect 587176 129062 587204 142394
rect 588556 138718 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 588544 138712 588596 138718
rect 588544 138654 588596 138660
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 134570 589504 136167
rect 590382 134600 590438 134609
rect 589464 134564 589516 134570
rect 590382 134535 590438 134544
rect 589464 134506 589516 134512
rect 589462 132968 589518 132977
rect 589462 132903 589518 132912
rect 589476 132530 589504 132903
rect 589464 132524 589516 132530
rect 589464 132466 589516 132472
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 588726 129704 588782 129713
rect 588726 129639 588782 129648
rect 587164 129056 587216 129062
rect 587164 128998 587216 129004
rect 587808 127016 587860 127022
rect 587808 126958 587860 126964
rect 587820 124914 587848 126958
rect 587808 124908 587860 124914
rect 587808 124850 587860 124856
rect 587348 121508 587400 121514
rect 587348 121450 587400 121456
rect 585968 112872 586020 112878
rect 585968 112814 586020 112820
rect 586152 112464 586204 112470
rect 586152 112406 586204 112412
rect 586164 93430 586192 112406
rect 587164 104916 587216 104922
rect 587164 104858 587216 104864
rect 586152 93424 586204 93430
rect 586152 93366 586204 93372
rect 585784 91180 585836 91186
rect 585784 91122 585836 91128
rect 587176 82142 587204 104858
rect 587360 100026 587388 121450
rect 588542 103592 588598 103601
rect 588542 103527 588598 103536
rect 587348 100020 587400 100026
rect 587348 99962 587400 99968
rect 587164 82136 587216 82142
rect 587164 82078 587216 82084
rect 587164 76560 587216 76566
rect 587164 76502 587216 76508
rect 584404 71596 584456 71602
rect 584404 71538 584456 71544
rect 587176 62082 587204 76502
rect 588556 73166 588584 103527
rect 588740 103426 588768 129639
rect 590396 129198 590424 134535
rect 590384 129192 590436 129198
rect 590384 129134 590436 129140
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 590106 126440 590162 126449
rect 590106 126375 590162 126384
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 590120 122058 590148 126375
rect 590566 124808 590622 124817
rect 590566 124743 590622 124752
rect 590108 122052 590160 122058
rect 590108 121994 590160 122000
rect 589278 121544 589334 121553
rect 589278 121479 589280 121488
rect 589332 121479 589334 121488
rect 589280 121450 589332 121456
rect 590580 120766 590608 124743
rect 590568 120760 590620 120766
rect 590568 120702 590620 120708
rect 589646 119912 589702 119921
rect 589646 119847 589702 119856
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589660 115258 589688 119847
rect 590106 118280 590162 118289
rect 590106 118215 590162 118224
rect 589648 115252 589700 115258
rect 589648 115194 589700 115200
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 590120 112470 590148 118215
rect 667216 116113 667244 280298
rect 667388 280220 667440 280226
rect 667388 280162 667440 280168
rect 667400 134609 667428 280162
rect 668768 237040 668820 237046
rect 668768 236982 668820 236988
rect 668216 235136 668268 235142
rect 668216 235078 668268 235084
rect 668032 224664 668084 224670
rect 668032 224606 668084 224612
rect 667848 224256 667900 224262
rect 667848 224198 667900 224204
rect 667860 220697 667888 224198
rect 668044 221785 668072 224606
rect 668030 221776 668086 221785
rect 668030 221711 668086 221720
rect 667846 220688 667902 220697
rect 667846 220623 667902 220632
rect 668030 219736 668086 219745
rect 668030 219671 668086 219680
rect 667754 219464 667810 219473
rect 667754 219399 667810 219408
rect 667572 209092 667624 209098
rect 667572 209034 667624 209040
rect 667386 134600 667442 134609
rect 667386 134535 667442 134544
rect 667584 133385 667612 209034
rect 667768 175001 667796 219399
rect 668044 213217 668072 219671
rect 668030 213208 668086 213217
rect 668030 213143 668086 213152
rect 668030 207632 668086 207641
rect 668030 207567 668086 207576
rect 668044 204105 668072 207567
rect 668030 204096 668086 204105
rect 668030 204031 668086 204040
rect 668044 200114 668072 204031
rect 667952 200086 668072 200114
rect 667952 199209 667980 200086
rect 667938 199200 667994 199209
rect 667938 199135 667994 199144
rect 667938 194168 667994 194177
rect 667938 194103 667994 194112
rect 667952 189689 667980 194103
rect 667938 189680 667994 189689
rect 667938 189615 667994 189624
rect 668030 184376 668086 184385
rect 668030 184311 668086 184320
rect 668044 179489 668072 184311
rect 668030 179480 668086 179489
rect 668030 179415 668086 179424
rect 667754 174992 667810 175001
rect 667754 174927 667810 174936
rect 667570 133376 667626 133385
rect 667570 133311 667626 133320
rect 668044 125361 668072 179415
rect 668228 173097 668256 235078
rect 668400 234864 668452 234870
rect 668400 234806 668452 234812
rect 668214 173088 668270 173097
rect 668214 173023 668270 173032
rect 668412 169697 668440 234806
rect 668584 227180 668636 227186
rect 668584 227122 668636 227128
rect 668596 219434 668624 227122
rect 668596 219406 668716 219434
rect 668398 169688 668454 169697
rect 668398 169623 668454 169632
rect 668216 165232 668268 165238
rect 668216 165174 668268 165180
rect 668228 164937 668256 165174
rect 668214 164928 668270 164937
rect 668214 164863 668270 164872
rect 668216 163328 668268 163334
rect 668214 163296 668216 163305
rect 668268 163296 668270 163305
rect 668214 163231 668270 163240
rect 668688 161474 668716 219406
rect 668596 161446 668716 161474
rect 668216 160064 668268 160070
rect 668214 160032 668216 160041
rect 668268 160032 668270 160041
rect 668214 159967 668270 159976
rect 668596 158409 668624 161446
rect 668582 158400 668638 158409
rect 668582 158335 668638 158344
rect 668308 155168 668360 155174
rect 668306 155136 668308 155145
rect 668360 155136 668362 155145
rect 668306 155071 668362 155080
rect 668216 148776 668268 148782
rect 668216 148718 668268 148724
rect 668228 148617 668256 148718
rect 668214 148608 668270 148617
rect 668214 148543 668270 148552
rect 668216 136264 668268 136270
rect 668216 136206 668268 136212
rect 668228 135561 668256 136206
rect 668214 135552 668270 135561
rect 668214 135487 668270 135496
rect 668780 130665 668808 236982
rect 668952 227792 669004 227798
rect 668952 227734 669004 227740
rect 668964 224210 668992 227734
rect 668872 224182 668992 224210
rect 668872 219434 668900 224182
rect 669044 224052 669096 224058
rect 669044 223994 669096 224000
rect 669056 223825 669084 223994
rect 669042 223816 669098 223825
rect 669042 223751 669098 223760
rect 669044 223168 669096 223174
rect 669044 223110 669096 223116
rect 669056 222601 669084 223110
rect 669042 222592 669098 222601
rect 669042 222527 669098 222536
rect 668872 219406 668992 219434
rect 668964 138825 668992 219406
rect 669240 143721 669268 393479
rect 670606 392320 670662 392329
rect 670606 392255 670662 392264
rect 669962 345672 670018 345681
rect 669962 345607 670018 345616
rect 669596 235340 669648 235346
rect 669596 235282 669648 235288
rect 669412 234524 669464 234530
rect 669412 234466 669464 234472
rect 669424 174729 669452 234466
rect 669410 174720 669466 174729
rect 669410 174655 669466 174664
rect 669410 172000 669466 172009
rect 669410 171935 669466 171944
rect 669424 149025 669452 171935
rect 669608 165238 669636 235282
rect 669778 234288 669834 234297
rect 669778 234223 669834 234232
rect 669596 165232 669648 165238
rect 669596 165174 669648 165180
rect 669792 163334 669820 234223
rect 669780 163328 669832 163334
rect 669780 163270 669832 163276
rect 669410 149016 669466 149025
rect 669410 148951 669466 148960
rect 669226 143712 669282 143721
rect 669226 143647 669282 143656
rect 668950 138816 669006 138825
rect 668950 138751 669006 138760
rect 669976 136270 670004 345607
rect 670422 261352 670478 261361
rect 670422 261287 670478 261296
rect 670238 259720 670294 259729
rect 670238 259655 670294 259664
rect 670252 245585 670280 259655
rect 670436 247217 670464 261287
rect 670422 247208 670478 247217
rect 670422 247143 670478 247152
rect 670238 245576 670294 245585
rect 670238 245511 670294 245520
rect 670148 235816 670200 235822
rect 670148 235758 670200 235764
rect 670160 148782 670188 235758
rect 670424 234660 670476 234666
rect 670424 234602 670476 234608
rect 670436 234025 670464 234602
rect 670422 234016 670478 234025
rect 670422 233951 670478 233960
rect 670332 233232 670384 233238
rect 670332 233174 670384 233180
rect 670344 160070 670372 233174
rect 670620 171057 670648 392255
rect 672000 372609 672028 397151
rect 671986 372600 672042 372609
rect 671986 372535 672042 372544
rect 672828 357513 672856 401639
rect 673182 401296 673238 401305
rect 673182 401231 673238 401240
rect 672998 394768 673054 394777
rect 672998 394703 673054 394712
rect 673012 381041 673040 394703
rect 672998 381032 673054 381041
rect 672998 380967 673054 380976
rect 672814 357504 672870 357513
rect 672814 357439 672870 357448
rect 672354 357096 672410 357105
rect 672354 357031 672410 357040
rect 672170 355464 672226 355473
rect 672170 355399 672226 355408
rect 671986 350160 672042 350169
rect 671986 350095 672042 350104
rect 672000 332353 672028 350095
rect 671986 332344 672042 332353
rect 671986 332279 672042 332288
rect 672184 310865 672212 355399
rect 672368 312497 672396 357031
rect 673196 356833 673224 401231
rect 673366 400616 673422 400625
rect 673366 400551 673422 400560
rect 673182 356824 673238 356833
rect 673182 356759 673238 356768
rect 672538 356280 672594 356289
rect 672538 356215 672594 356224
rect 672354 312488 672410 312497
rect 672354 312423 672410 312432
rect 672552 311681 672580 356215
rect 673380 355881 673408 400551
rect 673918 399800 673974 399809
rect 673918 399735 673974 399744
rect 673734 393136 673790 393145
rect 673734 393071 673790 393080
rect 673748 376689 673776 393071
rect 673734 376680 673790 376689
rect 673734 376615 673790 376624
rect 673366 355872 673422 355881
rect 673366 355807 673422 355816
rect 673932 355065 673960 399735
rect 674378 396536 674434 396545
rect 674378 396471 674434 396480
rect 674392 394618 674420 396471
rect 674576 395321 674604 403407
rect 676048 402665 676076 410479
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 676586 402928 676642 402937
rect 676586 402863 676642 402872
rect 676034 402656 676090 402665
rect 676034 402591 676090 402600
rect 674838 402248 674894 402257
rect 674838 402183 674894 402192
rect 674852 401713 674880 402183
rect 674838 401704 674894 401713
rect 674838 401639 674894 401648
rect 676600 400897 676628 402863
rect 676586 400888 676642 400897
rect 676586 400823 676642 400832
rect 674838 399392 674894 399401
rect 674838 399327 674894 399336
rect 674852 395842 674880 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675022 398168 675078 398177
rect 675022 398103 675078 398112
rect 674852 395814 674972 395842
rect 674746 395720 674802 395729
rect 674746 395655 674802 395664
rect 674562 395312 674618 395321
rect 674562 395247 674618 395256
rect 674392 394590 674512 394618
rect 674286 394496 674342 394505
rect 674286 394431 674342 394440
rect 674300 379514 674328 394431
rect 674484 393314 674512 394590
rect 674760 393314 674788 395655
rect 674944 393314 674972 395814
rect 674392 393286 674512 393314
rect 674668 393286 674788 393314
rect 674852 393286 674972 393314
rect 674392 389174 674420 393286
rect 674392 389146 674512 389174
rect 674484 382226 674512 389146
rect 674472 382220 674524 382226
rect 674472 382162 674524 382168
rect 674300 379486 674420 379514
rect 674392 378146 674420 379486
rect 674380 378140 674432 378146
rect 674380 378082 674432 378088
rect 674668 375238 674696 393286
rect 674852 385626 674880 393286
rect 674840 385620 674892 385626
rect 674840 385562 674892 385568
rect 675036 382582 675064 398103
rect 676232 395978 676260 398375
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 675312 395950 676260 395978
rect 675312 386414 675340 395950
rect 676034 394088 676090 394097
rect 676034 394023 676090 394032
rect 676048 393145 676076 394023
rect 676034 393136 676090 393145
rect 676034 393071 676090 393080
rect 681016 388521 681044 397559
rect 683026 392728 683082 392737
rect 683026 392663 683082 392672
rect 683040 389881 683068 392663
rect 683026 389872 683082 389881
rect 683026 389807 683082 389816
rect 681002 388512 681058 388521
rect 681002 388447 681058 388456
rect 675128 386386 675340 386414
rect 675128 385710 675156 386386
rect 675404 386073 675432 386275
rect 675390 386064 675446 386073
rect 675390 385999 675446 386008
rect 675312 385750 675432 385778
rect 675312 385710 675340 385750
rect 675128 385682 675340 385710
rect 675404 385696 675432 385750
rect 675300 385620 675352 385626
rect 675300 385562 675352 385568
rect 675312 384449 675340 385562
rect 675758 385384 675814 385393
rect 675758 385319 675814 385328
rect 675772 385084 675800 385319
rect 675312 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675392 382220 675444 382226
rect 675392 382162 675444 382168
rect 675404 382024 675432 382162
rect 675758 381712 675814 381721
rect 675758 381647 675814 381656
rect 675772 381412 675800 381647
rect 675390 381032 675446 381041
rect 675390 380967 675446 380976
rect 675404 380732 675432 380967
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675116 378140 675168 378146
rect 675116 378082 675168 378088
rect 675128 377754 675156 378082
rect 675128 377726 675340 377754
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675114 376680 675170 376689
rect 675114 376615 675170 376624
rect 675128 376462 675156 376615
rect 675128 376434 675340 376462
rect 675312 376394 675340 376434
rect 675404 376394 675432 376448
rect 675312 376366 675432 376394
rect 674668 375210 675418 375238
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675666 373008 675722 373017
rect 675666 372943 675722 372952
rect 675680 372776 675708 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675574 358320 675630 358329
rect 675574 358255 675630 358264
rect 673918 355056 673974 355065
rect 673918 354991 673974 355000
rect 674102 354648 674158 354657
rect 674102 354583 674158 354592
rect 673734 352608 673790 352617
rect 673734 352543 673790 352552
rect 672998 351384 673054 351393
rect 672998 351319 673054 351328
rect 672722 348528 672778 348537
rect 672722 348463 672778 348472
rect 672538 311672 672594 311681
rect 672538 311607 672594 311616
rect 672170 310856 672226 310865
rect 672170 310791 672226 310800
rect 672538 304328 672594 304337
rect 672538 304263 672594 304272
rect 671526 302288 671582 302297
rect 671526 302223 671582 302232
rect 671342 258496 671398 258505
rect 671342 258431 671398 258440
rect 670790 256456 670846 256465
rect 670790 256391 670846 256400
rect 670804 210497 670832 256391
rect 670974 250880 671030 250889
rect 670974 250815 671030 250824
rect 670988 248033 671016 250815
rect 670974 248024 671030 248033
rect 670974 247959 671030 247968
rect 670976 235952 671028 235958
rect 670976 235894 671028 235900
rect 670988 224954 671016 235894
rect 671160 234252 671212 234258
rect 671160 234194 671212 234200
rect 670896 224926 671016 224954
rect 670896 215294 670924 224926
rect 671172 224777 671200 234194
rect 671356 224954 671384 258431
rect 671540 237046 671568 302223
rect 672552 287881 672580 304263
rect 672736 302234 672764 348463
rect 673012 337249 673040 351319
rect 673366 349752 673422 349761
rect 673366 349687 673422 349696
rect 672998 337240 673054 337249
rect 672998 337175 673054 337184
rect 673380 335617 673408 349687
rect 673550 349344 673606 349353
rect 673550 349279 673606 349288
rect 673366 335608 673422 335617
rect 673366 335543 673422 335552
rect 673564 332761 673592 349279
rect 673748 333985 673776 352543
rect 673918 348936 673974 348945
rect 673918 348871 673974 348880
rect 673734 333976 673790 333985
rect 673734 333911 673790 333920
rect 673550 332752 673606 332761
rect 673550 332687 673606 332696
rect 673932 331265 673960 348871
rect 673918 331256 673974 331265
rect 673918 331191 673974 331200
rect 674116 325694 674144 354583
rect 674746 354240 674802 354249
rect 674746 354175 674802 354184
rect 674286 350976 674342 350985
rect 674286 350911 674342 350920
rect 674300 345014 674328 350911
rect 674562 350568 674618 350577
rect 674562 350503 674618 350512
rect 674576 345014 674604 350503
rect 674300 344986 674420 345014
rect 674576 344986 674696 345014
rect 674392 336598 674420 344986
rect 674380 336592 674432 336598
rect 674380 336534 674432 336540
rect 674668 330049 674696 344986
rect 674760 339402 674788 354175
rect 675588 352889 675616 358255
rect 675942 357912 675998 357921
rect 675942 357847 675998 357856
rect 675956 356561 675984 357847
rect 675942 356552 675998 356561
rect 675942 356487 675998 356496
rect 675850 353832 675906 353841
rect 675850 353767 675906 353776
rect 675574 352880 675630 352889
rect 675574 352815 675630 352824
rect 675864 351937 675892 353767
rect 675850 351928 675906 351937
rect 675850 351863 675906 351872
rect 676034 351792 676090 351801
rect 676034 351727 676090 351736
rect 676048 347478 676076 351727
rect 683118 347712 683174 347721
rect 683118 347647 683174 347656
rect 676036 347472 676088 347478
rect 676036 347414 676088 347420
rect 676496 347472 676548 347478
rect 676496 347414 676548 347420
rect 676034 347304 676090 347313
rect 676034 347239 676090 347248
rect 676048 345681 676076 347239
rect 676508 346633 676536 347414
rect 676494 346624 676550 346633
rect 676494 346559 676550 346568
rect 683132 346497 683160 347647
rect 683118 346488 683174 346497
rect 683118 346423 683174 346432
rect 676034 345672 676090 345681
rect 676034 345607 676090 345616
rect 675128 341074 675418 341102
rect 674760 339386 674880 339402
rect 674760 339380 674892 339386
rect 674760 339374 674840 339380
rect 674840 339322 674892 339328
rect 675128 338745 675156 341074
rect 675574 340776 675630 340785
rect 675574 340711 675630 340720
rect 675588 340544 675616 340711
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675772 339864 675800 340167
rect 675484 339380 675536 339386
rect 675484 339322 675536 339328
rect 675496 339252 675524 339322
rect 675114 338736 675170 338745
rect 675114 338671 675170 338680
rect 675666 337784 675722 337793
rect 675666 337719 675722 337728
rect 675680 337416 675708 337719
rect 675114 337240 675170 337249
rect 675114 337175 675170 337184
rect 675128 336857 675156 337175
rect 675128 336829 675418 336857
rect 675392 336592 675444 336598
rect 675392 336534 675444 336540
rect 675404 336192 675432 336534
rect 675114 335608 675170 335617
rect 675170 335566 675340 335594
rect 675114 335543 675170 335552
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675312 335430 675432 335458
rect 675114 333976 675170 333985
rect 675114 333911 675170 333920
rect 675128 333078 675156 333911
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 675114 332344 675170 332353
rect 675114 332279 675170 332288
rect 675128 331889 675156 332279
rect 675128 331861 675418 331889
rect 675114 331256 675170 331265
rect 675170 331214 675418 331242
rect 675114 331191 675170 331200
rect 674668 330021 675418 330049
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675128 327542 675418 327570
rect 674116 325666 674420 325694
rect 673366 312760 673422 312769
rect 673366 312695 673422 312704
rect 673182 311264 673238 311273
rect 673182 311199 673238 311208
rect 672998 305552 673054 305561
rect 672998 305487 673054 305496
rect 672736 302206 672856 302234
rect 672538 287872 672594 287881
rect 672538 287807 672594 287816
rect 672264 287088 672316 287094
rect 672264 287030 672316 287036
rect 672080 284368 672132 284374
rect 672080 284310 672132 284316
rect 671894 262168 671950 262177
rect 671894 262103 671950 262112
rect 671710 260944 671766 260953
rect 671710 260879 671766 260888
rect 671724 246945 671752 260879
rect 671710 246936 671766 246945
rect 671710 246871 671766 246880
rect 671528 237040 671580 237046
rect 671528 236982 671580 236988
rect 671528 236632 671580 236638
rect 671528 236574 671580 236580
rect 671356 224926 671476 224954
rect 671158 224768 671214 224777
rect 671158 224703 671214 224712
rect 671252 224460 671304 224466
rect 671252 224402 671304 224408
rect 671264 224233 671292 224402
rect 671250 224224 671306 224233
rect 671250 224159 671306 224168
rect 671252 223848 671304 223854
rect 671250 223816 671252 223825
rect 671304 223816 671306 223825
rect 671448 223802 671476 224926
rect 671540 223938 671568 236574
rect 671712 236496 671764 236502
rect 671712 236438 671764 236444
rect 671724 224954 671752 236438
rect 671908 234394 671936 262103
rect 672092 246265 672120 284310
rect 672078 246256 672134 246265
rect 672078 246191 672134 246200
rect 672276 244274 672304 287030
rect 672828 285002 672856 302206
rect 673012 285569 673040 305487
rect 672998 285560 673054 285569
rect 672998 285495 673054 285504
rect 672644 284974 672856 285002
rect 672644 277394 672672 284974
rect 672814 283928 672870 283937
rect 672814 283863 672870 283872
rect 672828 277394 672856 283863
rect 672644 277366 672764 277394
rect 672828 277366 672948 277394
rect 672736 244274 672764 277366
rect 672920 244274 672948 277366
rect 673196 266665 673224 311199
rect 673380 267481 673408 312695
rect 674194 310448 674250 310457
rect 674194 310383 674250 310392
rect 674010 303920 674066 303929
rect 674010 303855 674066 303864
rect 673642 303512 673698 303521
rect 673642 303447 673698 303456
rect 673366 267472 673422 267481
rect 673366 267407 673422 267416
rect 673182 266656 673238 266665
rect 673182 266591 673238 266600
rect 673366 260536 673422 260545
rect 673366 260471 673422 260480
rect 673182 258904 673238 258913
rect 673182 258839 673238 258848
rect 672276 244246 672488 244274
rect 672736 244246 672856 244274
rect 672920 244246 673040 244274
rect 672080 236836 672132 236842
rect 672080 236778 672132 236784
rect 672092 235822 672120 236778
rect 672080 235816 672132 235822
rect 672080 235758 672132 235764
rect 671896 234388 671948 234394
rect 671896 234330 671948 234336
rect 671894 232520 671950 232529
rect 671894 232455 671896 232464
rect 671948 232455 671950 232464
rect 671896 232426 671948 232432
rect 671894 231568 671950 231577
rect 671894 231503 671896 231512
rect 671948 231503 671950 231512
rect 671896 231474 671948 231480
rect 672080 230648 672132 230654
rect 672080 230590 672132 230596
rect 672092 228410 672120 230590
rect 672080 228404 672132 228410
rect 672080 228346 672132 228352
rect 672262 226128 672318 226137
rect 672080 226092 672132 226098
rect 672262 226063 672318 226072
rect 672080 226034 672132 226040
rect 671896 225480 671948 225486
rect 672092 225457 672120 226034
rect 672276 225894 672304 226063
rect 672264 225888 672316 225894
rect 672264 225830 672316 225836
rect 672262 225720 672318 225729
rect 672262 225655 672264 225664
rect 672316 225655 672318 225664
rect 672264 225626 672316 225632
rect 671896 225422 671948 225428
rect 672078 225448 672134 225457
rect 671908 225298 671936 225422
rect 672078 225383 672134 225392
rect 672262 225312 672318 225321
rect 671908 225270 672262 225298
rect 672262 225247 672318 225256
rect 672032 225176 672088 225185
rect 672032 225111 672034 225120
rect 672086 225111 672088 225120
rect 672034 225082 672086 225088
rect 672460 224954 672488 244246
rect 672632 235748 672684 235754
rect 672632 235690 672684 235696
rect 672644 233238 672672 235690
rect 672632 233232 672684 233238
rect 672632 233174 672684 233180
rect 672828 227882 672856 244246
rect 673012 236858 673040 244246
rect 673196 241097 673224 258839
rect 673182 241088 673238 241097
rect 673182 241023 673238 241032
rect 673380 240281 673408 260471
rect 673656 244274 673684 303447
rect 674024 286521 674052 303855
rect 674010 286512 674066 286521
rect 674010 286447 674066 286456
rect 673918 267064 673974 267073
rect 673918 266999 673974 267008
rect 673564 244246 673684 244274
rect 673366 240272 673422 240281
rect 673366 240207 673422 240216
rect 673012 236830 673316 236858
rect 673090 236736 673146 236745
rect 672966 236706 673090 236722
rect 672954 236700 673090 236706
rect 673006 236694 673090 236700
rect 673090 236671 673146 236680
rect 672954 236642 673006 236648
rect 673288 236586 673316 236830
rect 672736 227854 672856 227882
rect 672920 236558 673316 236586
rect 672736 227798 672764 227854
rect 672724 227792 672776 227798
rect 672724 227734 672776 227740
rect 672724 226432 672776 226438
rect 672722 226400 672724 226409
rect 672776 226400 672778 226409
rect 672722 226335 672778 226344
rect 672604 226160 672656 226166
rect 672604 226102 672656 226108
rect 672616 225865 672644 226102
rect 672616 225856 672686 225865
rect 672616 225814 672630 225856
rect 672630 225791 672686 225800
rect 671724 224926 672028 224954
rect 671820 224732 671872 224738
rect 671820 224674 671872 224680
rect 671832 224505 671860 224674
rect 671818 224496 671874 224505
rect 671818 224431 671874 224440
rect 672000 223938 672028 224926
rect 671540 223910 671844 223938
rect 671448 223774 671568 223802
rect 671250 223751 671306 223760
rect 671160 223576 671212 223582
rect 671160 223518 671212 223524
rect 671022 223440 671074 223446
rect 671020 223408 671022 223417
rect 671074 223408 671076 223417
rect 671020 223343 671076 223352
rect 671172 223258 671200 223518
rect 671172 223230 671384 223258
rect 671158 223136 671214 223145
rect 671158 223071 671214 223080
rect 670896 215266 671016 215294
rect 670790 210488 670846 210497
rect 670790 210423 670846 210432
rect 670790 209944 670846 209953
rect 670790 209879 670846 209888
rect 670804 193225 670832 209879
rect 670790 193216 670846 193225
rect 670790 193151 670846 193160
rect 670606 171048 670662 171057
rect 670606 170983 670662 170992
rect 670606 170368 670662 170377
rect 670606 170303 670662 170312
rect 670332 160064 670384 160070
rect 670332 160006 670384 160012
rect 670148 148776 670200 148782
rect 670148 148718 670200 148724
rect 670620 147665 670648 170303
rect 670988 157334 671016 215266
rect 671172 177993 671200 223071
rect 671356 219745 671384 223230
rect 671342 219736 671398 219745
rect 671342 219671 671398 219680
rect 671540 218770 671568 223774
rect 671816 222194 671844 223910
rect 671356 218742 671568 218770
rect 671632 222166 671844 222194
rect 671908 223910 672028 223938
rect 672276 224926 672488 224954
rect 671158 177984 671214 177993
rect 671158 177919 671214 177928
rect 670804 157306 671016 157334
rect 670804 155174 670832 157306
rect 670792 155168 670844 155174
rect 670792 155110 670844 155116
rect 670606 147656 670662 147665
rect 670606 147591 670662 147600
rect 671356 138014 671384 218742
rect 671632 212534 671660 222166
rect 671908 219042 671936 223910
rect 672078 223816 672134 223825
rect 672078 223751 672134 223760
rect 672092 219065 672120 223751
rect 671540 212506 671660 212534
rect 671724 219014 671936 219042
rect 672078 219056 672134 219065
rect 671540 145353 671568 212506
rect 671724 150249 671752 219014
rect 672078 218991 672134 219000
rect 671894 216608 671950 216617
rect 671894 216543 671950 216552
rect 671908 204513 671936 216543
rect 671894 204504 671950 204513
rect 671894 204439 671950 204448
rect 672276 180305 672304 224926
rect 672722 224768 672778 224777
rect 672722 224703 672778 224712
rect 672446 223408 672502 223417
rect 672446 223343 672502 223352
rect 672460 217297 672488 223343
rect 672736 222873 672764 224703
rect 672722 222864 672778 222873
rect 672722 222799 672778 222808
rect 672630 220280 672686 220289
rect 672630 220215 672686 220224
rect 672446 217288 672502 217297
rect 672446 217223 672502 217232
rect 672644 215294 672672 220215
rect 672368 215266 672672 215294
rect 672368 190454 672396 215266
rect 672538 213752 672594 213761
rect 672538 213687 672594 213696
rect 672552 196353 672580 213687
rect 672722 213344 672778 213353
rect 672722 213279 672778 213288
rect 672538 196344 672594 196353
rect 672538 196279 672594 196288
rect 672368 190426 672580 190454
rect 672262 180296 672318 180305
rect 672262 180231 672318 180240
rect 672354 176080 672410 176089
rect 672354 176015 672410 176024
rect 671986 170776 672042 170785
rect 671986 170711 672042 170720
rect 672000 154465 672028 170711
rect 672170 169144 672226 169153
rect 672170 169079 672226 169088
rect 671986 154456 672042 154465
rect 671986 154391 672042 154400
rect 672184 153105 672212 169079
rect 672170 153096 672226 153105
rect 672170 153031 672226 153040
rect 671710 150240 671766 150249
rect 671710 150175 671766 150184
rect 671526 145344 671582 145353
rect 671526 145279 671582 145288
rect 670804 137986 671384 138014
rect 669964 136264 670016 136270
rect 669964 136206 670016 136212
rect 669226 133784 669282 133793
rect 669226 133719 669282 133728
rect 669240 132705 669268 133719
rect 669226 132696 669282 132705
rect 669226 132631 669282 132640
rect 668950 131200 669006 131209
rect 668950 131135 669006 131144
rect 668766 130656 668822 130665
rect 668766 130591 668822 130600
rect 668584 129736 668636 129742
rect 668584 129678 668636 129684
rect 668596 129033 668624 129678
rect 668582 129024 668638 129033
rect 668582 128959 668638 128968
rect 668582 127800 668638 127809
rect 668582 127735 668638 127744
rect 668030 125352 668086 125361
rect 668030 125287 668086 125296
rect 667202 116104 667258 116113
rect 667202 116039 667258 116048
rect 590290 115016 590346 115025
rect 590290 114951 590346 114960
rect 590108 112464 590160 112470
rect 590108 112406 590160 112412
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589476 110498 589504 111687
rect 589464 110492 589516 110498
rect 589464 110434 589516 110440
rect 589462 110120 589518 110129
rect 589462 110055 589518 110064
rect 589476 109138 589504 110055
rect 589464 109132 589516 109138
rect 589464 109074 589516 109080
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589830 105224 589886 105233
rect 589830 105159 589886 105168
rect 589844 104922 589872 105159
rect 589832 104916 589884 104922
rect 589832 104858 589884 104864
rect 590304 103514 590332 114951
rect 668216 111512 668268 111518
rect 668216 111454 668268 111460
rect 668228 111081 668256 111454
rect 668214 111072 668270 111081
rect 668214 111007 668270 111016
rect 666650 109372 666706 109381
rect 666650 109307 666706 109316
rect 666664 103514 666692 109307
rect 667940 108860 667992 108866
rect 667940 108802 667992 108808
rect 667952 107817 667980 108802
rect 667938 107808 667994 107817
rect 667938 107743 667994 107752
rect 668122 106176 668178 106185
rect 668122 106111 668178 106120
rect 589936 103486 590332 103514
rect 666572 103486 666692 103514
rect 588728 103420 588780 103426
rect 588728 103362 588780 103368
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100162 589504 101895
rect 589464 100156 589516 100162
rect 589464 100098 589516 100104
rect 589936 88330 589964 103486
rect 592684 100020 592736 100026
rect 592684 99962 592736 99968
rect 595272 100014 595608 100042
rect 591304 96076 591356 96082
rect 591304 96018 591356 96024
rect 589924 88324 589976 88330
rect 589924 88266 589976 88272
rect 588544 73160 588596 73166
rect 588544 73102 588596 73108
rect 587164 62076 587216 62082
rect 587164 62018 587216 62024
rect 591316 54505 591344 96018
rect 592696 64870 592724 99962
rect 595272 99142 595300 100014
rect 596330 99770 596358 100028
rect 596284 99742 596358 99770
rect 596468 100014 597080 100042
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 594064 95940 594116 95946
rect 594064 95882 594116 95888
rect 592684 64864 592736 64870
rect 592684 64806 592736 64812
rect 594076 57934 594104 95882
rect 595272 93854 595300 99078
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 594064 57928 594116 57934
rect 594064 57870 594116 57876
rect 591302 54496 591358 54505
rect 591302 54431 591358 54440
rect 596284 54398 596312 99742
rect 596468 55214 596496 100014
rect 597802 99770 597830 100028
rect 598216 100014 598552 100042
rect 599136 100014 599288 100042
rect 599688 100014 600024 100042
rect 600332 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602632 100014 602968 100042
rect 603092 100014 603704 100042
rect 597802 99742 597876 99770
rect 597652 96960 597704 96966
rect 597652 96902 597704 96908
rect 596456 55208 596508 55214
rect 596456 55150 596508 55156
rect 597664 54942 597692 96902
rect 597848 55078 597876 99742
rect 598216 96966 598244 100014
rect 598204 96960 598256 96966
rect 598204 96902 598256 96908
rect 598940 96960 598992 96966
rect 598940 96902 598992 96908
rect 598952 56030 598980 96902
rect 598940 56024 598992 56030
rect 598940 55966 598992 55972
rect 597836 55072 597888 55078
rect 597836 55014 597888 55020
rect 597652 54936 597704 54942
rect 597652 54878 597704 54884
rect 599136 54806 599164 100014
rect 599688 96966 599716 100014
rect 599676 96960 599728 96966
rect 599676 96902 599728 96908
rect 600332 57254 600360 100014
rect 600884 84194 600912 100014
rect 600516 84166 600912 84194
rect 600516 79354 600544 84166
rect 600504 79348 600556 79354
rect 600504 79290 600556 79296
rect 600320 57248 600372 57254
rect 600320 57190 600372 57196
rect 601896 55894 601924 100014
rect 602632 96082 602660 100014
rect 602620 96076 602672 96082
rect 602620 96018 602672 96024
rect 603092 58682 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613884 100042
rect 604426 99742 604500 99770
rect 604472 58818 604500 99742
rect 605484 97442 605512 100014
rect 605472 97436 605524 97442
rect 605472 97378 605524 97384
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606956 91798 606984 100014
rect 607128 96960 607180 96966
rect 607128 96902 607180 96908
rect 606944 91792 606996 91798
rect 606944 91734 606996 91740
rect 607140 75342 607168 96902
rect 607692 94518 607720 100014
rect 607680 94512 607732 94518
rect 607680 94454 607732 94460
rect 608520 84182 608548 100014
rect 609164 96762 609192 100014
rect 609152 96756 609204 96762
rect 609152 96698 609204 96704
rect 609704 96756 609756 96762
rect 609704 96698 609756 96704
rect 609716 93158 609744 96698
rect 609704 93152 609756 93158
rect 609704 93094 609756 93100
rect 609900 85542 609928 100014
rect 610636 96082 610664 100014
rect 610624 96076 610676 96082
rect 610624 96018 610676 96024
rect 611280 91050 611308 100014
rect 611912 97436 611964 97442
rect 611912 97378 611964 97384
rect 611924 93854 611952 97378
rect 612108 96898 612136 100014
rect 612660 97442 612688 100014
rect 612648 97436 612700 97442
rect 612648 97378 612700 97384
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 611924 93826 612044 93854
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 612016 76702 612044 93826
rect 612660 79354 612688 96834
rect 613856 80850 613884 100014
rect 613994 99770 614022 100028
rect 614744 100014 615264 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613994 99742 614068 99770
rect 613844 80844 613896 80850
rect 613844 80786 613896 80792
rect 614040 79490 614068 99742
rect 615236 93854 615264 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 94994 616552 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616512 94988 616564 94994
rect 616512 94930 616564 94936
rect 615236 93826 615448 93854
rect 615420 80986 615448 93826
rect 615408 80980 615460 80986
rect 615408 80922 615460 80928
rect 614028 79484 614080 79490
rect 614028 79426 614080 79432
rect 612648 79348 612700 79354
rect 612648 79290 612700 79296
rect 612004 76696 612056 76702
rect 612004 76638 612056 76644
rect 616800 75478 616828 96902
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91186 618208 96834
rect 619560 93838 619588 100014
rect 620204 97850 620232 100014
rect 620192 97844 620244 97850
rect 620192 97786 620244 97792
rect 620284 97436 620336 97442
rect 620284 97378 620336 97384
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 618628 93152 618680 93158
rect 618628 93094 618680 93100
rect 618168 91180 618220 91186
rect 618168 91122 618220 91128
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 618180 88194 618208 90986
rect 618168 88188 618220 88194
rect 618168 88130 618220 88136
rect 618640 85406 618668 93094
rect 618628 85400 618680 85406
rect 618628 85342 618680 85348
rect 620296 76838 620324 97378
rect 620940 95198 620968 100014
rect 621676 97442 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 621664 97436 621716 97442
rect 621664 97378 621716 97384
rect 623148 97306 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 624620 99074 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 624608 99068 624660 99074
rect 624608 99010 624660 99016
rect 625080 98938 625108 99742
rect 625068 98932 625120 98938
rect 625068 98874 625120 98880
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 623136 97300 623188 97306
rect 623136 97242 623188 97248
rect 621664 96076 621716 96082
rect 621664 96018 621716 96024
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620836 94512 620888 94518
rect 620836 94454 620888 94460
rect 620848 89690 620876 94454
rect 620836 89684 620888 89690
rect 620836 89626 620888 89632
rect 621676 86358 621704 96018
rect 625436 95192 625488 95198
rect 625436 95134 625488 95140
rect 624976 94988 625028 94994
rect 624976 94930 625028 94936
rect 622400 91792 622452 91798
rect 622400 91734 622452 91740
rect 622412 88330 622440 91734
rect 624988 88369 625016 94930
rect 625448 94489 625476 95134
rect 625434 94480 625490 94489
rect 625434 94415 625490 94424
rect 625816 92041 625844 97922
rect 626092 97170 626120 100014
rect 626356 97844 626408 97850
rect 626356 97786 626408 97792
rect 626080 97164 626132 97170
rect 626080 97106 626132 97112
rect 626172 93832 626224 93838
rect 626172 93774 626224 93780
rect 626184 92857 626212 93774
rect 626368 93673 626396 97786
rect 626828 96898 626856 100014
rect 627564 97578 627592 100014
rect 628300 97850 628328 100014
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 97986 629800 100014
rect 630508 98666 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 629760 97980 629812 97986
rect 629760 97922 629812 97928
rect 628288 97844 628340 97850
rect 628288 97786 628340 97792
rect 627552 97572 627604 97578
rect 627552 97514 627604 97520
rect 629300 97436 629352 97442
rect 629300 97378 629352 97384
rect 626816 96892 626868 96898
rect 626816 96834 626868 96840
rect 629312 95826 629340 97378
rect 630784 95826 630812 99282
rect 631244 97714 631272 100014
rect 631416 98320 631468 98326
rect 631416 98262 631468 98268
rect 631428 97850 631456 98262
rect 631416 97844 631468 97850
rect 631416 97786 631468 97792
rect 631232 97708 631284 97714
rect 631232 97650 631284 97656
rect 631980 97442 632008 100014
rect 632716 97850 632744 100014
rect 632704 97844 632756 97850
rect 632704 97786 632756 97792
rect 631968 97436 632020 97442
rect 631968 97378 632020 97384
rect 633268 97306 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 632060 97300 632112 97306
rect 632060 97242 632112 97248
rect 633256 97300 633308 97306
rect 633256 97242 633308 97248
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97242
rect 633452 95826 633480 99146
rect 633624 98184 633676 98190
rect 633624 98126 633676 98132
rect 633636 97578 633664 98126
rect 633624 97572 633676 97578
rect 633624 97514 633676 97520
rect 633808 97572 633860 97578
rect 633808 97514 633860 97520
rect 633820 97170 633848 97514
rect 634188 97170 634216 100014
rect 633808 97164 633860 97170
rect 633808 97106 633860 97112
rect 634176 97164 634228 97170
rect 634176 97106 634228 97112
rect 634740 97034 634768 100014
rect 635004 99068 635056 99074
rect 635004 99010 635056 99016
rect 634728 97028 634780 97034
rect 634728 96970 634780 96976
rect 635016 95826 635044 99010
rect 635568 96937 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635554 96928 635610 96937
rect 635554 96863 635610 96872
rect 635752 95985 635780 100014
rect 636292 98932 636344 98938
rect 636292 98874 636344 98880
rect 635738 95976 635794 95985
rect 635738 95911 635794 95920
rect 636304 95826 636332 98874
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96354 637620 99742
rect 637764 97572 637816 97578
rect 637764 97514 637816 97520
rect 637580 96348 637632 96354
rect 637580 96290 637632 96296
rect 637776 95826 637804 97514
rect 638604 96490 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 638592 96484 638644 96490
rect 638592 96426 638644 96432
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 639064 95810 639092 99742
rect 639236 96892 639288 96898
rect 639236 96834 639288 96840
rect 639248 95826 639276 96834
rect 640076 96626 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640064 96620 640116 96626
rect 640064 96562 640116 96568
rect 640536 96082 640564 99742
rect 640708 98184 640760 98190
rect 640708 98126 640760 98132
rect 640524 96076 640576 96082
rect 640524 96018 640576 96024
rect 640720 95826 640748 98126
rect 641548 96490 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96529 642036 99742
rect 642180 98320 642232 98326
rect 642180 98262 642232 98268
rect 641994 96520 642050 96529
rect 641352 96484 641404 96490
rect 641352 96426 641404 96432
rect 641536 96484 641588 96490
rect 641994 96455 642050 96464
rect 641536 96426 641588 96432
rect 639052 95804 639104 95810
rect 639248 95798 639584 95826
rect 640720 95798 641056 95826
rect 639052 95746 639104 95752
rect 641364 95470 641392 96426
rect 642192 95826 642220 98262
rect 643020 97578 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 643434 99742 643508 99770
rect 643008 97572 643060 97578
rect 643008 97514 643060 97520
rect 642192 95798 642528 95826
rect 643480 95470 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643664 95826 643692 98738
rect 644308 96830 644336 100014
rect 644906 99770 644934 100028
rect 645656 100014 645808 100042
rect 644906 99742 644980 99770
rect 644296 96824 644348 96830
rect 644296 96766 644348 96772
rect 644952 96218 644980 99742
rect 645308 98048 645360 98054
rect 645308 97990 645360 97996
rect 645124 96620 645176 96626
rect 645124 96562 645176 96568
rect 644940 96212 644992 96218
rect 644940 96154 644992 96160
rect 643664 95798 644000 95826
rect 645136 95674 645164 96562
rect 645320 95826 645348 97990
rect 645582 96112 645638 96121
rect 645582 96047 645584 96056
rect 645636 96047 645638 96056
rect 645584 96018 645636 96024
rect 645320 95798 645472 95826
rect 645124 95668 645176 95674
rect 645124 95610 645176 95616
rect 645780 95577 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648292 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 646424 96626 646452 99742
rect 647160 98802 647188 99742
rect 647148 98796 647200 98802
rect 647148 98738 647200 98744
rect 646596 98660 646648 98666
rect 646596 98602 646648 98608
rect 646412 96620 646464 96626
rect 646412 96562 646464 96568
rect 646608 95826 646636 98602
rect 647700 97844 647752 97850
rect 647700 97786 647752 97792
rect 647332 97708 647384 97714
rect 647332 97650 647384 97656
rect 647148 97028 647200 97034
rect 647148 96970 647200 96976
rect 646608 95798 646944 95826
rect 645766 95568 645822 95577
rect 645766 95503 645822 95512
rect 641352 95464 641404 95470
rect 641352 95406 641404 95412
rect 643468 95464 643520 95470
rect 643468 95406 643520 95412
rect 647160 95062 647188 96970
rect 647148 95056 647200 95062
rect 647344 95033 647372 97650
rect 647514 96112 647570 96121
rect 647514 96047 647516 96056
rect 647568 96047 647570 96056
rect 647516 96018 647568 96024
rect 647514 95568 647570 95577
rect 647514 95503 647570 95512
rect 647528 95334 647556 95503
rect 647516 95328 647568 95334
rect 647516 95270 647568 95276
rect 647516 95192 647568 95198
rect 647516 95134 647568 95140
rect 647148 94998 647200 95004
rect 647330 95024 647386 95033
rect 647330 94959 647386 94968
rect 626354 93664 626410 93673
rect 626354 93599 626410 93608
rect 626170 92848 626226 92857
rect 626170 92783 626226 92792
rect 647528 92478 647556 95134
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 647516 92472 647568 92478
rect 647516 92414 647568 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626460 91225 626488 92414
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 647712 89865 647740 97786
rect 648068 96212 648120 96218
rect 648068 96154 648120 96160
rect 648080 95538 648108 96154
rect 648068 95532 648120 95538
rect 648068 95474 648120 95480
rect 647884 95464 647936 95470
rect 647884 95406 647936 95412
rect 647698 89856 647754 89865
rect 647698 89791 647754 89800
rect 626448 89684 626500 89690
rect 626448 89626 626500 89632
rect 626262 89584 626318 89593
rect 626262 89519 626318 89528
rect 626276 88369 626304 89519
rect 626460 88777 626488 89626
rect 626446 88768 626502 88777
rect 626446 88703 626502 88712
rect 624974 88360 625030 88369
rect 622400 88324 622452 88330
rect 624974 88295 625030 88304
rect 626262 88360 626318 88369
rect 626262 88295 626318 88304
rect 626448 88324 626500 88330
rect 622400 88266 622452 88272
rect 626448 88266 626500 88272
rect 626264 88188 626316 88194
rect 626264 88130 626316 88136
rect 626276 87145 626304 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 626262 87136 626318 87145
rect 626262 87071 626318 87080
rect 647896 86358 647924 95406
rect 648264 87038 648292 100014
rect 648620 97436 648672 97442
rect 648620 97378 648672 97384
rect 648436 96484 648488 96490
rect 648436 96426 648488 96432
rect 648448 96218 648476 96426
rect 648632 96370 648660 97378
rect 648908 96490 648936 100014
rect 649080 97164 649132 97170
rect 649080 97106 649132 97112
rect 648896 96484 648948 96490
rect 648896 96426 648948 96432
rect 648632 96342 648844 96370
rect 648436 96212 648488 96218
rect 648436 96154 648488 96160
rect 648620 95804 648672 95810
rect 648620 95746 648672 95752
rect 648632 90846 648660 95746
rect 648816 92041 648844 96342
rect 648802 92032 648858 92041
rect 648802 91967 648858 91976
rect 648620 90840 648672 90846
rect 648620 90782 648672 90788
rect 649092 89714 649120 97106
rect 648632 89686 649120 89714
rect 648252 87032 648304 87038
rect 648252 86974 648304 86980
rect 621664 86352 621716 86358
rect 626448 86352 626500 86358
rect 621664 86294 621716 86300
rect 626446 86320 626448 86329
rect 647884 86352 647936 86358
rect 626500 86320 626502 86329
rect 647884 86294 647936 86300
rect 626446 86255 626502 86264
rect 626448 85536 626500 85542
rect 626446 85504 626448 85513
rect 626500 85504 626502 85513
rect 626446 85439 626502 85448
rect 625252 85400 625304 85406
rect 625252 85342 625304 85348
rect 625264 84697 625292 85342
rect 648632 84697 648660 89686
rect 649736 88806 649764 100014
rect 650380 97442 650408 100014
rect 650368 97436 650420 97442
rect 650368 97378 650420 97384
rect 650552 97300 650604 97306
rect 650552 97242 650604 97248
rect 650276 95192 650328 95198
rect 650276 95134 650328 95140
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 625250 84688 625306 84697
rect 625250 84623 625306 84632
rect 648618 84688 648674 84697
rect 648618 84623 648674 84632
rect 626448 84176 626500 84182
rect 626448 84118 626500 84124
rect 626460 83881 626488 84118
rect 626446 83872 626502 83881
rect 626446 83807 626502 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 81122 628788 83263
rect 650288 82249 650316 95134
rect 650564 87145 650592 97242
rect 651300 93634 651328 100014
rect 651852 97714 651880 100014
rect 651840 97708 651892 97714
rect 651840 97650 651892 97656
rect 652588 96626 652616 100014
rect 652208 96620 652260 96626
rect 652208 96562 652260 96568
rect 652576 96620 652628 96626
rect 652576 96562 652628 96568
rect 652024 95668 652076 95674
rect 652024 95610 652076 95616
rect 651288 93628 651340 93634
rect 651288 93570 651340 93576
rect 650550 87136 650606 87145
rect 650550 87071 650606 87080
rect 652036 86630 652064 95610
rect 652024 86624 652076 86630
rect 652024 86566 652076 86572
rect 652220 86494 652248 96562
rect 653324 95810 653352 100014
rect 653968 97850 653996 100014
rect 653956 97844 654008 97850
rect 653956 97786 654008 97792
rect 654324 97844 654376 97850
rect 654324 97786 654376 97792
rect 653312 95804 653364 95810
rect 653312 95746 653364 95752
rect 652392 95668 652444 95674
rect 652392 95610 652444 95616
rect 652404 95334 652432 95610
rect 652392 95328 652444 95334
rect 652392 95270 652444 95276
rect 654336 94217 654364 97786
rect 654796 96966 654824 100014
rect 655440 97850 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97844 655480 97850
rect 655428 97786 655480 97792
rect 654784 96960 654836 96966
rect 654784 96902 654836 96908
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 654322 94208 654378 94217
rect 654322 94143 654378 94152
rect 655440 93854 655468 96902
rect 655256 93826 655468 93854
rect 654692 93628 654744 93634
rect 654692 93570 654744 93576
rect 654704 93401 654732 93570
rect 654690 93392 654746 93401
rect 654690 93327 654746 93336
rect 655256 88330 655284 93826
rect 655428 92472 655480 92478
rect 655428 92414 655480 92420
rect 655440 91497 655468 92414
rect 655426 91488 655482 91497
rect 655426 91423 655482 91432
rect 655428 90840 655480 90846
rect 655428 90782 655480 90788
rect 655440 90681 655468 90782
rect 655426 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656820 97238 656848 100014
rect 656808 97232 656860 97238
rect 656808 97174 656860 97180
rect 656716 96960 656768 96966
rect 656716 96902 656768 96908
rect 656348 95668 656400 95674
rect 656348 95610 656400 95616
rect 656164 95532 656216 95538
rect 656164 95474 656216 95480
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 656176 86766 656204 95474
rect 656360 88670 656388 95610
rect 656348 88664 656400 88670
rect 656348 88606 656400 88612
rect 656728 86902 656756 96902
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658154 99742 658228 99770
rect 658200 97578 658228 99742
rect 659212 97986 659240 100014
rect 659200 97980 659252 97986
rect 659200 97922 659252 97928
rect 659948 97850 659976 100014
rect 660132 100014 660376 100042
rect 659936 97844 659988 97850
rect 659936 97786 659988 97792
rect 659568 97708 659620 97714
rect 659568 97650 659620 97656
rect 658004 97572 658056 97578
rect 658004 97514 658056 97520
rect 658188 97572 658240 97578
rect 658188 97514 658240 97520
rect 658016 97102 658044 97514
rect 658280 97436 658332 97442
rect 658280 97378 658332 97384
rect 658004 97096 658056 97102
rect 658004 97038 658056 97044
rect 658292 95132 658320 97378
rect 658832 96824 658884 96830
rect 658832 96766 658884 96772
rect 658844 95132 658872 96766
rect 659580 95132 659608 97650
rect 659844 97096 659896 97102
rect 659844 97038 659896 97044
rect 659856 95146 659884 97038
rect 660132 96966 660160 100014
rect 661960 98796 662012 98802
rect 661960 98738 662012 98744
rect 661408 97232 661460 97238
rect 661408 97174 661460 97180
rect 660120 96960 660172 96966
rect 660120 96902 660172 96908
rect 660672 96348 660724 96354
rect 660672 96290 660724 96296
rect 659856 95118 660146 95146
rect 660684 95132 660712 96290
rect 661420 95132 661448 97174
rect 661972 95132 662000 98738
rect 664168 97980 664220 97986
rect 664168 97922 664220 97928
rect 662512 97708 662564 97714
rect 662512 97650 662564 97656
rect 662524 95132 662552 97650
rect 663064 97572 663116 97578
rect 663064 97514 663116 97520
rect 663076 95132 663104 97514
rect 663800 96212 663852 96218
rect 663800 96154 663852 96160
rect 663812 93129 663840 96154
rect 663984 96076 664036 96082
rect 663984 96018 664036 96024
rect 663798 93120 663854 93129
rect 663798 93055 663854 93064
rect 663996 91769 664024 96018
rect 663982 91760 664038 91769
rect 663982 91695 664038 91704
rect 664180 88806 664208 97922
rect 665364 97844 665416 97850
rect 665364 97786 665416 97792
rect 664352 96620 664404 96626
rect 664352 96562 664404 96568
rect 664364 90681 664392 96562
rect 664536 96484 664588 96490
rect 664536 96426 664588 96432
rect 664350 90672 664406 90681
rect 664350 90607 664406 90616
rect 664548 89865 664576 96426
rect 665180 95804 665232 95810
rect 665180 95746 665232 95752
rect 664534 89856 664590 89865
rect 664534 89791 664590 89800
rect 665192 89049 665220 95746
rect 665376 93401 665404 97786
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665178 89040 665234 89049
rect 665178 88975 665234 88984
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 664168 88800 664220 88806
rect 664168 88742 664220 88748
rect 661986 88726 662368 88742
rect 657452 88664 657504 88670
rect 657504 88612 657754 88618
rect 657452 88606 657754 88612
rect 657464 88590 657754 88606
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656716 86896 656768 86902
rect 656716 86838 656768 86844
rect 656164 86760 656216 86766
rect 656164 86702 656216 86708
rect 657188 86494 657216 88196
rect 659580 86902 659608 88196
rect 659568 86896 659620 86902
rect 659568 86838 659620 86844
rect 660132 86630 660160 88196
rect 660684 86766 660712 88196
rect 660672 86760 660724 86766
rect 660672 86702 660724 86708
rect 660120 86624 660172 86630
rect 660120 86566 660172 86572
rect 652208 86488 652260 86494
rect 652208 86430 652260 86436
rect 657176 86488 657228 86494
rect 657176 86430 657228 86436
rect 661420 86358 661448 88196
rect 662524 87038 662552 88196
rect 662512 87032 662564 87038
rect 662512 86974 662564 86980
rect 661408 86352 661460 86358
rect 661408 86294 661460 86300
rect 650274 82240 650330 82249
rect 650274 82175 650330 82184
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 81116 628800 81122
rect 628748 81058 628800 81064
rect 629220 80034 629248 81631
rect 642456 81116 642508 81122
rect 642456 81058 642508 81064
rect 632808 80974 633144 81002
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 77988 631100 77994
rect 631048 77930 631100 77936
rect 628472 77716 628524 77722
rect 628472 77658 628524 77664
rect 628484 77450 628512 77658
rect 624424 77444 624476 77450
rect 624424 77386 624476 77392
rect 628472 77444 628524 77450
rect 628472 77386 628524 77392
rect 623042 77344 623098 77353
rect 623042 77279 623098 77288
rect 620284 76832 620336 76838
rect 620284 76774 620336 76780
rect 616788 75472 616840 75478
rect 616788 75414 616840 75420
rect 607128 75336 607180 75342
rect 607128 75278 607180 75284
rect 604460 58812 604512 58818
rect 604460 58754 604512 58760
rect 603080 58676 603132 58682
rect 603080 58618 603132 58624
rect 601884 55888 601936 55894
rect 601884 55830 601936 55836
rect 599124 54800 599176 54806
rect 599124 54742 599176 54748
rect 623056 54670 623084 77279
rect 624436 60042 624464 77386
rect 625804 77308 625856 77314
rect 625804 77250 625856 77256
rect 624424 60036 624476 60042
rect 624424 59978 624476 59984
rect 623044 54664 623096 54670
rect 623044 54606 623096 54612
rect 625816 54534 625844 77250
rect 628484 75290 628512 77386
rect 631060 77314 631088 77930
rect 632808 77722 632836 80974
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78130 633480 79970
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633440 78124 633492 78130
rect 633440 78066 633492 78072
rect 632796 77716 632848 77722
rect 632796 77658 632848 77664
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 631048 77308 631100 77314
rect 633898 77279 633954 77288
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75290 633940 77279
rect 636764 75290 636792 80650
rect 639602 77616 639658 77625
rect 639602 77551 639658 77560
rect 639616 75290 639644 77551
rect 642468 75290 642496 81058
rect 643080 80974 643140 81002
rect 643112 77994 643140 80974
rect 646320 80980 646372 80986
rect 646320 80922 646372 80928
rect 646044 79484 646096 79490
rect 646044 79426 646096 79432
rect 645308 78124 645360 78130
rect 645308 78066 645360 78072
rect 643100 77988 643152 77994
rect 643100 77930 643152 77936
rect 645320 75290 645348 78066
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 646056 74534 646084 79426
rect 646056 74506 646176 74534
rect 646148 67153 646176 74506
rect 646332 69193 646360 80922
rect 647332 80844 647384 80850
rect 647332 80786 647384 80792
rect 646688 75472 646740 75478
rect 646688 75414 646740 75420
rect 646504 75336 646556 75342
rect 646504 75278 646556 75284
rect 646516 74225 646544 75278
rect 646502 74216 646558 74225
rect 646502 74151 646558 74160
rect 646700 71777 646728 75414
rect 646686 71768 646742 71777
rect 646686 71703 646742 71712
rect 646318 69184 646374 69193
rect 646318 69119 646374 69128
rect 646134 67144 646190 67153
rect 646134 67079 646190 67088
rect 625988 66904 626040 66910
rect 625988 66846 626040 66852
rect 625804 54528 625856 54534
rect 625804 54470 625856 54476
rect 596272 54392 596324 54398
rect 596272 54334 596324 54340
rect 583024 54256 583076 54262
rect 583024 54198 583076 54204
rect 580448 54120 580500 54126
rect 580448 54062 580500 54068
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459834 53680 459890 53689
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 461674 53615 461730 53624
rect 462594 53680 462650 53689
rect 470322 53680 470378 53689
rect 462594 53615 462650 53624
rect 463332 53644 463384 53650
rect 130384 53372 130436 53378
rect 130384 53314 130436 53320
rect 129004 53236 129056 53242
rect 129004 53178 129056 53184
rect 51724 49156 51776 49162
rect 51724 49098 51776 49104
rect 45468 49020 45520 49026
rect 45468 48962 45520 48968
rect 128820 49020 128872 49026
rect 128820 48962 128872 48968
rect 128832 47870 128860 48962
rect 128820 47864 128872 47870
rect 128820 47806 128872 47812
rect 129016 46102 129044 53178
rect 129188 53100 129240 53106
rect 129188 53042 129240 53048
rect 129004 46096 129056 46102
rect 129004 46038 129056 46044
rect 43812 45212 43864 45218
rect 43812 45154 43864 45160
rect 129200 44538 129228 53042
rect 129372 51876 129424 51882
rect 129372 51818 129424 51824
rect 129384 45082 129412 51818
rect 129648 49156 129700 49162
rect 129648 49098 129700 49104
rect 129660 45422 129688 49098
rect 129648 45416 129700 45422
rect 129648 45358 129700 45364
rect 129372 45076 129424 45082
rect 129372 45018 129424 45024
rect 129188 44532 129240 44538
rect 129188 44474 129240 44480
rect 43628 44328 43680 44334
rect 129096 44328 129148 44334
rect 43628 44270 43680 44276
rect 129094 44296 129096 44305
rect 129148 44296 129150 44305
rect 129094 44231 129150 44240
rect 43444 44192 43496 44198
rect 43444 44134 43496 44140
rect 130396 44062 130424 53314
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 306024 51746 306052 53108
rect 130568 51740 130620 51746
rect 130568 51682 130620 51688
rect 145380 51740 145432 51746
rect 145380 51682 145432 51688
rect 306012 51740 306064 51746
rect 306012 51682 306064 51688
rect 130580 45966 130608 51682
rect 145392 50810 145420 51682
rect 145084 50782 145420 50810
rect 131028 50380 131080 50386
rect 131028 50322 131080 50328
rect 130752 47864 130804 47870
rect 130752 47806 130804 47812
rect 130568 45960 130620 45966
rect 130568 45902 130620 45908
rect 130764 44334 130792 47806
rect 131040 45370 131068 50322
rect 308048 50289 308076 53108
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459146 52828 459198 52834
rect 459146 52770 459198 52776
rect 459158 52564 459186 52770
rect 459848 52578 459876 53615
rect 460388 53508 460440 53514
rect 460388 53450 460440 53456
rect 460400 52578 460428 53450
rect 460768 52578 460796 53615
rect 461308 53100 461360 53106
rect 461308 53042 461360 53048
rect 461320 52578 461348 53042
rect 461688 52578 461716 53615
rect 462228 53372 462280 53378
rect 462228 53314 462280 53320
rect 462240 52578 462268 53314
rect 462608 52578 462636 53615
rect 463332 53586 463384 53592
rect 463516 53644 463568 53650
rect 463516 53586 463568 53592
rect 463884 53644 463936 53650
rect 463884 53586 463936 53592
rect 464068 53644 464120 53650
rect 464068 53586 464120 53592
rect 465908 53644 465960 53650
rect 471978 53680 472034 53689
rect 470322 53615 470324 53624
rect 465908 53586 465960 53592
rect 470376 53615 470378 53624
rect 470968 53644 471020 53650
rect 470324 53586 470376 53592
rect 470968 53586 471020 53592
rect 471152 53644 471204 53650
rect 471152 53586 471204 53592
rect 471704 53644 471756 53650
rect 471978 53615 471980 53624
rect 471704 53586 471756 53592
rect 472032 53615 472034 53624
rect 476764 53644 476816 53650
rect 471980 53586 472032 53592
rect 476764 53586 476816 53592
rect 479616 53644 479668 53650
rect 479616 53586 479668 53592
rect 479984 53644 480036 53650
rect 479984 53586 480036 53592
rect 480168 53644 480220 53650
rect 480168 53586 480220 53592
rect 463148 53236 463200 53242
rect 463148 53178 463200 53184
rect 463160 52578 463188 53178
rect 463344 52970 463372 53586
rect 463332 52964 463384 52970
rect 463332 52906 463384 52912
rect 463528 52578 463556 53586
rect 463896 53145 463924 53586
rect 463882 53136 463938 53145
rect 463882 53071 463938 53080
rect 463792 52964 463844 52970
rect 463792 52906 463844 52912
rect 459632 52550 459876 52578
rect 460092 52550 460428 52578
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461932 52550 462268 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463556 52578
rect 463804 52442 463832 52906
rect 464080 52578 464108 53586
rect 464988 53508 465040 53514
rect 464988 53450 465040 53456
rect 465000 52578 465028 53450
rect 465126 52828 465178 52834
rect 465126 52770 465178 52776
rect 464080 52550 464232 52578
rect 464692 52550 465028 52578
rect 465138 52564 465166 52770
rect 465920 52578 465948 53586
rect 470980 53417 471008 53586
rect 470966 53408 471022 53417
rect 470966 53343 471022 53352
rect 471164 53145 471192 53586
rect 471150 53136 471206 53145
rect 471150 53071 471206 53080
rect 471716 52698 471744 53586
rect 476776 53417 476804 53586
rect 476762 53408 476818 53417
rect 476762 53343 476818 53352
rect 479628 53242 479656 53586
rect 479616 53236 479668 53242
rect 479616 53178 479668 53184
rect 479996 52834 480024 53586
rect 480180 53106 480208 53586
rect 480168 53100 480220 53106
rect 480168 53042 480220 53048
rect 479984 52828 480036 52834
rect 479984 52770 480036 52776
rect 471704 52692 471756 52698
rect 471704 52634 471756 52640
rect 465612 52550 465948 52578
rect 463772 52414 463832 52442
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461072 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 462392 47654 462728 47682
rect 462852 47654 462912 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 131764 46096 131816 46102
rect 131764 46038 131816 46044
rect 131040 45354 131436 45370
rect 131040 45348 131448 45354
rect 131040 45342 131396 45348
rect 131396 45290 131448 45296
rect 131132 45218 131436 45234
rect 131120 45212 131448 45218
rect 131172 45206 131396 45212
rect 131120 45154 131172 45160
rect 131396 45154 131448 45160
rect 131580 44804 131632 44810
rect 131580 44746 131632 44752
rect 130752 44328 130804 44334
rect 130752 44270 130804 44276
rect 131592 44198 131620 44746
rect 131776 44702 131804 46038
rect 132500 45960 132552 45966
rect 132500 45902 132552 45908
rect 131764 44696 131816 44702
rect 131764 44638 131816 44644
rect 131948 44668 132000 44674
rect 131948 44610 132000 44616
rect 131960 44305 131988 44610
rect 132512 44402 132540 45902
rect 132960 45348 133012 45354
rect 132960 45290 133012 45296
rect 132500 44396 132552 44402
rect 132500 44338 132552 44344
rect 132972 44310 133000 45290
rect 133144 45212 133196 45218
rect 133144 45154 133196 45160
rect 131946 44296 132002 44305
rect 132960 44304 133012 44310
rect 132960 44246 133012 44252
rect 131946 44231 132002 44240
rect 133156 44198 133184 45154
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 458178 44432 458234 44441
rect 458178 44367 458234 44376
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 131580 44192 131632 44198
rect 131580 44134 131632 44140
rect 133144 44192 133196 44198
rect 133144 44134 133196 44140
rect 307298 44160 307354 44169
rect 307298 44095 307354 44104
rect 130384 44056 130436 44062
rect 130384 43998 130436 44004
rect 187332 42764 187384 42770
rect 187332 42706 187384 42712
rect 187344 42092 187372 42706
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 44095
rect 440240 43648 440292 43654
rect 419722 43616 419778 43625
rect 419722 43551 419778 43560
rect 440238 43616 440240 43625
rect 441068 43648 441120 43654
rect 440292 43616 440294 43625
rect 440238 43551 440294 43560
rect 441066 43616 441068 43625
rect 441120 43616 441122 43625
rect 441066 43551 441122 43560
rect 416594 42392 416650 42401
rect 419736 42364 419764 43551
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 441068 42764 441120 42770
rect 441068 42706 441120 42712
rect 449164 42764 449216 42770
rect 449164 42706 449216 42712
rect 416594 42327 416650 42336
rect 307004 42078 307340 42106
rect 404634 42120 404690 42129
rect 194322 42055 194378 42064
rect 404634 42055 404690 42064
rect 405186 42120 405242 42129
rect 415582 42120 415638 42129
rect 405242 42078 405582 42106
rect 415426 42078 415582 42106
rect 405186 42055 405242 42064
rect 416608 42092 416636 42327
rect 415582 42055 415638 42064
rect 404648 41886 404676 42055
rect 431236 42022 431264 42706
rect 441080 42022 441108 42706
rect 449176 42022 449204 42706
rect 454500 42356 454552 42362
rect 454500 42298 454552 42304
rect 431224 42016 431276 42022
rect 431224 41958 431276 41964
rect 441068 42016 441120 42022
rect 441068 41958 441120 41964
rect 449164 42016 449216 42022
rect 449164 41958 449216 41964
rect 404636 41880 404688 41886
rect 310426 41848 310482 41857
rect 310132 41806 310426 41834
rect 310426 41783 310482 41792
rect 311070 41848 311126 41857
rect 361946 41848 362002 41857
rect 361790 41806 361946 41834
rect 311070 41783 311126 41792
rect 365166 41848 365222 41857
rect 364918 41806 365166 41834
rect 361946 41783 362002 41792
rect 404636 41822 404688 41828
rect 365166 41783 365222 41792
rect 311084 41614 311112 41783
rect 420736 41744 420788 41750
rect 420736 41686 420788 41692
rect 427084 41744 427136 41750
rect 427084 41686 427136 41692
rect 311072 41608 311124 41614
rect 311072 41550 311124 41556
rect 420748 41478 420776 41686
rect 427096 41478 427124 41686
rect 454512 41614 454540 42298
rect 454500 41608 454552 41614
rect 454500 41550 454552 41556
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 427084 41472 427136 41478
rect 427084 41414 427136 41420
rect 458192 41177 458220 44367
rect 459204 41750 459232 47654
rect 459560 42492 459612 42498
rect 459560 42434 459612 42440
rect 459376 42016 459428 42022
rect 459572 41970 459600 42434
rect 459940 42106 459968 47654
rect 460124 42498 460152 47654
rect 460860 43897 460888 47654
rect 461044 44441 461072 47654
rect 461030 44432 461086 44441
rect 461030 44367 461086 44376
rect 460846 43888 460902 43897
rect 460846 43823 460902 43832
rect 461780 42945 461808 47654
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 460112 42492 460164 42498
rect 460112 42434 460164 42440
rect 459940 42078 460368 42106
rect 459428 41964 459600 41970
rect 459376 41958 459600 41964
rect 459388 41942 459600 41958
rect 461964 41857 461992 47654
rect 462700 43217 462728 47654
rect 462884 43625 462912 47654
rect 463068 47654 463312 47682
rect 462870 43616 462926 43625
rect 462870 43551 462926 43560
rect 462686 43208 462742 43217
rect 462686 43143 462742 43152
rect 463068 42362 463096 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463896 47654 464232 47682
rect 464692 47654 464752 47682
rect 463712 44441 463740 47382
rect 463698 44432 463754 44441
rect 463698 44367 463754 44376
rect 463896 44169 463924 47654
rect 464724 44577 464752 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46753 465120 47382
rect 465276 47025 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 465078 46744 465134 46753
rect 465078 46679 465134 46688
rect 626000 46510 626028 66846
rect 647344 64433 647372 80786
rect 648620 79348 648672 79354
rect 648620 79290 648672 79296
rect 647514 78160 647570 78169
rect 647514 78095 647570 78104
rect 647330 64424 647386 64433
rect 647330 64359 647386 64368
rect 647528 57361 647556 78095
rect 648632 59265 648660 79290
rect 648988 76832 649040 76838
rect 648988 76774 649040 76780
rect 649000 62121 649028 76774
rect 662420 76696 662472 76702
rect 662420 76638 662472 76644
rect 648986 62112 649042 62121
rect 648986 62047 649042 62056
rect 648618 59256 648674 59265
rect 648618 59191 648674 59200
rect 647514 57352 647570 57361
rect 647514 57287 647570 57296
rect 661590 48510 661646 48519
rect 661590 48445 661646 48454
rect 625988 46504 626040 46510
rect 625988 46446 626040 46452
rect 661604 45554 661632 48445
rect 661774 47789 661830 47798
rect 661774 47724 661830 47733
rect 661788 46510 661816 47724
rect 662432 47433 662460 76638
rect 666572 75206 666600 103486
rect 667938 102776 667994 102785
rect 667938 102711 667994 102720
rect 667952 100026 667980 102711
rect 667940 100020 667992 100026
rect 667940 99962 667992 99968
rect 668136 95962 668164 106111
rect 668306 104816 668362 104825
rect 668306 104751 668362 104760
rect 668320 104417 668348 104751
rect 668306 104408 668362 104417
rect 668306 104343 668362 104352
rect 668320 103514 668348 104343
rect 668044 95946 668164 95962
rect 668032 95940 668164 95946
rect 668084 95934 668164 95940
rect 668228 103486 668348 103514
rect 668032 95882 668084 95888
rect 668228 76566 668256 103486
rect 668596 102785 668624 127735
rect 668766 120048 668822 120057
rect 668766 119983 668822 119992
rect 668780 104825 668808 119983
rect 668964 119241 668992 131135
rect 669962 130928 670018 130937
rect 669962 130863 670018 130872
rect 669226 126032 669282 126041
rect 669226 125967 669282 125976
rect 669240 124137 669268 125967
rect 669226 124128 669282 124137
rect 669226 124063 669282 124072
rect 668950 119232 669006 119241
rect 668950 119167 669006 119176
rect 669226 117056 669282 117065
rect 669226 116991 669282 117000
rect 669240 114345 669268 116991
rect 669226 114336 669282 114345
rect 669226 114271 669282 114280
rect 669976 108866 670004 130863
rect 670804 129742 670832 137986
rect 672170 131744 672226 131753
rect 672170 131679 672226 131688
rect 670792 129736 670844 129742
rect 670792 129678 670844 129684
rect 672184 128354 672212 131679
rect 672368 131481 672396 176015
rect 672552 175681 672580 190426
rect 672538 175672 672594 175681
rect 672538 175607 672594 175616
rect 672538 168328 672594 168337
rect 672538 168263 672594 168272
rect 672354 131472 672410 131481
rect 672354 131407 672410 131416
rect 672552 131209 672580 168263
rect 672538 131200 672594 131209
rect 672538 131135 672594 131144
rect 672184 128326 672396 128354
rect 671986 126848 672042 126857
rect 671986 126783 672042 126792
rect 671526 122768 671582 122777
rect 671526 122703 671582 122712
rect 670698 121408 670754 121417
rect 670698 121343 670754 121352
rect 670712 111518 670740 121343
rect 671540 112713 671568 122703
rect 671526 112704 671582 112713
rect 671526 112639 671582 112648
rect 670700 111512 670752 111518
rect 670700 111454 670752 111460
rect 669964 108860 670016 108866
rect 669964 108802 670016 108808
rect 668766 104816 668822 104825
rect 668766 104751 668822 104760
rect 668582 102776 668638 102785
rect 668582 102711 668638 102720
rect 672000 99385 672028 126783
rect 672368 106185 672396 128326
rect 672736 126041 672764 213279
rect 672920 177721 672948 236558
rect 673184 236292 673236 236298
rect 673184 236234 673236 236240
rect 673196 236178 673224 236234
rect 673196 236150 673500 236178
rect 673276 235952 673328 235958
rect 673276 235894 673328 235900
rect 673092 235544 673144 235550
rect 673092 235486 673144 235492
rect 673104 224954 673132 235486
rect 673288 234977 673316 235894
rect 673274 234968 673330 234977
rect 673274 234903 673330 234912
rect 673472 234682 673500 236150
rect 673564 234818 673592 244246
rect 673932 239442 673960 266999
rect 674208 265849 674236 310383
rect 674392 310049 674420 325666
rect 675128 325281 675156 327542
rect 675312 326454 675432 326482
rect 675312 325553 675340 326454
rect 675404 326332 675432 326454
rect 675298 325544 675354 325553
rect 675298 325479 675354 325488
rect 675114 325272 675170 325281
rect 675114 325207 675170 325216
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676218 313984 676274 313993
rect 676218 313919 676274 313928
rect 674654 313032 674710 313041
rect 674654 312967 674710 312976
rect 674668 311953 674696 312967
rect 674838 312760 674894 312769
rect 674838 312695 674894 312704
rect 674852 312089 674880 312695
rect 674838 312080 674894 312089
rect 674838 312015 674894 312024
rect 674654 311944 674710 311953
rect 674654 311879 674710 311888
rect 674378 310040 674434 310049
rect 674378 309975 674434 309984
rect 674562 309632 674618 309641
rect 674562 309567 674618 309576
rect 674378 305144 674434 305153
rect 674378 305079 674434 305088
rect 674392 287026 674420 305079
rect 674380 287020 674432 287026
rect 674380 286962 674432 286968
rect 674378 283520 674434 283529
rect 674378 283455 674434 283464
rect 674392 267889 674420 283455
rect 674378 267880 674434 267889
rect 674378 267815 674434 267824
rect 674378 266248 674434 266257
rect 674378 266183 674434 266192
rect 674194 265840 674250 265849
rect 674194 265775 674250 265784
rect 674102 265432 674158 265441
rect 674102 265367 674158 265376
rect 674116 241913 674144 265367
rect 674392 263594 674420 266183
rect 674576 265033 674604 309567
rect 675850 309360 675906 309369
rect 676232 309346 676260 313919
rect 675906 309318 676260 309346
rect 675850 309295 675906 309304
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 675114 308000 675170 308009
rect 675114 307935 675170 307944
rect 674930 301880 674986 301889
rect 674930 301815 674986 301824
rect 674944 293570 674972 301815
rect 675128 297106 675156 307935
rect 676232 307834 676260 308366
rect 676220 307828 676272 307834
rect 676220 307770 676272 307776
rect 676864 307828 676916 307834
rect 676864 307770 676916 307776
rect 676034 307592 676090 307601
rect 676090 307550 676260 307578
rect 676034 307527 676090 307536
rect 676034 304736 676090 304745
rect 676034 304671 676090 304680
rect 675852 304156 675904 304162
rect 675852 304098 675904 304104
rect 675864 301889 675892 304098
rect 675850 301880 675906 301889
rect 675850 301815 675906 301824
rect 676048 300665 676076 304671
rect 676232 304162 676260 307550
rect 676494 305960 676550 305969
rect 676494 305895 676550 305904
rect 676220 304156 676272 304162
rect 676220 304098 676272 304104
rect 676508 301617 676536 305895
rect 676494 301608 676550 301617
rect 676494 301543 676550 301552
rect 676034 300656 676090 300665
rect 676034 300591 676090 300600
rect 676876 298110 676904 307770
rect 679622 306776 679678 306785
rect 679622 306711 679678 306720
rect 677598 306368 677654 306377
rect 677598 306303 677654 306312
rect 675852 298104 675904 298110
rect 675036 297078 675156 297106
rect 675496 298064 675852 298092
rect 675036 293706 675064 297078
rect 675496 296410 675524 298064
rect 675852 298046 675904 298052
rect 676864 298104 676916 298110
rect 676864 298046 676916 298052
rect 676128 297968 676180 297974
rect 676128 297910 676180 297916
rect 675944 297492 675996 297498
rect 675944 297434 675996 297440
rect 675956 296585 675984 297434
rect 676140 296857 676168 297910
rect 677612 297498 677640 306303
rect 679636 297974 679664 306711
rect 683026 302696 683082 302705
rect 683026 302631 683082 302640
rect 683040 299441 683068 302631
rect 683026 299432 683082 299441
rect 683026 299367 683082 299376
rect 679624 297968 679676 297974
rect 679624 297910 679676 297916
rect 677600 297492 677652 297498
rect 677600 297434 677652 297440
rect 676126 296848 676182 296857
rect 676126 296783 676182 296792
rect 675942 296576 675998 296585
rect 675942 296511 675998 296520
rect 675484 296404 675536 296410
rect 675484 296346 675536 296352
rect 675220 296058 675418 296086
rect 675220 293865 675248 296058
rect 675484 295792 675536 295798
rect 675484 295734 675536 295740
rect 675496 295528 675524 295734
rect 675574 295352 675630 295361
rect 675574 295287 675630 295296
rect 675588 294879 675616 295287
rect 675758 294536 675814 294545
rect 675758 294471 675814 294480
rect 675772 294236 675800 294471
rect 675206 293856 675262 293865
rect 675206 293791 675262 293800
rect 675036 293678 675340 293706
rect 674944 293542 675064 293570
rect 675036 288062 675064 293542
rect 675312 292574 675340 293678
rect 675312 292546 675432 292574
rect 675404 292400 675432 292546
rect 675574 292224 675630 292233
rect 675574 292159 675630 292168
rect 675588 291856 675616 292159
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675758 290864 675814 290873
rect 675758 290799 675814 290808
rect 675772 290564 675800 290799
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 675036 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675116 287020 675168 287026
rect 675116 286962 675168 286968
rect 675128 286906 675156 286962
rect 675128 286878 675340 286906
rect 675312 286770 675340 286878
rect 675404 286770 675432 286892
rect 675312 286742 675432 286770
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675666 283656 675722 283665
rect 675666 283591 675722 283600
rect 675680 283220 675708 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675772 281217 675800 281355
rect 675758 281208 675814 281217
rect 675758 281143 675814 281152
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 683132 268569 683160 271079
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683118 268560 683174 268569
rect 683118 268495 683174 268504
rect 674562 265024 674618 265033
rect 674562 264959 674618 264968
rect 674654 264616 674710 264625
rect 674654 264551 674710 264560
rect 674668 263594 674696 264551
rect 674392 263566 674512 263594
rect 674286 262576 674342 262585
rect 674286 262511 674342 262520
rect 674300 243681 674328 262511
rect 674484 253934 674512 263566
rect 674392 253906 674512 253934
rect 674576 263566 674696 263594
rect 674392 244274 674420 253906
rect 674392 244246 674512 244274
rect 674286 243672 674342 243681
rect 674286 243607 674342 243616
rect 674484 242533 674512 244246
rect 674392 242505 674512 242533
rect 674102 241904 674158 241913
rect 674102 241839 674158 241848
rect 674392 241641 674420 242505
rect 674378 241632 674434 241641
rect 674378 241567 674434 241576
rect 673932 239414 674236 239442
rect 673918 236736 673974 236745
rect 673918 236671 673974 236680
rect 673564 234790 673684 234818
rect 673472 234654 673592 234682
rect 673564 229922 673592 234654
rect 673288 229894 673592 229922
rect 673288 227186 673316 229894
rect 673460 229832 673512 229838
rect 673460 229774 673512 229780
rect 673472 229129 673500 229774
rect 673458 229120 673514 229129
rect 673458 229055 673514 229064
rect 673460 228948 673512 228954
rect 673460 228890 673512 228896
rect 673276 227180 673328 227186
rect 673276 227122 673328 227128
rect 673472 227089 673500 228890
rect 673458 227080 673514 227089
rect 673458 227015 673514 227024
rect 673460 226840 673512 226846
rect 673458 226808 673460 226817
rect 673512 226808 673514 226817
rect 673458 226743 673514 226752
rect 673276 226568 673328 226574
rect 673276 226510 673328 226516
rect 673012 224926 673132 224954
rect 673288 224954 673316 226510
rect 673288 224926 673408 224954
rect 673012 215914 673040 224926
rect 673380 224777 673408 224926
rect 673366 224768 673422 224777
rect 673366 224703 673422 224712
rect 673458 224224 673514 224233
rect 673458 224159 673514 224168
rect 673472 216073 673500 224159
rect 673458 216064 673514 216073
rect 673458 215999 673514 216008
rect 673012 215886 673408 215914
rect 673182 215792 673238 215801
rect 673182 215727 673238 215736
rect 673196 212650 673224 215727
rect 673104 212622 673224 212650
rect 673104 201385 673132 212622
rect 673380 212534 673408 215886
rect 673656 215257 673684 234790
rect 673932 233458 673960 236671
rect 674088 234728 674140 234734
rect 674088 234670 674140 234676
rect 674100 234614 674128 234670
rect 674208 234614 674236 239414
rect 674576 235249 674604 263566
rect 681002 263256 681058 263265
rect 681002 263191 681058 263200
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 259622 676260 262783
rect 676036 259616 676088 259622
rect 676036 259558 676088 259564
rect 676220 259616 676272 259622
rect 676220 259558 676272 259564
rect 674746 259312 674802 259321
rect 674746 259247 674802 259256
rect 674760 253934 674788 259247
rect 675298 254960 675354 254969
rect 675298 254895 675354 254904
rect 675022 254688 675078 254697
rect 675022 254623 675078 254632
rect 675036 254402 675064 254623
rect 675036 254374 675248 254402
rect 675024 254312 675076 254318
rect 675024 254254 675076 254260
rect 674668 253906 674788 253934
rect 674668 243085 674696 253906
rect 675036 249914 675064 254254
rect 674852 249886 675064 249914
rect 674852 246378 674880 249886
rect 675022 249248 675078 249257
rect 675022 249183 675078 249192
rect 674852 246350 674972 246378
rect 674668 243057 674788 243085
rect 674760 242758 674788 243057
rect 674748 242752 674800 242758
rect 674748 242694 674800 242700
rect 674944 237538 674972 246350
rect 675036 243085 675064 249183
rect 675220 247398 675248 254374
rect 675312 250526 675340 254895
rect 676048 254697 676076 259558
rect 676218 257136 676274 257145
rect 676218 257071 676274 257080
rect 676232 256465 676260 257071
rect 676218 256456 676274 256465
rect 676218 256391 676274 256400
rect 681016 254969 681044 263191
rect 683026 257544 683082 257553
rect 683026 257479 683082 257488
rect 681002 254960 681058 254969
rect 681002 254895 681058 254904
rect 676034 254688 676090 254697
rect 675852 254652 675904 254658
rect 683040 254658 683068 257479
rect 676034 254623 676090 254632
rect 683028 254652 683080 254658
rect 675852 254594 675904 254600
rect 683028 254594 683080 254600
rect 675864 254402 675892 254594
rect 675496 254374 675892 254402
rect 675496 254318 675524 254374
rect 675484 254312 675536 254318
rect 675484 254254 675536 254260
rect 675496 250889 675524 251056
rect 675482 250880 675538 250889
rect 675482 250815 675538 250824
rect 675312 250498 675418 250526
rect 675758 250200 675814 250209
rect 675758 250135 675814 250144
rect 675772 249900 675800 250135
rect 675390 249520 675446 249529
rect 675390 249455 675446 249464
rect 675404 249220 675432 249455
rect 675220 247370 675418 247398
rect 675298 247208 675354 247217
rect 675298 247143 675354 247152
rect 675312 247058 675340 247143
rect 675312 247030 675432 247058
rect 675206 246936 675262 246945
rect 675206 246871 675262 246880
rect 675220 246213 675248 246871
rect 675404 246840 675432 247030
rect 675220 246185 675418 246213
rect 675206 245576 675262 245585
rect 675262 245534 675418 245562
rect 675206 245511 675262 245520
rect 675206 243672 675262 243681
rect 675206 243607 675262 243616
rect 675220 243085 675248 243607
rect 675036 243057 675156 243085
rect 675220 243057 675418 243085
rect 675128 242533 675156 243057
rect 675300 242752 675352 242758
rect 675300 242694 675352 242700
rect 675036 242505 675156 242533
rect 675312 242533 675340 242694
rect 675312 242505 675418 242533
rect 675036 241514 675064 242505
rect 675758 242312 675814 242321
rect 675758 242247 675814 242256
rect 675772 241876 675800 242247
rect 675036 241486 675248 241514
rect 675220 238218 675248 241486
rect 675404 241097 675432 241231
rect 675390 241088 675446 241097
rect 675390 241023 675446 241032
rect 675390 240272 675446 240281
rect 675390 240207 675446 240216
rect 675404 240040 675432 240207
rect 675220 238190 675418 238218
rect 675312 237646 675432 237674
rect 675312 237538 675340 237646
rect 674944 237510 675340 237538
rect 675404 237524 675432 237646
rect 675128 236354 675418 236382
rect 674562 235240 674618 235249
rect 674562 235175 674618 235184
rect 674838 234696 674894 234705
rect 674838 234631 674894 234640
rect 674100 234586 674144 234614
rect 674208 234586 674328 234614
rect 674116 234258 674144 234586
rect 674104 234252 674156 234258
rect 674104 234194 674156 234200
rect 674102 233880 674158 233889
rect 674102 233815 674104 233824
rect 674156 233815 674158 233824
rect 674104 233786 674156 233792
rect 673932 233430 674052 233458
rect 674024 229786 674052 233430
rect 673748 229758 674052 229786
rect 673748 224954 673776 229758
rect 673920 229628 673972 229634
rect 673920 229570 673972 229576
rect 673748 224926 673868 224954
rect 673642 215248 673698 215257
rect 673642 215183 673698 215192
rect 673642 214976 673698 214985
rect 673642 214911 673698 214920
rect 673288 212506 673408 212534
rect 673090 201376 673146 201385
rect 673090 201311 673146 201320
rect 673288 200114 673316 212506
rect 673656 200569 673684 214911
rect 673642 200560 673698 200569
rect 673642 200495 673698 200504
rect 673840 200114 673868 224926
rect 673932 214010 673960 229570
rect 674104 229356 674156 229362
rect 674104 229298 674156 229304
rect 674116 228585 674144 229298
rect 674102 228576 674158 228585
rect 674102 228511 674158 228520
rect 674102 226808 674158 226817
rect 674102 226743 674158 226752
rect 674116 217410 674144 226743
rect 674300 224954 674328 234586
rect 674852 234546 674880 234631
rect 674852 234518 674972 234546
rect 675128 234530 675156 236354
rect 675850 235240 675906 235249
rect 675850 235175 675906 235184
rect 674944 234410 674972 234518
rect 675116 234524 675168 234530
rect 675116 234466 675168 234472
rect 674944 234382 675432 234410
rect 674932 231668 674984 231674
rect 674932 231610 674984 231616
rect 674944 231146 674972 231610
rect 675116 231396 675168 231402
rect 675116 231338 675168 231344
rect 674944 231118 674996 231146
rect 674968 230858 674996 231118
rect 675128 231062 675156 231338
rect 675116 231056 675168 231062
rect 675116 230998 675168 231004
rect 674956 230852 675008 230858
rect 674956 230794 675008 230800
rect 674674 230480 674730 230489
rect 674674 230415 674676 230424
rect 674728 230415 674730 230424
rect 674838 230480 674894 230489
rect 674838 230415 674894 230424
rect 674676 230386 674728 230392
rect 674852 230330 674880 230415
rect 674576 230302 674880 230330
rect 674576 230246 674604 230302
rect 674564 230240 674616 230246
rect 674564 230182 674616 230188
rect 674452 229968 674504 229974
rect 674452 229910 674504 229916
rect 674464 229650 674492 229910
rect 674464 229622 674512 229650
rect 674484 229401 674512 229622
rect 674470 229392 674526 229401
rect 674470 229327 674526 229336
rect 674838 226128 674894 226137
rect 674838 226063 674894 226072
rect 674300 224926 674420 224954
rect 674392 222329 674420 224926
rect 674378 222320 674434 222329
rect 674378 222255 674434 222264
rect 674852 221513 674880 226063
rect 675022 225856 675078 225865
rect 675022 225791 675078 225800
rect 674838 221504 674894 221513
rect 674838 221439 674894 221448
rect 675036 220561 675064 225791
rect 675206 225312 675262 225321
rect 675206 225247 675262 225256
rect 675022 220552 675078 220561
rect 675022 220487 675078 220496
rect 675220 218770 675248 225247
rect 675404 225162 675432 234382
rect 675864 233986 675892 235175
rect 675852 233980 675904 233986
rect 675852 233922 675904 233928
rect 683396 233980 683448 233986
rect 683396 233922 683448 233928
rect 676034 233880 676090 233889
rect 676034 233815 676036 233824
rect 676088 233815 676090 233824
rect 678244 233844 678296 233850
rect 676036 233786 676088 233792
rect 678244 233786 678296 233792
rect 675852 232552 675904 232558
rect 675850 232520 675852 232529
rect 675904 232520 675906 232529
rect 675850 232455 675906 232464
rect 675850 231568 675906 231577
rect 675850 231503 675852 231512
rect 675904 231503 675906 231512
rect 675852 231474 675904 231480
rect 676678 230480 676734 230489
rect 676678 230415 676734 230424
rect 676034 230208 676090 230217
rect 676034 230143 676090 230152
rect 675128 218742 675248 218770
rect 675312 225134 675432 225162
rect 675128 218657 675156 218742
rect 675114 218648 675170 218657
rect 675114 218583 675170 218592
rect 675022 217832 675078 217841
rect 675022 217767 675078 217776
rect 674116 217382 674236 217410
rect 674208 215370 674236 217382
rect 674654 217016 674710 217025
rect 674654 216951 674710 216960
rect 674378 216336 674434 216345
rect 674378 216271 674434 216280
rect 674392 215529 674420 216271
rect 674378 215520 674434 215529
rect 674378 215455 674434 215464
rect 674208 215342 674328 215370
rect 674102 214024 674158 214033
rect 673932 213982 674102 214010
rect 674102 213959 674158 213968
rect 674010 212800 674066 212809
rect 674010 212735 674066 212744
rect 674024 212534 674052 212735
rect 673196 200086 673316 200114
rect 673748 200086 673868 200114
rect 673932 212506 674052 212534
rect 672906 177712 672962 177721
rect 672906 177647 672962 177656
rect 673196 167929 673224 200086
rect 673366 176896 673422 176905
rect 673366 176831 673422 176840
rect 673182 167920 673238 167929
rect 673182 167855 673238 167864
rect 673090 166968 673146 166977
rect 673090 166903 673146 166912
rect 672906 165608 672962 165617
rect 672906 165543 672962 165552
rect 672722 126032 672778 126041
rect 672722 125967 672778 125976
rect 672722 123992 672778 124001
rect 672722 123927 672778 123936
rect 672736 106593 672764 123927
rect 672920 115841 672948 165543
rect 673104 117609 673132 166903
rect 673380 132161 673408 176831
rect 673748 153377 673776 200086
rect 673932 177313 673960 212506
rect 674102 209672 674158 209681
rect 674102 209607 674158 209616
rect 673918 177304 673974 177313
rect 673918 177239 673974 177248
rect 673918 168736 673974 168745
rect 673918 168671 673974 168680
rect 673734 153368 673790 153377
rect 673734 153303 673790 153312
rect 673932 151065 673960 168671
rect 673918 151056 673974 151065
rect 673918 150991 673974 151000
rect 673366 132152 673422 132161
rect 673366 132087 673422 132096
rect 673734 123584 673790 123593
rect 673734 123519 673790 123528
rect 673550 123176 673606 123185
rect 673550 123111 673606 123120
rect 673366 120728 673422 120737
rect 673366 120663 673422 120672
rect 673090 117600 673146 117609
rect 673090 117535 673146 117544
rect 672906 115832 672962 115841
rect 672906 115767 672962 115776
rect 672722 106584 672778 106593
rect 672722 106519 672778 106528
rect 672354 106176 672410 106185
rect 672354 106111 672410 106120
rect 673380 104553 673408 120663
rect 673564 117065 673592 123111
rect 673550 117056 673606 117065
rect 673550 116991 673606 117000
rect 673748 105822 673776 123519
rect 674116 120465 674144 209607
rect 674300 178129 674328 215342
rect 674668 215294 674696 216951
rect 674838 216200 674894 216209
rect 674838 216135 674894 216144
rect 674668 215266 674788 215294
rect 674470 214160 674526 214169
rect 674470 214095 674526 214104
rect 674484 200841 674512 214095
rect 674470 200832 674526 200841
rect 674470 200767 674526 200776
rect 674760 191162 674788 215266
rect 674852 201634 674880 216135
rect 675036 205634 675064 217767
rect 675312 205889 675340 225134
rect 676048 221513 676076 230143
rect 676402 228576 676458 228585
rect 676402 228511 676458 228520
rect 676034 221504 676090 221513
rect 676034 221439 676090 221448
rect 676034 219056 676090 219065
rect 676090 219014 676260 219042
rect 676034 218991 676090 219000
rect 676232 218074 676260 219014
rect 676220 218068 676272 218074
rect 676220 218010 676272 218016
rect 675852 217592 675904 217598
rect 675574 217560 675630 217569
rect 675630 217540 675852 217546
rect 675630 217534 675904 217540
rect 675630 217518 675892 217534
rect 675574 217495 675630 217504
rect 675944 215552 675996 215558
rect 675942 215520 675944 215529
rect 675996 215520 675998 215529
rect 675942 215455 675998 215464
rect 676416 215294 676444 228511
rect 676692 217598 676720 230415
rect 677046 227080 677102 227089
rect 677046 227015 677102 227024
rect 676864 218068 676916 218074
rect 676864 218010 676916 218016
rect 676680 217592 676732 217598
rect 676680 217534 676732 217540
rect 676232 215266 676444 215294
rect 675942 214704 675998 214713
rect 676232 214690 676260 215266
rect 675998 214662 676260 214690
rect 675942 214639 675998 214648
rect 675850 212120 675906 212129
rect 675850 212055 675906 212064
rect 675864 209681 675892 212055
rect 675850 209672 675906 209681
rect 675850 209607 675906 209616
rect 676876 206961 676904 218010
rect 677060 215558 677088 227015
rect 678256 223825 678284 233786
rect 683212 232552 683264 232558
rect 683212 232494 683264 232500
rect 678242 223816 678298 223825
rect 678242 223751 678298 223760
rect 683224 222737 683252 232494
rect 683210 222728 683266 222737
rect 683210 222663 683266 222672
rect 683408 219881 683436 233922
rect 683580 231532 683632 231538
rect 683580 231474 683632 231480
rect 683592 223145 683620 231474
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683578 223136 683634 223145
rect 683578 223071 683634 223080
rect 683394 219872 683450 219881
rect 683394 219807 683450 219816
rect 683302 218648 683358 218657
rect 683302 218583 683358 218592
rect 677048 215552 677100 215558
rect 677048 215494 677100 215500
rect 683118 212936 683174 212945
rect 683118 212871 683174 212880
rect 678978 211440 679034 211449
rect 678978 211375 679034 211384
rect 678992 207641 679020 211375
rect 683132 211206 683160 212871
rect 680360 211200 680412 211206
rect 680360 211142 680412 211148
rect 683120 211200 683172 211206
rect 683120 211142 683172 211148
rect 680372 210633 680400 211142
rect 680358 210624 680414 210633
rect 680358 210559 680414 210568
rect 683316 210361 683344 218583
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 678978 207632 679034 207641
rect 678978 207567 679034 207576
rect 676862 206952 676918 206961
rect 676862 206887 676918 206896
rect 675312 205861 675418 205889
rect 674944 205606 675064 205634
rect 674944 202209 674972 205606
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675128 204666 675418 204694
rect 675128 204513 675156 204666
rect 675114 204504 675170 204513
rect 675114 204439 675170 204448
rect 675758 204232 675814 204241
rect 675758 204167 675814 204176
rect 675772 204035 675800 204167
rect 674944 202181 675418 202209
rect 675312 201742 675432 201770
rect 675312 201634 675340 201742
rect 674852 201606 675340 201634
rect 675404 201620 675432 201742
rect 675114 201376 675170 201385
rect 675114 201311 675170 201320
rect 675128 201022 675156 201311
rect 675128 200994 675418 201022
rect 675298 200832 675354 200841
rect 675298 200767 675354 200776
rect 675114 200560 675170 200569
rect 675114 200495 675170 200504
rect 675128 196670 675156 200495
rect 675312 197282 675340 200767
rect 675758 200696 675814 200705
rect 675758 200631 675814 200640
rect 675772 200328 675800 200631
rect 675758 198384 675814 198393
rect 675758 198319 675814 198328
rect 675772 197880 675800 198319
rect 675404 197282 675432 197336
rect 675312 197254 675432 197282
rect 675312 196710 675432 196738
rect 675312 196670 675340 196710
rect 675128 196642 675340 196670
rect 675404 196656 675432 196710
rect 675114 196344 675170 196353
rect 675114 196279 675170 196288
rect 675128 196058 675156 196279
rect 675128 196030 675418 196058
rect 675298 195800 675354 195809
rect 675298 195735 675354 195744
rect 675312 194834 675340 195735
rect 675312 194806 675418 194834
rect 675114 193216 675170 193225
rect 675114 193151 675170 193160
rect 675128 192998 675156 193151
rect 675128 192970 675418 192998
rect 675666 192672 675722 192681
rect 675666 192607 675722 192616
rect 675680 192372 675708 192607
rect 674760 191134 675418 191162
rect 676862 189680 676918 189689
rect 676862 189615 676918 189624
rect 674286 178120 674342 178129
rect 674286 178055 674342 178064
rect 674654 175264 674710 175273
rect 674654 175199 674710 175208
rect 674378 174448 674434 174457
rect 674378 174383 674434 174392
rect 674392 129713 674420 174383
rect 674668 130529 674696 175199
rect 675206 174040 675262 174049
rect 675206 173975 675262 173984
rect 674838 169416 674894 169425
rect 674838 169351 674894 169360
rect 674852 160585 674880 169351
rect 675220 164234 675248 173975
rect 676034 173224 676090 173233
rect 676090 173182 676260 173210
rect 676034 173159 676090 173168
rect 675390 171184 675446 171193
rect 675390 171119 675446 171128
rect 675404 166994 675432 171119
rect 675942 169416 675998 169425
rect 676232 169402 676260 173182
rect 676586 169960 676642 169969
rect 676586 169895 676642 169904
rect 675998 169374 676260 169402
rect 675942 169351 675998 169360
rect 675850 167920 675906 167929
rect 675850 167855 675906 167864
rect 675036 164206 675248 164234
rect 675312 166966 675432 166994
rect 675864 166977 675892 167855
rect 676034 167104 676090 167113
rect 676034 167039 676090 167048
rect 675850 166968 675906 166977
rect 674838 160576 674894 160585
rect 674838 160511 674894 160520
rect 675036 159497 675064 164206
rect 675312 161650 675340 166966
rect 675850 166903 675906 166912
rect 676048 165617 676076 167039
rect 676600 166433 676628 169895
rect 676876 166433 676904 189615
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 678242 171592 678298 171601
rect 678242 171527 678298 171536
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676862 166424 676918 166433
rect 676862 166359 676918 166368
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 678256 162858 678284 171527
rect 675852 162852 675904 162858
rect 675220 161622 675340 161650
rect 675404 162812 675852 162840
rect 675220 159610 675248 161622
rect 675404 161474 675432 162812
rect 675852 162794 675904 162800
rect 678244 162852 678296 162858
rect 678244 162794 678296 162800
rect 675312 161446 675432 161474
rect 675312 160154 675340 161446
rect 675482 161392 675538 161401
rect 675482 161327 675538 161336
rect 675496 160888 675524 161327
rect 675482 160576 675538 160585
rect 675482 160511 675538 160520
rect 675496 160344 675524 160511
rect 675312 160126 675432 160154
rect 675404 159664 675432 160126
rect 675220 159582 675340 159610
rect 675022 159488 675078 159497
rect 675022 159423 675078 159432
rect 675312 156657 675340 159582
rect 675482 159488 675538 159497
rect 675482 159423 675538 159432
rect 675496 159052 675524 159423
rect 675772 157049 675800 157216
rect 675758 157040 675814 157049
rect 675758 156975 675814 156984
rect 675312 156629 675418 156657
rect 675128 155978 675418 156006
rect 675128 154465 675156 155978
rect 675758 155680 675814 155689
rect 675758 155615 675814 155624
rect 675772 155380 675800 155615
rect 675114 154456 675170 154465
rect 675114 154391 675170 154400
rect 675114 153096 675170 153105
rect 675114 153031 675170 153040
rect 675666 153096 675722 153105
rect 675666 153031 675722 153040
rect 675128 152334 675156 153031
rect 675680 152864 675708 153031
rect 675128 152306 675418 152334
rect 675772 151473 675800 151675
rect 675758 151464 675814 151473
rect 675758 151399 675814 151408
rect 675114 151056 675170 151065
rect 675170 151014 675418 151042
rect 675114 150991 675170 151000
rect 675128 149821 675418 149849
rect 675128 147665 675156 149821
rect 675298 149016 675354 149025
rect 675298 148951 675354 148960
rect 675114 147656 675170 147665
rect 675114 147591 675170 147600
rect 675312 146690 675340 148951
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675312 146662 675432 146690
rect 675404 146132 675432 146662
rect 676034 134600 676090 134609
rect 676034 134535 676090 134544
rect 676048 132569 676076 134535
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676034 132560 676090 132569
rect 676034 132495 676090 132504
rect 674654 130520 674710 130529
rect 674654 130455 674710 130464
rect 676218 130248 676274 130257
rect 676218 130183 676274 130192
rect 674378 129704 674434 129713
rect 674378 129639 674434 129648
rect 674286 129296 674342 129305
rect 674286 129231 674342 129240
rect 674102 120456 674158 120465
rect 674102 120391 674158 120400
rect 674300 120057 674328 129231
rect 675206 128888 675262 128897
rect 675206 128823 675262 128832
rect 674470 125624 674526 125633
rect 674470 125559 674526 125568
rect 674286 120048 674342 120057
rect 674286 119983 674342 119992
rect 674484 111353 674512 125559
rect 674654 124808 674710 124817
rect 674654 124743 674710 124752
rect 674470 111344 674526 111353
rect 674470 111279 674526 111288
rect 674668 106434 674696 124743
rect 675220 118694 675248 128823
rect 676232 127809 676260 130183
rect 676678 128208 676734 128217
rect 676678 128143 676734 128152
rect 676218 127800 676274 127809
rect 676218 127735 676274 127744
rect 676402 127800 676458 127809
rect 676402 127735 676458 127744
rect 675942 125352 675998 125361
rect 675942 125287 675944 125296
rect 675996 125287 675998 125296
rect 676126 125352 676182 125361
rect 676126 125287 676182 125296
rect 675944 125258 675996 125264
rect 675852 123412 675904 123418
rect 675852 123354 675904 123360
rect 674852 118666 675248 118694
rect 674852 114345 674880 118666
rect 675864 118561 675892 123354
rect 676140 120737 676168 125287
rect 676416 123418 676444 127735
rect 676692 126177 676720 128143
rect 676678 126168 676734 126177
rect 676678 126103 676734 126112
rect 683118 126168 683174 126177
rect 683118 126103 683174 126112
rect 676862 125760 676918 125769
rect 676862 125695 676918 125704
rect 676586 125352 676642 125361
rect 676586 125287 676588 125296
rect 676640 125287 676642 125296
rect 676588 125258 676640 125264
rect 676404 123412 676456 123418
rect 676404 123354 676456 123360
rect 676126 120728 676182 120737
rect 676126 120663 676182 120672
rect 675298 118552 675354 118561
rect 675298 118487 675354 118496
rect 675850 118552 675906 118561
rect 675850 118487 675906 118496
rect 675022 116376 675078 116385
rect 675022 116311 675078 116320
rect 675036 115934 675064 116311
rect 675036 115906 675156 115934
rect 674838 114336 674894 114345
rect 674838 114271 674894 114280
rect 675128 111466 675156 115906
rect 675312 115138 675340 118487
rect 676876 116550 676904 125695
rect 678978 125352 679034 125361
rect 678978 125287 679034 125296
rect 677598 122088 677654 122097
rect 677598 122023 677654 122032
rect 675852 116544 675904 116550
rect 675852 116486 675904 116492
rect 676864 116544 676916 116550
rect 676864 116486 676916 116492
rect 675864 116385 675892 116486
rect 675850 116376 675906 116385
rect 675850 116311 675906 116320
rect 677612 116113 677640 122023
rect 678992 121689 679020 125287
rect 683132 122913 683160 126103
rect 683118 122904 683174 122913
rect 683118 122839 683174 122848
rect 678978 121680 679034 121689
rect 678978 121615 679034 121624
rect 675482 116104 675538 116113
rect 675482 116039 675538 116048
rect 677598 116104 677654 116113
rect 677598 116039 677654 116048
rect 675496 115668 675524 116039
rect 675312 115110 675418 115138
rect 675772 114345 675800 114479
rect 675390 114336 675446 114345
rect 675390 114271 675446 114280
rect 675758 114336 675814 114345
rect 675758 114271 675814 114280
rect 675404 113832 675432 114271
rect 675758 112432 675814 112441
rect 675758 112367 675814 112376
rect 675772 111996 675800 112367
rect 675128 111438 675418 111466
rect 675390 111344 675446 111353
rect 675390 111279 675446 111288
rect 675404 110772 675432 111279
rect 675758 110392 675814 110401
rect 675758 110327 675814 110336
rect 675772 110160 675800 110327
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106593 675156 107086
rect 675114 106584 675170 106593
rect 675114 106519 675170 106528
rect 675312 106474 675418 106502
rect 675312 106434 675340 106474
rect 674668 106406 675340 106434
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 673748 105794 675340 105822
rect 675404 105808 675432 105862
rect 675128 104638 675340 104666
rect 675128 104553 675156 104638
rect 673366 104544 673422 104553
rect 673366 104479 673422 104488
rect 675114 104544 675170 104553
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 675114 104479 675170 104488
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 675666 102640 675722 102649
rect 675666 102575 675722 102584
rect 675680 102136 675708 102575
rect 675404 100450 675432 100980
rect 675312 100422 675432 100450
rect 675312 99385 675340 100422
rect 671986 99376 672042 99385
rect 671986 99311 672042 99320
rect 675298 99376 675354 99385
rect 675298 99311 675354 99320
rect 668216 76560 668268 76566
rect 668216 76502 668268 76508
rect 666560 75200 666612 75206
rect 666560 75142 666612 75148
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661776 46504 661828 46510
rect 661776 46446 661828 46452
rect 661420 45526 661632 45554
rect 464710 44568 464766 44577
rect 464710 44503 464766 44512
rect 463882 44160 463938 44169
rect 463882 44095 463938 44104
rect 471058 43888 471114 43897
rect 471058 43823 471114 43832
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 463974 42936 464030 42945
rect 463974 42871 464030 42880
rect 463988 42514 464016 42871
rect 463988 42486 464050 42514
rect 463056 42356 463108 42362
rect 463056 42298 463108 42304
rect 464022 42228 464050 42486
rect 465828 42364 465856 43143
rect 471072 42106 471100 43823
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42228 518848 42735
rect 661420 42187 661448 45526
rect 661408 42181 661460 42187
rect 515402 42120 515458 42129
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 661408 42123 661460 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 461950 41848 462006 41857
rect 461950 41783 462006 41792
rect 459192 41744 459244 41750
rect 459192 41686 459244 41692
rect 458178 41168 458234 41177
rect 458178 41103 458234 41112
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 676034 897116 676090 897152
rect 676034 897096 676036 897116
rect 676036 897096 676088 897116
rect 676088 897096 676090 897116
rect 651470 868536 651526 868592
rect 675850 896688 675906 896744
rect 676034 896280 676090 896336
rect 652022 867584 652078 867640
rect 651470 866224 651526 866280
rect 651378 865172 651380 865192
rect 651380 865172 651432 865192
rect 651432 865172 651434 865192
rect 651378 865136 651434 865172
rect 651470 863812 651472 863832
rect 651472 863812 651524 863832
rect 651524 863812 651526 863832
rect 651470 863776 651526 863812
rect 651470 862280 651526 862336
rect 35622 817944 35678 818000
rect 35806 817264 35862 817320
rect 35622 816856 35678 816912
rect 35806 816040 35862 816096
rect 35622 815224 35678 815280
rect 35806 814408 35862 814464
rect 41326 813592 41382 813648
rect 41142 812776 41198 812832
rect 40498 812368 40554 812424
rect 39302 811552 39358 811608
rect 33046 811144 33102 811200
rect 31022 809920 31078 809976
rect 31758 806676 31814 806712
rect 31758 806656 31760 806676
rect 31760 806656 31812 806676
rect 31812 806656 31814 806676
rect 33782 809512 33838 809568
rect 40682 809104 40738 809160
rect 40498 805568 40554 805624
rect 40130 800808 40186 800864
rect 40958 808288 41014 808344
rect 41142 807880 41198 807936
rect 41326 806248 41382 806304
rect 41786 810736 41842 810792
rect 41970 810328 42026 810384
rect 41786 808696 41842 808752
rect 41786 805160 41842 805216
rect 41970 804888 42026 804944
rect 41602 804616 41658 804672
rect 40682 800536 40738 800592
rect 41970 800264 42026 800320
rect 42890 807472 42946 807528
rect 42154 797272 42210 797328
rect 41786 796184 41842 796240
rect 41786 794416 41842 794472
rect 42062 792920 42118 792976
rect 42246 791288 42302 791344
rect 41786 790608 41842 790664
rect 42614 791560 42670 791616
rect 42246 788160 42302 788216
rect 41786 786800 41842 786856
rect 41786 786120 41842 786176
rect 40498 776600 40554 776656
rect 35806 774696 35862 774752
rect 35162 773880 35218 773936
rect 35346 773472 35402 773528
rect 35530 773100 35532 773120
rect 35532 773100 35584 773120
rect 35584 773100 35586 773120
rect 35530 773064 35586 773100
rect 35806 773064 35862 773120
rect 40498 773100 40500 773120
rect 40500 773100 40552 773120
rect 40552 773100 40554 773120
rect 40498 773064 40554 773100
rect 35622 772248 35678 772304
rect 41326 772248 41382 772304
rect 35806 771860 35862 771896
rect 35806 771840 35808 771860
rect 35808 771840 35860 771860
rect 35860 771840 35862 771860
rect 35806 771452 35862 771488
rect 35806 771432 35808 771452
rect 35808 771432 35860 771452
rect 35860 771432 35862 771452
rect 39578 771432 39634 771488
rect 35622 771024 35678 771080
rect 35806 770616 35862 770672
rect 40038 770616 40094 770672
rect 35806 770208 35862 770264
rect 35346 769392 35402 769448
rect 35530 768984 35586 769040
rect 35806 769004 35862 769040
rect 35806 768984 35808 769004
rect 35808 768984 35860 769004
rect 35860 768984 35862 769004
rect 39762 768576 39818 768632
rect 35622 768168 35678 768224
rect 33046 767760 33102 767816
rect 35806 767760 35862 767816
rect 35162 766944 35218 767000
rect 35806 766536 35862 766592
rect 35806 765720 35862 765776
rect 35806 764532 35808 764552
rect 35808 764532 35860 764552
rect 35860 764532 35862 764552
rect 35806 764496 35862 764532
rect 35806 764088 35862 764144
rect 35806 762864 35862 762920
rect 40314 766944 40370 767000
rect 39302 764496 39358 764552
rect 40406 764088 40462 764144
rect 37094 763700 37150 763736
rect 37094 763680 37096 763700
rect 37096 763680 37148 763700
rect 37148 763680 37150 763700
rect 36542 759056 36598 759112
rect 40498 759500 40500 759520
rect 40500 759500 40552 759520
rect 40552 759500 40554 759520
rect 40498 759464 40554 759500
rect 41694 763680 41750 763736
rect 41694 763292 41750 763328
rect 41694 763272 41696 763292
rect 41696 763272 41748 763292
rect 41748 763272 41750 763292
rect 42706 768576 42762 768632
rect 42430 759464 42486 759520
rect 42154 758920 42210 758976
rect 40682 757696 40738 757752
rect 39946 757424 40002 757480
rect 41786 757016 41842 757072
rect 41878 755384 41934 755440
rect 42154 754840 42210 754896
rect 42062 754024 42118 754080
rect 42062 752936 42118 752992
rect 42062 751712 42118 751768
rect 41786 750352 41842 750408
rect 42338 749536 42394 749592
rect 41786 746680 41842 746736
rect 42062 744776 42118 744832
rect 41786 743688 41842 743744
rect 42522 745048 42578 745104
rect 39578 732264 39634 732320
rect 35806 731312 35862 731368
rect 35622 730904 35678 730960
rect 35438 730496 35494 730552
rect 35254 729680 35310 729736
rect 35806 730088 35862 730144
rect 35622 729272 35678 729328
rect 35806 728864 35862 728920
rect 39946 731992 40002 732048
rect 40406 731584 40462 731640
rect 35622 728456 35678 728512
rect 35806 728048 35862 728104
rect 35806 727640 35862 727696
rect 41694 730260 41696 730280
rect 41696 730260 41748 730280
rect 41748 730260 41750 730280
rect 41694 730224 41750 730260
rect 41694 728628 41696 728648
rect 41696 728628 41748 728648
rect 41748 728628 41750 728648
rect 41694 728592 41750 728628
rect 35806 727268 35808 727288
rect 35808 727268 35860 727288
rect 35860 727268 35862 727288
rect 35806 727232 35862 727268
rect 41694 726960 41750 727016
rect 41142 726824 41198 726880
rect 39302 726178 39358 726234
rect 35162 724784 35218 724840
rect 31666 724376 31722 724432
rect 33046 723968 33102 724024
rect 31666 718256 31722 718312
rect 33782 723152 33838 723208
rect 41326 726232 41382 726234
rect 41326 726180 41328 726232
rect 41328 726180 41380 726232
rect 41380 726180 41382 726232
rect 41326 726178 41382 726180
rect 41786 725736 41842 725792
rect 41326 725600 41382 725656
rect 41142 725192 41198 725248
rect 41326 720296 41382 720352
rect 41142 719208 41198 719264
rect 41970 722336 42026 722392
rect 41786 721928 41842 721984
rect 41510 718936 41566 718992
rect 41786 718528 41842 718584
rect 41970 717984 42026 718040
rect 39302 716080 39358 716136
rect 39854 715556 39910 715592
rect 39854 715536 39856 715556
rect 39856 715536 39908 715556
rect 39908 715536 39910 715556
rect 37738 714448 37794 714504
rect 42614 719208 42670 719264
rect 42614 718936 42670 718992
rect 42430 715536 42486 715592
rect 42062 714448 42118 714504
rect 41234 714176 41290 714232
rect 41786 712136 41842 712192
rect 42154 710776 42210 710832
rect 42062 708464 42118 708520
rect 42062 707648 42118 707704
rect 41786 707376 41842 707432
rect 42246 706152 42302 706208
rect 42062 703432 42118 703488
rect 42338 701800 42394 701856
rect 41786 700440 41842 700496
rect 42706 702072 42762 702128
rect 42706 688064 42762 688120
rect 40866 686840 40922 686896
rect 41142 686432 41198 686488
rect 41050 685854 41106 685910
rect 40866 684800 40922 684856
rect 41694 684700 41696 684720
rect 41696 684700 41748 684720
rect 41748 684700 41750 684720
rect 41694 684664 41750 684700
rect 41326 683460 41382 683462
rect 41326 683408 41328 683460
rect 41328 683408 41380 683460
rect 41380 683408 41382 683460
rect 41326 683406 41382 683408
rect 40958 682760 41014 682816
rect 35162 681944 35218 682000
rect 32402 681128 32458 681184
rect 33782 680720 33838 680776
rect 42522 682352 42578 682408
rect 42246 681536 42302 681592
rect 41142 679904 41198 679960
rect 41786 678816 41842 678872
rect 41786 678272 41842 678328
rect 40958 677748 41014 677750
rect 40958 677696 40960 677748
rect 40960 677696 41012 677748
rect 41012 677696 41014 677748
rect 40958 677694 41014 677696
rect 39946 677048 40002 677104
rect 43074 771432 43130 771488
rect 43442 797272 43498 797328
rect 43258 770616 43314 770672
rect 43626 764088 43682 764144
rect 43258 757424 43314 757480
rect 43074 732264 43130 732320
rect 43074 686024 43130 686080
rect 43074 677864 43130 677920
rect 39946 672968 40002 673024
rect 32402 672696 32458 672752
rect 38934 671200 38990 671256
rect 38198 670928 38254 670984
rect 41786 669024 41842 669080
rect 43442 752936 43498 752992
rect 43442 723560 43498 723616
rect 43626 710776 43682 710832
rect 43626 707648 43682 707704
rect 43442 703432 43498 703488
rect 43442 687248 43498 687304
rect 43626 680312 43682 680368
rect 43442 676640 43498 676696
rect 43258 671880 43314 671936
rect 42798 671200 42854 671256
rect 42154 666576 42210 666632
rect 42062 665896 42118 665952
rect 42430 665488 42486 665544
rect 42246 665216 42302 665272
rect 41786 663992 41842 664048
rect 42062 662768 42118 662824
rect 42706 660864 42762 660920
rect 41786 658280 41842 658336
rect 42522 658552 42578 658608
rect 35806 644680 35862 644736
rect 40130 644680 40186 644736
rect 38566 644272 38622 644328
rect 35346 643864 35402 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 35622 642640 35678 642696
rect 39946 643048 40002 643104
rect 35806 642232 35862 642288
rect 35438 641416 35494 641472
rect 35806 641008 35862 641064
rect 39762 641008 39818 641064
rect 35622 640600 35678 640656
rect 40038 640192 40094 640248
rect 35806 639784 35862 639840
rect 35806 638988 35862 639024
rect 35806 638968 35808 638988
rect 35808 638968 35860 638988
rect 35860 638968 35862 638988
rect 35622 638560 35678 638616
rect 35162 637744 35218 637800
rect 31942 636928 31998 636984
rect 35806 638152 35862 638208
rect 35530 636540 35586 636576
rect 35530 636520 35532 636540
rect 35532 636520 35584 636540
rect 35584 636520 35586 636540
rect 35806 636520 35862 636576
rect 35806 635704 35862 635760
rect 35622 634480 35678 634536
rect 35806 633700 35808 633720
rect 35808 633700 35860 633720
rect 35860 633700 35862 633720
rect 35806 633664 35862 633700
rect 40682 636520 40738 636576
rect 39854 636112 39910 636168
rect 38566 633664 38622 633720
rect 37922 631352 37978 631408
rect 35162 629856 35218 629912
rect 42706 636520 42762 636576
rect 41602 634924 41604 634944
rect 41604 634924 41656 634944
rect 41656 634924 41658 634944
rect 41602 634888 41658 634924
rect 41418 632848 41474 632904
rect 40130 631896 40186 631952
rect 42614 631352 42670 631408
rect 39578 630672 39634 630728
rect 40222 629176 40278 629232
rect 40498 628260 40500 628280
rect 40500 628260 40552 628280
rect 40552 628260 40554 628280
rect 40498 628224 40554 628260
rect 42154 629176 42210 629232
rect 42338 628258 42394 628314
rect 42246 625640 42302 625696
rect 42062 623736 42118 623792
rect 42062 623328 42118 623384
rect 42062 622104 42118 622160
rect 41786 620880 41842 620936
rect 42706 624552 42762 624608
rect 42522 619792 42578 619848
rect 41786 616392 41842 616448
rect 42614 616120 42670 616176
rect 42338 615712 42394 615768
rect 42614 615168 42670 615224
rect 43258 666512 43314 666568
rect 42890 613808 42946 613864
rect 43258 612176 43314 612232
rect 43626 631896 43682 631952
rect 44270 772248 44326 772304
rect 62210 790472 62266 790528
rect 62118 789148 62120 789168
rect 62120 789148 62172 789168
rect 62172 789148 62174 789168
rect 62118 789112 62174 789148
rect 62118 787344 62174 787400
rect 62762 787072 62818 787128
rect 61382 786120 61438 786176
rect 62118 784896 62174 784952
rect 651470 778368 651526 778424
rect 652022 777008 652078 777064
rect 45006 776600 45062 776656
rect 651470 776056 651526 776112
rect 651378 775276 651380 775296
rect 651380 775276 651432 775296
rect 651432 775276 651434 775296
rect 651378 775240 651434 775276
rect 44914 773064 44970 773120
rect 44546 766944 44602 767000
rect 44730 754024 44786 754080
rect 45098 764496 45154 764552
rect 45282 763680 45338 763736
rect 45558 763272 45614 763328
rect 45098 751712 45154 751768
rect 44914 731992 44970 732048
rect 44546 731584 44602 731640
rect 45190 728592 45246 728648
rect 44270 726960 44326 727016
rect 44454 722744 44510 722800
rect 44638 721520 44694 721576
rect 44454 708464 44510 708520
rect 44822 687656 44878 687712
rect 44270 685208 44326 685264
rect 44454 684664 44510 684720
rect 44270 683984 44326 684040
rect 43994 679496 44050 679552
rect 44454 644680 44510 644736
rect 45006 684392 45062 684448
rect 45006 667392 45062 667448
rect 44730 643048 44786 643104
rect 44270 641008 44326 641064
rect 43994 636112 44050 636168
rect 44362 634888 44418 634944
rect 45098 640192 45154 640248
rect 43994 623328 44050 623384
rect 44178 622104 44234 622160
rect 44086 613808 44142 613864
rect 43764 612196 43820 612232
rect 43764 612176 43766 612196
rect 43766 612176 43818 612196
rect 43818 612176 43820 612196
rect 44086 612060 44142 612096
rect 44086 612040 44088 612060
rect 44088 612040 44140 612060
rect 44140 612040 44142 612060
rect 43994 611788 44050 611824
rect 43994 611768 43996 611788
rect 43996 611768 44048 611788
rect 44048 611768 44050 611788
rect 44086 611532 44088 611552
rect 44088 611532 44140 611552
rect 44140 611532 44142 611552
rect 44086 611496 44142 611532
rect 35806 601724 35862 601760
rect 35806 601704 35808 601724
rect 35808 601704 35860 601724
rect 35860 601704 35862 601724
rect 33046 595346 33102 595402
rect 35438 595346 35494 595402
rect 31022 594360 31078 594416
rect 33782 593544 33838 593600
rect 38566 601296 38622 601352
rect 39946 600888 40002 600944
rect 44914 630672 44970 630728
rect 44638 600480 44694 600536
rect 44914 600072 44970 600128
rect 42982 597624 43038 597680
rect 42614 596808 42670 596864
rect 42338 595992 42394 596048
rect 41694 595756 41696 595776
rect 41696 595756 41748 595776
rect 41748 595756 41750 595776
rect 41694 595720 41750 595756
rect 39302 594768 39358 594824
rect 41786 594224 41842 594280
rect 41694 592900 41696 592920
rect 41696 592900 41748 592920
rect 41748 592900 41750 592920
rect 41694 592864 41750 592900
rect 41234 589600 41290 589656
rect 40682 587308 40738 587344
rect 40682 587288 40684 587308
rect 40684 587288 40736 587308
rect 40736 587288 40738 587308
rect 40130 585948 40186 585984
rect 40130 585928 40132 585948
rect 40132 585928 40184 585948
rect 40184 585928 40186 585948
rect 41234 585792 41290 585848
rect 39302 585112 39358 585168
rect 40590 584568 40646 584624
rect 42154 585792 42210 585848
rect 42614 587560 42670 587616
rect 42706 587288 42762 587344
rect 42706 584568 42762 584624
rect 42154 581848 42210 581904
rect 42154 580624 42210 580680
rect 41786 580216 41842 580272
rect 42062 578720 42118 578776
rect 42246 578448 42302 578504
rect 42062 578040 42118 578096
rect 41786 577768 41842 577824
rect 42246 575592 42302 575648
rect 41786 574640 41842 574696
rect 42614 572736 42670 572792
rect 42062 571512 42118 571568
rect 42430 571376 42486 571432
rect 41786 570152 41842 570208
rect 43166 596944 43222 597000
rect 44362 593136 44418 593192
rect 44178 591912 44234 591968
rect 43350 591504 43406 591560
rect 43626 590280 43682 590336
rect 42338 558048 42394 558104
rect 40038 553352 40094 553408
rect 40958 553352 41014 553408
rect 34426 551928 34482 551984
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 43074 556416 43130 556472
rect 42798 554784 42854 554840
rect 42338 552608 42394 552664
rect 42982 552336 43038 552392
rect 42798 551112 42854 551168
rect 41878 550296 41934 550352
rect 41326 546352 41382 546408
rect 42062 549888 42118 549944
rect 41878 545672 41934 545728
rect 42062 545400 42118 545456
rect 41326 541320 41382 541376
rect 41786 540640 41842 540696
rect 42522 539552 42578 539608
rect 42614 538056 42670 538112
rect 43166 549480 43222 549536
rect 42430 537376 42486 537432
rect 41786 536968 41842 537024
rect 42246 536424 42302 536480
rect 42062 535608 42118 535664
rect 42706 532752 42762 532808
rect 42614 530712 42670 530768
rect 42430 529488 42486 529544
rect 41786 528944 41842 529000
rect 42246 528808 42302 528864
rect 42614 527176 42670 527232
rect 35806 430072 35862 430128
rect 41970 427080 42026 427136
rect 41326 425992 41382 426048
rect 41142 425584 41198 425640
rect 40958 425176 41014 425232
rect 32034 424360 32090 424416
rect 41878 424224 41934 424280
rect 41142 418784 41198 418840
rect 42798 423544 42854 423600
rect 42522 419872 42578 419928
rect 42062 411848 42118 411904
rect 42522 411848 42578 411904
rect 41786 409400 41842 409456
rect 41970 408040 42026 408096
rect 42430 407768 42486 407824
rect 42246 407496 42302 407552
rect 42062 406680 42118 406736
rect 41786 406272 41842 406328
rect 42246 405592 42302 405648
rect 42430 405592 42486 405648
rect 43258 420688 43314 420744
rect 43074 419464 43130 419520
rect 42338 402872 42394 402928
rect 41786 401784 41842 401840
rect 42430 400152 42486 400208
rect 41786 400016 41842 400072
rect 41786 398792 41842 398848
rect 42154 395664 42210 395720
rect 41142 387096 41198 387152
rect 40774 385872 40830 385928
rect 41326 386688 41382 386744
rect 41326 385872 41382 385928
rect 41326 382608 41382 382664
rect 40958 381792 41014 381848
rect 41142 381792 41198 381848
rect 40222 381384 40278 381440
rect 40774 381384 40830 381440
rect 35162 380976 35218 381032
rect 33782 379752 33838 379808
rect 33782 371864 33838 371920
rect 37922 380160 37978 380216
rect 35806 379344 35862 379400
rect 35806 376488 35862 376544
rect 35806 374584 35862 374640
rect 40958 379752 41014 379808
rect 40590 379344 40646 379400
rect 37922 372680 37978 372736
rect 41786 368464 41842 368520
rect 42890 379344 42946 379400
rect 42062 366152 42118 366208
rect 42062 364792 42118 364848
rect 42246 364112 42302 364168
rect 41786 363704 41842 363760
rect 42890 366152 42946 366208
rect 42246 362888 42302 362944
rect 42706 363160 42762 363216
rect 42430 361528 42486 361584
rect 41786 360032 41842 360088
rect 41786 359216 41842 359272
rect 41786 358672 41842 358728
rect 41786 356088 41842 356144
rect 42430 354320 42486 354376
rect 43074 353912 43130 353968
rect 42154 353232 42210 353288
rect 44178 578720 44234 578776
rect 44638 580624 44694 580680
rect 44362 578040 44418 578096
rect 45098 598848 45154 598904
rect 45098 598440 45154 598496
rect 44914 558728 44970 558784
rect 44546 556824 44602 556880
rect 44270 556008 44326 556064
rect 43810 548256 43866 548312
rect 43994 547032 44050 547088
rect 43810 355136 43866 355192
rect 43626 354864 43682 354920
rect 651470 774172 651526 774208
rect 651470 774152 651472 774172
rect 651472 774152 651524 774172
rect 651524 774152 651526 774172
rect 651470 773336 651526 773392
rect 62762 747632 62818 747688
rect 62118 746136 62174 746192
rect 62118 744096 62174 744152
rect 62118 743724 62120 743744
rect 62120 743724 62172 743744
rect 62172 743724 62174 743744
rect 62118 743688 62174 743724
rect 62118 742364 62120 742384
rect 62120 742364 62172 742384
rect 62172 742364 62174 742384
rect 62118 742328 62174 742364
rect 62394 741784 62450 741840
rect 651470 734168 651526 734224
rect 651470 732944 651526 733000
rect 651470 731720 651526 731776
rect 46202 730224 46258 730280
rect 47214 721112 47270 721168
rect 47030 719888 47086 719944
rect 45742 665896 45798 665952
rect 45558 612040 45614 612096
rect 47030 611768 47086 611824
rect 651470 731040 651526 731096
rect 651470 729816 651526 729872
rect 62118 704384 62174 704440
rect 62118 703296 62174 703352
rect 62210 701256 62266 701312
rect 651470 728492 651472 728512
rect 651472 728492 651524 728512
rect 651524 728492 651526 728512
rect 651470 728456 651526 728492
rect 62762 700848 62818 700904
rect 61382 699624 61438 699680
rect 62118 698164 62120 698184
rect 62120 698164 62172 698184
rect 62172 698164 62174 698184
rect 62118 698128 62174 698164
rect 651654 689424 651710 689480
rect 651470 688744 651526 688800
rect 652022 687248 652078 687304
rect 651470 686840 651526 686896
rect 62118 660900 62120 660920
rect 62120 660900 62172 660920
rect 62172 660900 62174 660920
rect 62118 660864 62174 660900
rect 62118 659540 62120 659560
rect 62120 659540 62172 659560
rect 62172 659540 62174 659560
rect 62118 659504 62174 659540
rect 62118 658280 62174 658336
rect 651470 685208 651526 685264
rect 62762 657600 62818 657656
rect 61382 656512 61438 656568
rect 62118 655288 62174 655344
rect 652574 684392 652630 684448
rect 651470 643184 651526 643240
rect 62118 616528 62174 616584
rect 62118 614624 62174 614680
rect 61382 613808 61438 613864
rect 62118 612620 62120 612640
rect 62120 612620 62172 612640
rect 62172 612620 62174 612640
rect 62118 612584 62174 612620
rect 652022 641824 652078 641880
rect 651470 640736 651526 640792
rect 651378 640092 651380 640112
rect 651380 640092 651432 640112
rect 651432 640092 651434 640112
rect 651378 640056 651434 640092
rect 651470 638560 651526 638616
rect 651654 638152 651710 638208
rect 62946 618024 63002 618080
rect 62762 612040 62818 612096
rect 47214 611496 47270 611552
rect 45282 598032 45338 598088
rect 651470 597896 651526 597952
rect 651470 596672 651526 596728
rect 62946 595720 63002 595776
rect 62762 594088 62818 594144
rect 45558 578448 45614 578504
rect 62118 574776 62174 574832
rect 62118 573552 62174 573608
rect 651470 595448 651526 595504
rect 651654 595176 651710 595232
rect 651470 594088 651526 594144
rect 63130 592864 63186 592920
rect 62946 571104 63002 571160
rect 651470 592728 651526 592784
rect 63130 569880 63186 569936
rect 62762 568520 62818 568576
rect 61382 557504 61438 557560
rect 45098 555600 45154 555656
rect 45650 555192 45706 555248
rect 45190 551520 45246 551576
rect 45006 549072 45062 549128
rect 44730 548664 44786 548720
rect 45006 538056 45062 538112
rect 44730 536832 44786 536888
rect 44730 535608 44786 535664
rect 45374 550704 45430 550760
rect 45374 532752 45430 532808
rect 45190 528808 45246 528864
rect 45098 527176 45154 527232
rect 44546 429664 44602 429720
rect 44638 429256 44694 429312
rect 44270 428848 44326 428904
rect 44270 428440 44326 428496
rect 44454 422320 44510 422376
rect 44454 407496 44510 407552
rect 45834 554376 45890 554432
rect 45650 428032 45706 428088
rect 45558 427624 45614 427680
rect 45006 423136 45062 423192
rect 44822 405592 44878 405648
rect 45374 421504 45430 421560
rect 45190 421096 45246 421152
rect 45190 408040 45246 408096
rect 45374 406680 45430 406736
rect 45006 402872 45062 402928
rect 44638 386416 44694 386472
rect 44270 385600 44326 385656
rect 45098 385192 45154 385248
rect 44362 379072 44418 379128
rect 44178 376216 44234 376272
rect 44546 378664 44602 378720
rect 44362 364112 44418 364168
rect 44730 377848 44786 377904
rect 44914 377440 44970 377496
rect 44730 364792 44786 364848
rect 60002 539552 60058 539608
rect 63406 556688 63462 556744
rect 62946 552608 63002 552664
rect 62118 531276 62174 531312
rect 62118 531256 62120 531276
rect 62120 531256 62172 531276
rect 62172 531256 62174 531276
rect 62118 530576 62174 530632
rect 62118 528572 62120 528592
rect 62120 528572 62172 528592
rect 62172 528572 62174 528592
rect 62118 528536 62174 528572
rect 61382 527040 61438 527096
rect 651470 553424 651526 553480
rect 651470 552336 651526 552392
rect 652022 550976 652078 551032
rect 651378 550332 651380 550352
rect 651380 550332 651432 550352
rect 651432 550332 651434 550352
rect 651378 550296 651434 550332
rect 651470 549092 651526 549128
rect 651470 549072 651472 549092
rect 651472 549072 651524 549092
rect 651524 549072 651526 549092
rect 651470 548392 651526 548448
rect 63406 527992 63462 528048
rect 62946 525680 63002 525736
rect 668398 685480 668454 685536
rect 667570 595448 667626 595504
rect 669042 733760 669098 733816
rect 669410 698264 669466 698320
rect 669226 697312 669282 697368
rect 669042 647808 669098 647864
rect 668858 638696 668914 638752
rect 668398 616800 668454 616856
rect 668398 555192 668454 555248
rect 671618 779320 671674 779376
rect 669226 607960 669282 608016
rect 669042 562264 669098 562320
rect 670422 600344 670478 600400
rect 670790 688472 670846 688528
rect 671802 714856 671858 714912
rect 671158 643592 671214 643648
rect 670974 593544 671030 593600
rect 672170 712136 672226 712192
rect 672170 690512 672226 690568
rect 671986 652840 672042 652896
rect 671802 641688 671858 641744
rect 671342 594768 671398 594824
rect 675850 895464 675906 895520
rect 676034 894648 676090 894704
rect 672538 715264 672594 715320
rect 672538 694592 672594 694648
rect 675850 893832 675906 893888
rect 676034 893036 676090 893072
rect 676034 893016 676036 893036
rect 676036 893016 676088 893036
rect 676088 893016 676090 893036
rect 676034 892608 676090 892664
rect 676034 891384 676090 891440
rect 675206 890976 675262 891032
rect 674746 888528 674802 888584
rect 676034 890160 676090 890216
rect 676034 889344 676090 889400
rect 676034 888956 676090 888992
rect 676034 888936 676036 888956
rect 676036 888936 676088 888956
rect 676088 888936 676090 888956
rect 676034 887324 676090 887360
rect 676034 887304 676036 887324
rect 676036 887304 676088 887324
rect 676088 887304 676090 887324
rect 676034 886916 676090 886952
rect 676034 886896 676036 886916
rect 676036 886896 676088 886916
rect 676088 886896 676090 886916
rect 676034 885692 676090 885728
rect 676034 885672 676036 885692
rect 676036 885672 676088 885692
rect 676088 885672 676090 885692
rect 675758 878464 675814 878520
rect 679622 891792 679678 891848
rect 678242 889752 678298 889808
rect 681002 890568 681058 890624
rect 683118 888120 683174 888176
rect 681002 880640 681058 880696
rect 683118 880368 683174 880424
rect 675574 874112 675630 874168
rect 675022 873024 675078 873080
rect 675758 872752 675814 872808
rect 675022 869388 675024 869408
rect 675024 869388 675076 869408
rect 675076 869388 675078 869408
rect 675022 869352 675078 869388
rect 674286 868536 674342 868592
rect 675022 868944 675078 869000
rect 675390 868536 675446 868592
rect 675298 865680 675354 865736
rect 675758 865408 675814 865464
rect 675666 865000 675722 865056
rect 675758 786664 675814 786720
rect 673734 778776 673790 778832
rect 674470 777416 674526 777472
rect 674102 775648 674158 775704
rect 673274 715708 673276 715728
rect 673276 715708 673328 715728
rect 673328 715708 673330 715728
rect 673274 715672 673330 715708
rect 673090 714448 673146 714504
rect 673274 714040 673330 714096
rect 672906 709144 672962 709200
rect 673458 712952 673514 713008
rect 675482 783808 675538 783864
rect 675114 782448 675170 782504
rect 675482 779320 675538 779376
rect 675482 778776 675538 778832
rect 675482 777416 675538 777472
rect 675482 775648 675538 775704
rect 673826 735664 673882 735720
rect 674102 734984 674158 735040
rect 674286 728048 674342 728104
rect 673550 712680 673606 712736
rect 672998 695544 673054 695600
rect 672722 663856 672778 663912
rect 672722 651344 672778 651400
rect 672538 618976 672594 619032
rect 672538 606464 672594 606520
rect 672262 603472 672318 603528
rect 671986 553424 672042 553480
rect 673182 685752 673238 685808
rect 673550 701020 673552 701040
rect 673552 701020 673604 701040
rect 673604 701020 673606 701040
rect 673550 700984 673606 701020
rect 673550 697076 673552 697096
rect 673552 697076 673604 697096
rect 673604 697076 673606 697096
rect 673550 697040 673606 697076
rect 673550 690004 673552 690024
rect 673552 690004 673604 690024
rect 673604 690004 673606 690024
rect 673550 689968 673606 690004
rect 673550 687656 673606 687712
rect 673918 727232 673974 727288
rect 675758 739744 675814 739800
rect 675298 738112 675354 738168
rect 675482 735664 675538 735720
rect 675482 734984 675538 735040
rect 674654 727776 674710 727832
rect 674470 727232 674526 727288
rect 674838 722200 674894 722256
rect 674654 721928 674710 721984
rect 675574 733760 675630 733816
rect 675850 728048 675906 728104
rect 676034 727776 676090 727832
rect 681002 726824 681058 726880
rect 673642 682488 673698 682544
rect 674010 716488 674066 716544
rect 674010 716080 674066 716136
rect 674010 713668 674012 713688
rect 674012 713668 674064 713688
rect 674064 713668 674066 713688
rect 674010 713632 674066 713668
rect 674010 713244 674066 713280
rect 674010 713224 674012 713244
rect 674012 713224 674064 713244
rect 674064 713224 674066 713244
rect 674010 712428 674066 712464
rect 674010 712408 674012 712428
rect 674012 712408 674064 712428
rect 674064 712408 674066 712428
rect 674010 711184 674066 711240
rect 674010 710404 674012 710424
rect 674012 710404 674064 710424
rect 674064 710404 674066 710424
rect 674010 710368 674066 710404
rect 674010 709996 674012 710016
rect 674012 709996 674064 710016
rect 674064 709996 674066 710016
rect 674010 709960 674066 709996
rect 674010 709588 674012 709608
rect 674012 709588 674064 709608
rect 674064 709588 674066 709608
rect 674010 709552 674066 709588
rect 674010 707956 674012 707976
rect 674012 707956 674064 707976
rect 674064 707956 674066 707976
rect 674010 707920 674066 707956
rect 674010 705356 674066 705392
rect 674010 705336 674012 705356
rect 674012 705336 674064 705356
rect 674064 705336 674066 705356
rect 674010 705064 674066 705120
rect 674746 712952 674802 713008
rect 674378 712680 674434 712736
rect 674930 712816 674986 712872
rect 674930 712136 674986 712192
rect 683118 726416 683174 726472
rect 681002 712000 681058 712056
rect 675390 710776 675446 710832
rect 683302 711592 683358 711648
rect 683118 708736 683174 708792
rect 683486 708328 683542 708384
rect 674746 707104 674802 707160
rect 674378 706696 674434 706752
rect 683118 705472 683174 705528
rect 675850 705336 675906 705392
rect 673642 682216 673698 682272
rect 675114 700984 675170 701040
rect 675114 698264 675170 698320
rect 675114 697312 675170 697368
rect 675114 697040 675170 697096
rect 674930 695544 674986 695600
rect 675390 696768 675446 696824
rect 675114 694592 675170 694648
rect 674102 689152 674158 689208
rect 673642 671336 673698 671392
rect 673642 670520 673698 670576
rect 673366 669432 673422 669488
rect 673642 668888 673698 668944
rect 673642 667256 673698 667312
rect 673642 666032 673698 666088
rect 673642 664808 673698 664864
rect 673366 664128 673422 664184
rect 673642 663856 673698 663912
rect 674010 670928 674066 670984
rect 674010 670132 674066 670168
rect 674010 670112 674012 670132
rect 674012 670112 674064 670132
rect 674064 670112 674066 670132
rect 674010 669704 674066 669760
rect 674010 668516 674012 668536
rect 674012 668516 674064 668536
rect 674064 668516 674066 668536
rect 674010 668480 674066 668516
rect 674010 668072 674066 668128
rect 674010 667664 674066 667720
rect 674010 665644 674066 665680
rect 674010 665624 674012 665644
rect 674012 665624 674064 665644
rect 674064 665624 674066 665644
rect 674010 663584 674066 663640
rect 674010 662768 674066 662824
rect 673826 661952 673882 662008
rect 674010 661580 674012 661600
rect 674012 661580 674064 661600
rect 674064 661580 674066 661600
rect 674010 661544 674066 661580
rect 674010 661156 674066 661192
rect 674010 661136 674012 661156
rect 674012 661136 674064 661156
rect 674064 661136 674066 661156
rect 674010 660084 674012 660104
rect 674012 660084 674064 660104
rect 674064 660084 674066 660104
rect 674010 660048 674066 660084
rect 673274 659640 673330 659696
rect 673090 620200 673146 620256
rect 673090 619828 673092 619848
rect 673092 619828 673144 619848
rect 673144 619828 673146 619848
rect 673090 619792 673146 619828
rect 672906 618568 672962 618624
rect 673090 604288 673146 604344
rect 672906 599664 672962 599720
rect 672722 576408 672778 576464
rect 674010 655580 674066 655616
rect 674010 655560 674012 655580
rect 674012 655560 674064 655580
rect 674064 655560 674066 655580
rect 674010 654100 674012 654120
rect 674012 654100 674064 654120
rect 674064 654100 674066 654120
rect 674010 654064 674066 654100
rect 673642 649168 673698 649224
rect 673458 625912 673514 625968
rect 673458 620608 673514 620664
rect 673458 619384 673514 619440
rect 673458 616564 673460 616584
rect 673460 616564 673512 616584
rect 673512 616564 673514 616584
rect 673458 616528 673514 616564
rect 673458 614916 673514 614952
rect 673458 614896 673460 614916
rect 673460 614896 673512 614916
rect 673512 614896 673514 614916
rect 673458 611380 673514 611416
rect 673458 611360 673460 611380
rect 673460 611360 673512 611380
rect 673512 611360 673514 611380
rect 673458 600072 673514 600128
rect 673458 599004 673514 599040
rect 673458 598984 673460 599004
rect 673460 598984 673512 599004
rect 673512 598984 673514 599004
rect 674010 647284 674066 647320
rect 674010 647264 674012 647284
rect 674012 647264 674064 647284
rect 674064 647264 674066 647284
rect 673826 644680 673882 644736
rect 674010 643084 674012 643104
rect 674012 643084 674064 643104
rect 674064 643084 674066 643104
rect 674010 643048 674066 643084
rect 675114 690512 675170 690568
rect 674930 689968 674986 690024
rect 675114 689152 675170 689208
rect 675114 688472 675170 688528
rect 675298 687656 675354 687712
rect 674930 687112 674986 687168
rect 675758 686160 675814 686216
rect 675114 685752 675170 685808
rect 675482 685480 675538 685536
rect 675850 682524 675852 682544
rect 675852 682524 675904 682544
rect 675904 682524 675906 682544
rect 675850 682488 675906 682524
rect 675666 682216 675722 682272
rect 682382 682080 682438 682136
rect 678242 681808 678298 681864
rect 675298 676368 675354 676424
rect 678242 666984 678298 667040
rect 682382 666576 682438 666632
rect 683210 665352 683266 665408
rect 683394 663312 683450 663368
rect 675850 660048 675906 660104
rect 683118 660048 683174 660104
rect 675114 655560 675170 655616
rect 674930 654064 674986 654120
rect 675390 652840 675446 652896
rect 675114 651344 675170 651400
rect 674562 644000 674618 644056
rect 674102 636792 674158 636848
rect 674010 626320 674066 626376
rect 674010 625540 674012 625560
rect 674012 625540 674064 625560
rect 674064 625540 674066 625560
rect 674010 625504 674066 625540
rect 674010 625116 674066 625152
rect 674010 625096 674012 625116
rect 674012 625096 674064 625116
rect 674064 625096 674066 625116
rect 674010 624708 674066 624744
rect 674010 624688 674012 624708
rect 674012 624688 674064 624708
rect 674064 624688 674066 624708
rect 674010 624316 674012 624336
rect 674012 624316 674064 624336
rect 674064 624316 674066 624336
rect 674010 624280 674066 624316
rect 674010 623892 674066 623928
rect 674010 623872 674012 623892
rect 674012 623872 674064 623892
rect 674064 623872 674066 623892
rect 674010 623500 674012 623520
rect 674012 623500 674064 623520
rect 674064 623500 674066 623520
rect 674010 623464 674066 623500
rect 674010 623076 674066 623112
rect 674010 623056 674012 623076
rect 674012 623056 674064 623076
rect 674064 623056 674066 623076
rect 674010 622684 674012 622704
rect 674012 622684 674064 622704
rect 674064 622684 674066 622704
rect 674010 622648 674066 622684
rect 674010 622260 674066 622296
rect 674010 622240 674012 622260
rect 674012 622240 674064 622260
rect 674064 622240 674066 622260
rect 674010 621188 674012 621208
rect 674012 621188 674064 621208
rect 674064 621188 674066 621208
rect 674010 621152 674066 621188
rect 674470 640192 674526 640248
rect 675390 649712 675446 649768
rect 675390 649168 675446 649224
rect 675758 648624 675814 648680
rect 675390 647808 675446 647864
rect 675114 647264 675170 647320
rect 675298 644680 675354 644736
rect 675390 643592 675446 643648
rect 675114 643048 675170 643104
rect 675298 641688 675354 641744
rect 674746 626592 674802 626648
rect 675482 638696 675538 638752
rect 675850 636828 675852 636848
rect 675852 636828 675904 636848
rect 675904 636828 675906 636848
rect 675850 636792 675906 636828
rect 675482 636520 675538 636576
rect 683210 636520 683266 636576
rect 681002 636112 681058 636168
rect 674470 618160 674526 618216
rect 673918 602928 673974 602984
rect 673642 591776 673698 591832
rect 673458 591232 673514 591288
rect 673642 580624 673698 580680
rect 673458 579400 673514 579456
rect 673642 578176 673698 578232
rect 673458 576680 673514 576736
rect 673642 574504 673698 574560
rect 673642 572464 673698 572520
rect 673642 558048 673698 558104
rect 673274 557504 673330 557560
rect 673458 549208 673514 549264
rect 672906 527584 672962 527640
rect 672906 491272 672962 491328
rect 671986 474816 672042 474872
rect 669410 455368 669466 455424
rect 672446 453736 672502 453792
rect 60002 430616 60058 430672
rect 45834 427352 45890 427408
rect 45834 426808 45890 426864
rect 45558 384784 45614 384840
rect 46018 423952 46074 424008
rect 53838 407768 53894 407824
rect 46018 400152 46074 400208
rect 61382 429256 61438 429312
rect 63130 427080 63186 427136
rect 62118 404096 62174 404152
rect 62118 402600 62174 402656
rect 62118 400560 62174 400616
rect 657542 403280 657598 403336
rect 652022 400832 652078 400888
rect 63130 400152 63186 400208
rect 62118 399336 62174 399392
rect 61382 398248 61438 398304
rect 51078 395664 51134 395720
rect 61382 386416 61438 386472
rect 46018 384376 46074 384432
rect 45834 383968 45890 384024
rect 45650 383560 45706 383616
rect 45282 381384 45338 381440
rect 44546 361528 44602 361584
rect 44822 355136 44878 355192
rect 44638 354864 44694 354920
rect 43258 353640 43314 353696
rect 42338 352960 42394 353016
rect 35806 344256 35862 344312
rect 35622 343848 35678 343904
rect 35806 343440 35862 343496
rect 40406 343848 40462 343904
rect 35806 341808 35862 341864
rect 39670 341808 39726 341864
rect 39854 341808 39910 341864
rect 35806 341028 35808 341048
rect 35808 341028 35860 341048
rect 35860 341028 35862 341048
rect 35806 340992 35862 341028
rect 40222 342236 40278 342272
rect 40222 342216 40224 342236
rect 40224 342216 40276 342236
rect 40276 342216 40278 342236
rect 45374 362888 45430 362944
rect 45190 343304 45246 343360
rect 45006 342488 45062 342544
rect 45466 342236 45522 342272
rect 45466 342216 45468 342236
rect 45468 342216 45520 342236
rect 45520 342216 45522 342236
rect 42246 341264 42302 341320
rect 40130 341028 40132 341048
rect 40132 341028 40184 341048
rect 40184 341028 40186 341048
rect 40130 340992 40186 341028
rect 45834 353932 45890 353968
rect 45834 353912 45836 353932
rect 45836 353912 45888 353932
rect 45888 353912 45890 353932
rect 45834 353676 45836 353696
rect 45836 353676 45888 353696
rect 45888 353676 45890 353696
rect 45834 353640 45890 353676
rect 47122 383152 47178 383208
rect 46938 382336 46994 382392
rect 46570 363160 46626 363216
rect 47122 354320 47178 354376
rect 63406 385872 63462 385928
rect 62946 381792 63002 381848
rect 62118 360848 62174 360904
rect 62118 359760 62174 359816
rect 62118 357720 62174 357776
rect 61382 355952 61438 356008
rect 651470 373224 651526 373280
rect 652206 395256 652262 395312
rect 654782 382880 654838 382936
rect 652206 373904 652262 373960
rect 652022 372136 652078 372192
rect 673458 535200 673514 535256
rect 673274 529080 673330 529136
rect 673090 483112 673146 483168
rect 674838 600072 674894 600128
rect 674562 599392 674618 599448
rect 674378 598304 674434 598360
rect 674194 597352 674250 597408
rect 674010 581576 674066 581632
rect 674010 581052 674066 581088
rect 674010 581032 674012 581052
rect 674012 581032 674064 581052
rect 674064 581032 674066 581052
rect 674010 580252 674012 580272
rect 674012 580252 674064 580272
rect 674064 580252 674066 580272
rect 674010 580216 674066 580252
rect 674010 579808 674066 579864
rect 674010 578992 674066 579048
rect 674010 578584 674066 578640
rect 674010 577396 674012 577416
rect 674012 577396 674064 577416
rect 674064 577396 674066 577416
rect 674010 577360 674066 577396
rect 674010 576972 674066 577008
rect 674010 576952 674012 576972
rect 674012 576952 674064 576972
rect 674064 576952 674066 576972
rect 674010 575728 674066 575784
rect 674010 574096 674066 574152
rect 674010 572892 674066 572928
rect 674010 572872 674012 572892
rect 674012 572872 674064 572892
rect 674064 572872 674066 572892
rect 674010 572056 674066 572112
rect 674010 565836 674012 565856
rect 674012 565836 674064 565856
rect 674064 565836 674066 565856
rect 674010 565800 674066 565836
rect 673918 555464 673974 555520
rect 674010 554648 674066 554704
rect 674102 552880 674158 552936
rect 674838 598576 674894 598632
rect 675850 626592 675906 626648
rect 681002 621968 681058 622024
rect 683394 617888 683450 617944
rect 683118 617480 683174 617536
rect 683302 617072 683358 617128
rect 675850 616800 675906 616856
rect 683118 615476 683120 615496
rect 683120 615476 683172 615496
rect 683172 615476 683174 615496
rect 683118 615440 683174 615476
rect 675390 611360 675446 611416
rect 675390 608232 675446 608288
rect 675390 607960 675446 608016
rect 675390 606464 675446 606520
rect 675482 604560 675538 604616
rect 675390 604288 675446 604344
rect 675482 603472 675538 603528
rect 675390 602928 675446 602984
rect 675482 600344 675538 600400
rect 675758 599800 675814 599856
rect 675482 599664 675538 599720
rect 675482 599120 675538 599176
rect 675298 598984 675354 599040
rect 675482 598576 675538 598632
rect 675758 598576 675814 598632
rect 675482 597352 675538 597408
rect 675298 596264 675354 596320
rect 674746 592864 674802 592920
rect 675390 595448 675446 595504
rect 675482 594768 675538 594824
rect 675390 593544 675446 593600
rect 675850 592884 675906 592920
rect 675850 592864 675852 592884
rect 675852 592864 675904 592884
rect 675904 592864 675906 592884
rect 675482 592048 675538 592104
rect 674930 589192 674986 589248
rect 675850 591776 675906 591832
rect 675850 591268 675852 591288
rect 675852 591268 675904 591288
rect 675904 591268 675906 591288
rect 675850 591232 675906 591268
rect 675850 589228 675852 589248
rect 675852 589228 675904 589248
rect 675904 589228 675906 589248
rect 675850 589192 675906 589228
rect 675114 586200 675170 586256
rect 675482 586200 675538 586256
rect 673826 536016 673882 536072
rect 674010 535644 674012 535664
rect 674012 535644 674064 535664
rect 674064 535644 674066 535664
rect 674010 535608 674066 535644
rect 674010 534792 674066 534848
rect 673826 534384 673882 534440
rect 674010 534112 674066 534168
rect 674010 533588 674066 533624
rect 674010 533568 674012 533588
rect 674012 533568 674064 533588
rect 674064 533568 674066 533588
rect 674010 533332 674012 533352
rect 674012 533332 674064 533352
rect 674064 533332 674066 533352
rect 674010 533296 674066 533332
rect 674010 532772 674066 532808
rect 674010 532752 674012 532772
rect 674012 532752 674064 532772
rect 674064 532752 674066 532772
rect 674010 532516 674012 532536
rect 674012 532516 674064 532536
rect 674064 532516 674066 532536
rect 674010 532480 674066 532516
rect 674010 531956 674066 531992
rect 674010 531936 674012 531956
rect 674012 531936 674064 531956
rect 674064 531936 674066 531956
rect 674010 531700 674012 531720
rect 674012 531700 674064 531720
rect 674064 531700 674066 531720
rect 674010 531664 674066 531700
rect 674010 531120 674066 531176
rect 673826 530068 673828 530088
rect 673828 530068 673880 530088
rect 673880 530068 673882 530088
rect 673826 530032 673882 530068
rect 674010 529660 674012 529680
rect 674012 529660 674064 529680
rect 674064 529660 674066 529680
rect 674010 529624 674066 529660
rect 674654 581576 674710 581632
rect 675850 577768 675906 577824
rect 675850 576680 675906 576736
rect 684038 592592 684094 592648
rect 678242 576408 678298 576464
rect 674654 571376 674710 571432
rect 684038 575592 684094 575648
rect 684222 573960 684278 574016
rect 683394 571920 683450 571976
rect 683118 570696 683174 570752
rect 676218 569472 676274 569528
rect 675390 565800 675446 565856
rect 676218 565528 676274 565584
rect 675758 562672 675814 562728
rect 675114 562264 675170 562320
rect 675390 561856 675446 561912
rect 674470 537104 674526 537160
rect 674010 529080 674066 529136
rect 674010 528436 674012 528456
rect 674012 528436 674064 528456
rect 674064 528436 674066 528456
rect 674010 528400 674066 528436
rect 674010 524628 674012 524648
rect 674012 524628 674064 524648
rect 674064 524628 674066 524648
rect 674010 524592 674066 524628
rect 674378 492360 674434 492416
rect 673826 492088 673882 492144
rect 674010 491680 674066 491736
rect 674010 490900 674012 490920
rect 674012 490900 674064 490920
rect 674064 490900 674066 490920
rect 674010 490864 674066 490900
rect 674010 490084 674012 490104
rect 674012 490084 674064 490104
rect 674064 490084 674066 490104
rect 674010 490048 674066 490084
rect 674010 489660 674066 489696
rect 674010 489640 674012 489660
rect 674012 489640 674064 489660
rect 674064 489640 674066 489660
rect 674010 489268 674012 489288
rect 674012 489268 674064 489288
rect 674064 489268 674066 489288
rect 674010 489232 674066 489268
rect 674010 488452 674012 488472
rect 674012 488452 674064 488472
rect 674064 488452 674066 488472
rect 674010 488416 674066 488452
rect 674010 485968 674066 486024
rect 673826 485560 673882 485616
rect 674010 485152 674066 485208
rect 673642 484336 673698 484392
rect 675390 558048 675446 558104
rect 675390 557504 675446 557560
rect 675114 555464 675170 555520
rect 675390 555192 675446 555248
rect 675114 554648 675170 554704
rect 674838 549752 674894 549808
rect 674654 482704 674710 482760
rect 674010 482332 674012 482352
rect 674012 482332 674064 482352
rect 674064 482332 674066 482352
rect 674010 482296 674066 482332
rect 675758 553832 675814 553888
rect 675390 553424 675446 553480
rect 675206 552880 675262 552936
rect 675758 552064 675814 552120
rect 675390 549752 675446 549808
rect 675390 549208 675446 549264
rect 675482 547596 675538 547632
rect 675482 547576 675484 547596
rect 675484 547576 675536 547596
rect 675536 547576 675538 547596
rect 676034 547576 676090 547632
rect 677414 547576 677470 547632
rect 675298 544448 675354 544504
rect 675850 537104 675906 537160
rect 675850 524612 675906 524648
rect 675850 524592 675852 524612
rect 675852 524592 675904 524612
rect 675904 524592 675906 524612
rect 675574 513712 675630 513768
rect 675206 508816 675262 508872
rect 675022 501880 675078 501936
rect 675298 487600 675354 487656
rect 675114 481888 675170 481944
rect 674838 479984 674894 480040
rect 673458 464752 673514 464808
rect 673274 455388 673330 455424
rect 673274 455368 673276 455388
rect 673276 455368 673328 455388
rect 673328 455368 673330 455388
rect 673826 455812 673828 455832
rect 673828 455812 673880 455832
rect 673880 455812 673882 455832
rect 673826 455776 673882 455812
rect 673274 454996 673276 455016
rect 673276 454996 673328 455016
rect 673328 454996 673330 455016
rect 673274 454960 673330 454996
rect 673044 454588 673046 454608
rect 673046 454588 673098 454608
rect 673098 454588 673100 454608
rect 673044 454552 673100 454588
rect 672952 454316 672954 454336
rect 672954 454316 673006 454336
rect 673006 454316 673008 454336
rect 672952 454280 673008 454316
rect 674286 454316 674288 454336
rect 674288 454316 674340 454336
rect 674340 454316 674342 454336
rect 674286 454280 674342 454316
rect 672814 454044 672816 454064
rect 672816 454044 672868 454064
rect 672868 454044 672870 454064
rect 672814 454008 672870 454044
rect 675298 480664 675354 480720
rect 676034 513712 676090 513768
rect 676126 508816 676182 508872
rect 678242 547304 678298 547360
rect 681002 547032 681058 547088
rect 681002 530984 681058 531040
rect 678242 530576 678298 530632
rect 683210 527312 683266 527368
rect 684222 528128 684278 528184
rect 683578 526904 683634 526960
rect 683394 526496 683450 526552
rect 677874 525680 677930 525736
rect 677690 524456 677746 524512
rect 683118 524864 683174 524920
rect 675850 501880 675906 501936
rect 676034 492360 676090 492416
rect 675850 490456 675906 490512
rect 676034 488008 676090 488064
rect 675666 454552 675722 454608
rect 675298 454008 675354 454064
rect 675114 453736 675170 453792
rect 678242 487192 678298 487248
rect 676586 484506 676642 484562
rect 676126 479984 676182 480040
rect 676218 477400 676274 477456
rect 676126 455776 676182 455832
rect 675942 447752 675998 447808
rect 683394 486784 683450 486840
rect 681002 486376 681058 486432
rect 683118 481072 683174 481128
rect 677506 440272 677562 440328
rect 676034 410488 676090 410544
rect 674562 403416 674618 403472
rect 672630 401920 672686 401976
rect 672814 401648 672870 401704
rect 671986 397160 672042 397216
rect 669226 393488 669282 393544
rect 668858 386008 668914 386064
rect 668858 382880 668914 382936
rect 651470 370640 651526 370696
rect 654782 358536 654838 358592
rect 63406 357312 63462 357368
rect 652022 356632 652078 356688
rect 62946 354456 63002 354512
rect 51722 353232 51778 353288
rect 46938 352960 46994 353016
rect 46018 343848 46074 343904
rect 62946 341672 63002 341728
rect 62762 341400 62818 341456
rect 45650 340720 45706 340776
rect 39670 340176 39726 340232
rect 35530 339768 35586 339824
rect 35806 339768 35862 339824
rect 37094 336504 37150 336560
rect 46938 339224 46994 339280
rect 45558 338816 45614 338872
rect 45374 337864 45430 337920
rect 35806 335688 35862 335744
rect 38842 335688 38898 335744
rect 35806 334464 35862 334520
rect 44178 334600 44234 334656
rect 44362 334600 44418 334656
rect 40314 332832 40370 332888
rect 42890 332832 42946 332888
rect 39854 332424 39910 332480
rect 42430 326984 42486 327040
rect 41786 325352 41842 325408
rect 41786 324808 41842 324864
rect 42062 322768 42118 322824
rect 42062 321136 42118 321192
rect 42154 320456 42210 320512
rect 41878 319912 41934 319968
rect 42062 319912 42118 319968
rect 43074 332424 43130 332480
rect 42890 321136 42946 321192
rect 42614 320728 42670 320784
rect 43074 320456 43130 320512
rect 45282 326984 45338 327040
rect 44362 322768 44418 322824
rect 44178 319912 44234 319968
rect 42430 319640 42486 319696
rect 42246 318960 42302 319016
rect 41786 317328 41842 317384
rect 42154 315968 42210 316024
rect 42154 315424 42210 315480
rect 45558 315424 45614 315480
rect 42062 313656 42118 313712
rect 42430 312704 42486 312760
rect 51722 334056 51778 334112
rect 50342 333104 50398 333160
rect 42430 310392 42486 310448
rect 46938 310392 46994 310448
rect 42062 309032 42118 309088
rect 35622 300872 35678 300928
rect 46202 300464 46258 300520
rect 44178 299648 44234 299704
rect 35806 298832 35862 298888
rect 41786 298696 41842 298752
rect 41786 296520 41842 296576
rect 42798 296520 42854 296576
rect 35438 296384 35494 296440
rect 35622 295976 35678 296032
rect 35806 295604 35808 295624
rect 35808 295604 35860 295624
rect 35860 295604 35862 295624
rect 35806 295568 35862 295604
rect 35806 295160 35862 295216
rect 33782 294752 33838 294808
rect 32402 294344 32458 294400
rect 35806 293120 35862 293176
rect 35806 292712 35862 292768
rect 35806 291080 35862 291136
rect 35622 290264 35678 290320
rect 32402 284824 32458 284880
rect 41786 295296 41842 295352
rect 41786 292168 41842 292224
rect 41786 291896 41842 291952
rect 41786 290264 41842 290320
rect 41786 289176 41842 289232
rect 40682 284280 40738 284336
rect 41786 278432 41842 278488
rect 42062 277752 42118 277808
rect 41786 277072 41842 277128
rect 42062 276664 42118 276720
rect 42430 278704 42486 278760
rect 42614 276664 42670 276720
rect 42246 275848 42302 275904
rect 41786 274216 41842 274272
rect 42338 273128 42394 273184
rect 42430 272856 42486 272912
rect 41970 272312 42026 272368
rect 41786 270408 41842 270464
rect 41878 270000 41934 270056
rect 40682 267008 40738 267064
rect 35806 257080 35862 257136
rect 42154 266192 42210 266248
rect 43166 295296 43222 295352
rect 43626 292168 43682 292224
rect 43350 290264 43406 290320
rect 35806 255856 35862 255912
rect 39762 255856 39818 255912
rect 42798 255856 42854 255912
rect 35806 253816 35862 253872
rect 39578 253816 39634 253872
rect 42798 253816 42854 253872
rect 35622 253408 35678 253464
rect 35806 253000 35862 253056
rect 40958 253000 41014 253056
rect 35806 252184 35862 252240
rect 40498 252184 40554 252240
rect 35806 250552 35862 250608
rect 35806 249328 35862 249384
rect 39394 249328 39450 249384
rect 42430 252184 42486 252240
rect 35622 247696 35678 247752
rect 35806 246880 35862 246936
rect 41510 246880 41566 246936
rect 39210 244976 39266 245032
rect 42062 240080 42118 240136
rect 43258 253000 43314 253056
rect 43166 249328 43222 249384
rect 42982 244976 43038 245032
rect 42430 237360 42486 237416
rect 41786 236544 41842 236600
rect 42430 235864 42486 235920
rect 42430 233416 42486 233472
rect 42430 233144 42486 233200
rect 42246 233008 42302 233064
rect 42062 230968 42118 231024
rect 41970 228928 42026 228984
rect 42246 226072 42302 226128
rect 42614 225528 42670 225584
rect 42430 224848 42486 224904
rect 42154 223216 42210 223272
rect 35806 217912 35862 217968
rect 35806 214648 35862 214704
rect 35806 214240 35862 214296
rect 35438 212200 35494 212256
rect 43626 277752 43682 277808
rect 45006 298016 45062 298072
rect 44362 297200 44418 297256
rect 44178 256808 44234 256864
rect 44730 293936 44786 293992
rect 44546 293528 44602 293584
rect 44546 273128 44602 273184
rect 44730 272856 44786 272912
rect 44822 256400 44878 256456
rect 44638 254768 44694 254824
rect 44362 254360 44418 254416
rect 44362 252728 44418 252784
rect 44178 251504 44234 251560
rect 43626 246880 43682 246936
rect 35622 211792 35678 211848
rect 39578 211792 39634 211848
rect 42798 211792 42854 211848
rect 35806 211384 35862 211440
rect 35806 210160 35862 210216
rect 35622 208936 35678 208992
rect 35806 208548 35862 208584
rect 35806 208528 35808 208548
rect 35808 208528 35860 208548
rect 35860 208528 35862 208548
rect 40038 208120 40094 208176
rect 35806 207712 35862 207768
rect 35806 206080 35862 206136
rect 40498 207712 40554 207768
rect 40222 205672 40278 205728
rect 35622 204856 35678 204912
rect 35806 204040 35862 204096
rect 40406 204040 40462 204096
rect 28538 203632 28594 203688
rect 41694 208120 41750 208176
rect 42982 207712 43038 207768
rect 41326 206488 41382 206544
rect 40958 204448 41014 204504
rect 40774 203224 40830 203280
rect 42798 203224 42854 203280
rect 28538 199280 28594 199336
rect 42246 199280 42302 199336
rect 42062 196968 42118 197024
rect 41878 195200 41934 195256
rect 42246 194928 42302 194984
rect 41786 193160 41842 193216
rect 42062 191528 42118 191584
rect 42246 190848 42302 190904
rect 42430 186768 42486 186824
rect 41786 186360 41842 186416
rect 41786 185952 41842 186008
rect 41786 184048 41842 184104
rect 43166 204448 43222 204504
rect 43350 204348 43352 204368
rect 43352 204348 43404 204368
rect 43404 204348 43406 204368
rect 43350 204312 43406 204348
rect 42430 180648 42486 180704
rect 42062 179288 42118 179344
rect 44178 240080 44234 240136
rect 44362 226072 44418 226128
rect 48962 289856 49018 289912
rect 46202 258032 46258 258088
rect 45558 255584 45614 255640
rect 45006 255176 45062 255232
rect 45006 251912 45062 251968
rect 45190 249056 45246 249112
rect 45006 233144 45062 233200
rect 45190 230968 45246 231024
rect 44822 213696 44878 213752
rect 45926 251096 45982 251152
rect 45742 248648 45798 248704
rect 45742 233416 45798 233472
rect 46110 248240 46166 248296
rect 47582 246608 47638 246664
rect 46110 235864 46166 235920
rect 45926 224848 45982 224904
rect 45558 212880 45614 212936
rect 44638 212064 44694 212120
rect 46938 209616 46994 209672
rect 44362 208392 44418 208448
rect 44178 207168 44234 207224
rect 43994 204312 44050 204368
rect 43810 204040 43866 204096
rect 43994 191528 44050 191584
rect 44638 205264 44694 205320
rect 44362 196968 44418 197024
rect 44822 204856 44878 204912
rect 44638 190848 44694 190904
rect 44178 186768 44234 186824
rect 46202 203496 46258 203552
rect 46938 180648 46994 180704
rect 47766 214920 47822 214976
rect 47766 213288 47822 213344
rect 47950 210840 48006 210896
rect 48778 206488 48834 206544
rect 48318 194384 48374 194440
rect 48778 192344 48834 192400
rect 47766 190440 47822 190496
rect 49146 247424 49202 247480
rect 49514 208120 49570 208176
rect 49514 196424 49570 196480
rect 50526 290672 50582 290728
rect 50710 179288 50766 179344
rect 53838 320728 53894 320784
rect 53102 319640 53158 319696
rect 62118 317364 62120 317384
rect 62120 317364 62172 317384
rect 62172 317364 62174 317384
rect 62118 317328 62174 317364
rect 62118 315988 62174 316024
rect 62118 315968 62120 315988
rect 62120 315968 62172 315988
rect 62172 315968 62174 315988
rect 62118 314764 62174 314800
rect 62118 314744 62120 314764
rect 62120 314744 62172 314764
rect 62172 314744 62174 314764
rect 651378 328072 651434 328128
rect 652390 352552 652446 352608
rect 653402 338680 653458 338736
rect 652390 329704 652446 329760
rect 652022 326848 652078 326904
rect 651378 325644 651434 325680
rect 658922 346432 658978 346488
rect 651378 325624 651380 325644
rect 651380 325624 651432 325644
rect 651432 325624 651434 325644
rect 63130 314064 63186 314120
rect 653402 313248 653458 313304
rect 62946 312976 63002 313032
rect 62762 311752 62818 311808
rect 652298 309848 652354 309904
rect 59910 309032 59966 309088
rect 651378 303320 651434 303376
rect 652298 302096 652354 302152
rect 53102 301280 53158 301336
rect 654782 300872 654838 300928
rect 651470 300600 651526 300656
rect 62762 298696 62818 298752
rect 651470 298696 651526 298752
rect 62118 295452 62174 295488
rect 62118 295432 62120 295452
rect 62120 295432 62172 295452
rect 62172 295432 62174 295452
rect 54482 266192 54538 266248
rect 62118 294092 62174 294128
rect 62118 294072 62120 294092
rect 62120 294072 62172 294092
rect 62172 294072 62174 294092
rect 62302 292712 62358 292768
rect 62118 292460 62174 292496
rect 62118 292440 62120 292460
rect 62120 292440 62172 292460
rect 62172 292440 62174 292460
rect 62118 290944 62174 291000
rect 651470 297472 651526 297528
rect 652666 296792 652722 296848
rect 652114 295296 652170 295352
rect 651470 294208 651526 294264
rect 651470 292984 651526 293040
rect 651470 290400 651526 290456
rect 62762 289720 62818 289776
rect 651470 289176 651526 289232
rect 62118 288516 62174 288552
rect 62118 288496 62120 288516
rect 62120 288496 62172 288516
rect 62172 288496 62174 288516
rect 651746 288496 651802 288552
rect 651470 287408 651526 287464
rect 63130 287136 63186 287192
rect 62118 285912 62174 285968
rect 62118 284436 62174 284472
rect 62118 284416 62120 284436
rect 62120 284416 62172 284436
rect 62172 284416 62174 284436
rect 58622 278704 58678 278760
rect 57242 275848 57298 275904
rect 62762 283192 62818 283248
rect 62118 280880 62174 280936
rect 61382 280336 61438 280392
rect 60002 256672 60058 256728
rect 55862 223216 55918 223272
rect 61290 217912 61346 217968
rect 62946 282104 63002 282160
rect 651470 285912 651526 285968
rect 651470 284688 651526 284744
rect 652390 291488 652446 291544
rect 652114 283464 652170 283520
rect 651930 282104 651986 282160
rect 651654 280880 651710 280936
rect 651470 280356 651526 280392
rect 651470 280336 651472 280356
rect 651472 280336 651524 280356
rect 651524 280336 651526 280356
rect 63130 267008 63186 267064
rect 462226 272312 462282 272368
rect 470414 272620 470416 272640
rect 470416 272620 470468 272640
rect 470468 272620 470470 272640
rect 470414 272584 470470 272620
rect 470598 272620 470600 272640
rect 470600 272620 470652 272640
rect 470652 272620 470654 272640
rect 470598 272584 470654 272620
rect 470414 272312 470470 272368
rect 470598 271904 470654 271960
rect 478050 271904 478106 271960
rect 489918 272720 489974 272776
rect 495714 272720 495770 272776
rect 523866 271124 523868 271144
rect 523868 271124 523920 271144
rect 523920 271124 523922 271144
rect 523866 271088 523922 271124
rect 525338 271088 525394 271144
rect 530398 270136 530454 270192
rect 534078 270136 534134 270192
rect 537298 275032 537354 275088
rect 538126 275032 538182 275088
rect 537758 269900 537760 269920
rect 537760 269900 537812 269920
rect 537812 269900 537814 269920
rect 537758 269864 537814 269900
rect 538310 269864 538366 269920
rect 539322 274488 539378 274544
rect 542266 274760 542322 274816
rect 543186 274780 543242 274816
rect 543186 274760 543188 274780
rect 543188 274760 543240 274780
rect 543240 274760 543242 274780
rect 543830 274508 543886 274544
rect 543830 274488 543832 274508
rect 543832 274488 543884 274508
rect 543884 274488 543886 274508
rect 544014 273264 544070 273320
rect 552570 273264 552626 273320
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553490 255604 553546 255640
rect 553490 255584 553492 255604
rect 553492 255584 553544 255604
rect 553544 255584 553546 255604
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 554042 249056 554098 249112
rect 553858 246880 553914 246936
rect 553674 242528 553730 242584
rect 62946 225528 63002 225584
rect 140042 229064 140098 229120
rect 139306 228248 139362 228304
rect 141146 226108 141148 226128
rect 141148 226108 141200 226128
rect 141200 226108 141202 226128
rect 141146 226072 141202 226108
rect 142434 230444 142490 230480
rect 142434 230424 142436 230444
rect 142436 230424 142488 230444
rect 142488 230424 142490 230444
rect 142986 228248 143042 228304
rect 140778 220360 140834 220416
rect 142342 220360 142398 220416
rect 142158 220108 142214 220144
rect 142158 220088 142160 220108
rect 142160 220088 142212 220108
rect 142212 220088 142214 220108
rect 141974 219680 142030 219736
rect 144090 230424 144146 230480
rect 143998 229492 144054 229528
rect 143998 229472 144000 229492
rect 144000 229472 144052 229492
rect 144052 229472 144054 229492
rect 145378 229472 145434 229528
rect 146206 229336 146262 229392
rect 145194 226108 145196 226128
rect 145196 226108 145248 226128
rect 145248 226108 145250 226128
rect 145194 226072 145250 226108
rect 145930 222264 145986 222320
rect 144826 220360 144882 220416
rect 144182 219680 144238 219736
rect 147126 229064 147182 229120
rect 147586 229744 147642 229800
rect 147954 229744 148010 229800
rect 147770 229356 147826 229392
rect 147770 229336 147772 229356
rect 147772 229336 147824 229356
rect 147824 229336 147826 229356
rect 147310 222944 147366 223000
rect 147126 222300 147128 222320
rect 147128 222300 147180 222320
rect 147180 222300 147182 222320
rect 147126 222264 147182 222300
rect 150346 229336 150402 229392
rect 151910 223080 151966 223136
rect 151450 222944 151506 223000
rect 151634 222672 151690 222728
rect 152094 222672 152150 222728
rect 151726 220516 151782 220552
rect 151726 220496 151728 220516
rect 151728 220496 151780 220516
rect 151780 220496 151782 220516
rect 151450 220360 151506 220416
rect 150898 220088 150954 220144
rect 151082 220088 151138 220144
rect 151910 220088 151966 220144
rect 156694 229900 156750 229936
rect 156694 229880 156696 229900
rect 156696 229880 156748 229900
rect 156748 229880 156750 229900
rect 156694 227432 156750 227488
rect 157430 229880 157486 229936
rect 157062 229356 157118 229392
rect 157062 229336 157064 229356
rect 157064 229336 157116 229356
rect 157116 229336 157118 229356
rect 156786 223080 156842 223136
rect 156970 220516 157026 220552
rect 156970 220496 156972 220516
rect 156972 220496 157024 220516
rect 157024 220496 157026 220516
rect 158350 220904 158406 220960
rect 160006 228112 160062 228168
rect 161938 221604 161994 221640
rect 161938 221584 161940 221604
rect 161940 221584 161992 221604
rect 161992 221584 161994 221604
rect 164330 221584 164386 221640
rect 166814 228812 166870 228848
rect 166814 228792 166816 228812
rect 166816 228792 166868 228812
rect 166868 228792 166870 228812
rect 166814 228404 166870 228440
rect 166814 228384 166816 228404
rect 166816 228384 166868 228404
rect 166868 228384 166870 228404
rect 166814 228112 166870 228168
rect 166538 227432 166594 227488
rect 169298 228948 169354 228984
rect 169298 228928 169300 228948
rect 169300 228928 169352 228948
rect 169352 228928 169354 228948
rect 169114 228792 169170 228848
rect 169482 227316 169538 227352
rect 169482 227296 169484 227316
rect 169484 227296 169536 227316
rect 169536 227296 169538 227316
rect 166722 220904 166778 220960
rect 166906 220904 166962 220960
rect 166906 220224 166962 220280
rect 167090 220224 167146 220280
rect 171230 227568 171286 227624
rect 172150 228928 172206 228984
rect 172334 228384 172390 228440
rect 172150 227568 172206 227624
rect 171690 227296 171746 227352
rect 171046 218612 171102 218648
rect 171046 218592 171048 218612
rect 171048 218592 171100 218612
rect 171100 218592 171102 218612
rect 173162 228792 173218 228848
rect 174818 228812 174874 228848
rect 174818 228792 174820 228812
rect 174820 228792 174872 228812
rect 174872 228792 174874 228812
rect 172886 218592 172942 218648
rect 175462 220904 175518 220960
rect 176474 221332 176530 221368
rect 176474 221312 176476 221332
rect 176476 221312 176528 221332
rect 176528 221312 176530 221332
rect 177302 221312 177358 221368
rect 176474 220788 176530 220824
rect 176474 220768 176476 220788
rect 176476 220768 176528 220788
rect 176528 220768 176530 220788
rect 179878 220768 179934 220824
rect 180522 220088 180578 220144
rect 184662 221720 184718 221776
rect 185766 221740 185822 221776
rect 185766 221720 185768 221740
rect 185768 221720 185820 221740
rect 185820 221720 185822 221740
rect 185766 220088 185822 220144
rect 202602 226208 202658 226264
rect 202418 219816 202474 219872
rect 203154 219816 203210 219872
rect 205086 226244 205088 226264
rect 205088 226244 205140 226264
rect 205140 226244 205142 226264
rect 205086 226208 205142 226244
rect 219622 228656 219678 228712
rect 220542 228676 220598 228712
rect 220542 228656 220544 228676
rect 220544 228656 220596 228676
rect 220596 228656 220598 228676
rect 486974 219408 487030 219464
rect 487802 218048 487858 218104
rect 490378 218592 490434 218648
rect 492678 218864 492734 218920
rect 488676 217096 488732 217152
rect 493782 218864 493838 218920
rect 493782 217232 493838 217288
rect 494702 218864 494758 218920
rect 495346 217232 495402 217288
rect 497830 220904 497886 220960
rect 497462 218592 497518 218648
rect 498566 217232 498622 217288
rect 505650 217504 505706 217560
rect 508502 217776 508558 217832
rect 510158 217776 510214 217832
rect 513378 221604 513434 221640
rect 513378 221584 513380 221604
rect 513380 221584 513432 221604
rect 513432 221584 513434 221604
rect 515218 219680 515274 219736
rect 520186 221176 520242 221232
rect 522578 217776 522634 217832
rect 540886 221992 540942 222048
rect 543094 221720 543150 221776
rect 543830 221992 543886 222048
rect 544198 221992 544254 222048
rect 544014 221720 544070 221776
rect 546590 221992 546646 222048
rect 547142 221856 547198 221912
rect 554502 244704 554558 244760
rect 554502 240352 554558 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 557078 224748 557080 224768
rect 557080 224748 557132 224768
rect 557132 224748 557134 224768
rect 557078 224712 557134 224748
rect 552938 222128 552994 222184
rect 553582 222128 553638 222184
rect 552846 220224 552902 220280
rect 553950 220380 554006 220416
rect 553950 220360 553952 220380
rect 553952 220360 554004 220380
rect 554004 220360 554006 220380
rect 553214 219136 553270 219192
rect 555698 217776 555754 217832
rect 557906 222264 557962 222320
rect 558550 221856 558606 221912
rect 559562 221992 559618 222048
rect 561678 224712 561734 224768
rect 560206 219136 560262 219192
rect 563150 222264 563206 222320
rect 562874 221992 562930 222048
rect 562690 221756 562692 221776
rect 562692 221756 562744 221776
rect 562744 221756 562746 221776
rect 562690 221720 562746 221756
rect 563150 220632 563206 220688
rect 563334 220360 563390 220416
rect 562874 219952 562930 220008
rect 562690 217776 562746 217832
rect 562874 217776 562930 217832
rect 563518 219952 563574 220008
rect 563518 217776 563574 217832
rect 564806 220632 564862 220688
rect 565634 220360 565690 220416
rect 564806 219952 564862 220008
rect 567106 219136 567162 219192
rect 566922 217776 566978 217832
rect 568946 221720 569002 221776
rect 568302 219136 568358 219192
rect 569958 220380 570014 220416
rect 569958 220360 569960 220380
rect 569960 220360 570012 220380
rect 570012 220360 570014 220380
rect 572994 220496 573050 220552
rect 572626 220360 572682 220416
rect 572810 220360 572866 220416
rect 573362 220224 573418 220280
rect 572534 219952 572590 220008
rect 572994 220088 573050 220144
rect 572074 217776 572130 217832
rect 574098 217776 574154 217832
rect 574098 216688 574154 216744
rect 574834 217776 574890 217832
rect 574650 216688 574706 216744
rect 650642 256672 650698 256728
rect 589646 220496 589702 220552
rect 586334 220224 586390 220280
rect 586334 219988 586336 220008
rect 586336 219988 586388 220008
rect 586388 219988 586390 220008
rect 586334 219952 586390 219988
rect 589462 219952 589518 220008
rect 578882 213968 578938 214024
rect 578514 211656 578570 211712
rect 579526 209788 579528 209808
rect 579528 209788 579580 209808
rect 579580 209788 579582 209808
rect 579526 209752 579582 209788
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 598938 221448 598994 221504
rect 594798 218320 594854 218376
rect 595166 217504 595222 217560
rect 596362 217232 596418 217288
rect 595718 216960 595774 217016
rect 598478 215872 598534 215928
rect 600778 217096 600834 217152
rect 601514 217132 601516 217152
rect 601516 217132 601568 217152
rect 601568 217132 601570 217152
rect 601514 217096 601570 217132
rect 603354 218592 603410 218648
rect 611634 219408 611690 219464
rect 618258 221176 618314 221232
rect 617246 219680 617302 219736
rect 618902 215328 618958 215384
rect 627458 218048 627514 218104
rect 627918 216144 627974 216200
rect 631322 220904 631378 220960
rect 631138 218592 631194 218648
rect 650642 222808 650698 222864
rect 649906 221448 649962 221504
rect 644754 220360 644810 220416
rect 648526 218592 648582 218648
rect 651470 221720 651526 221776
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153992 578386 154048
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147464 579582 147520
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 578882 136584 578938 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578882 129648 578938 129704
rect 579526 127880 579582 127936
rect 578330 125296 578386 125352
rect 578698 123528 578754 123584
rect 578882 121352 578938 121408
rect 578514 118360 578570 118416
rect 578330 108296 578386 108352
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579526 112512 579582 112568
rect 579342 110064 579398 110120
rect 579066 105848 579122 105904
rect 578514 103128 578570 103184
rect 579158 101632 579214 101688
rect 578606 97416 578662 97472
rect 578330 94968 578386 95024
rect 579526 99220 579528 99240
rect 579528 99220 579580 99240
rect 579580 99220 579582 99240
rect 579526 99184 579582 99220
rect 579250 93064 579306 93120
rect 578606 90888 578662 90944
rect 579250 88032 579306 88088
rect 578330 86400 578386 86456
rect 579250 83988 579252 84008
rect 579252 83988 579304 84008
rect 579304 83988 579306 84008
rect 579250 83952 579306 83988
rect 578882 82184 578938 82240
rect 578238 77832 578294 77888
rect 579434 80008 579490 80064
rect 652574 283192 652630 283248
rect 656162 271088 656218 271144
rect 652574 229744 652630 229800
rect 654782 226344 654838 226400
rect 653402 225256 653458 225312
rect 653034 220632 653090 220688
rect 652850 215872 652906 215928
rect 656162 225528 656218 225584
rect 655426 218864 655482 218920
rect 657726 224984 657782 225040
rect 657542 223896 657598 223952
rect 656806 217232 656862 217288
rect 656530 213152 656586 213208
rect 664442 311888 664498 311944
rect 662418 293800 662474 293856
rect 668122 283872 668178 283928
rect 665822 268504 665878 268560
rect 664442 247968 664498 248024
rect 659106 222536 659162 222592
rect 658738 214512 658794 214568
rect 662050 217504 662106 217560
rect 661498 213424 661554 213480
rect 663706 229336 663762 229392
rect 664442 223760 664498 223816
rect 665822 230424 665878 230480
rect 665178 229064 665234 229120
rect 665546 216144 665602 216200
rect 667018 221040 667074 221096
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589462 204720 589518 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 667018 176432 667074 176488
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589646 170448 589702 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 580446 77832 580502 77888
rect 579250 75656 579306 75712
rect 578514 71168 578570 71224
rect 579526 73108 579528 73128
rect 579528 73108 579580 73128
rect 579580 73108 579582 73128
rect 579526 73072 579582 73108
rect 579526 66852 579528 66872
rect 579528 66852 579580 66872
rect 579580 66852 579582 66872
rect 579526 66816 579582 66852
rect 579526 64504 579582 64560
rect 579526 61784 579582 61840
rect 578882 60424 578938 60480
rect 574466 54712 574522 54768
rect 576122 54984 576178 55040
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 578330 56072 578386 56128
rect 577502 54168 577558 54224
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590382 134544 590438 134600
rect 589462 132912 589518 132968
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 588726 129648 588782 129704
rect 588542 103536 588598 103592
rect 589462 128016 589518 128072
rect 590106 126384 590162 126440
rect 589462 123120 589518 123176
rect 590566 124752 590622 124808
rect 589278 121508 589334 121544
rect 589278 121488 589280 121508
rect 589280 121488 589332 121508
rect 589332 121488 589334 121508
rect 589646 119856 589702 119912
rect 589462 116592 589518 116648
rect 590106 118224 590162 118280
rect 589462 113328 589518 113384
rect 668030 221720 668086 221776
rect 667846 220632 667902 220688
rect 668030 219680 668086 219736
rect 667754 219408 667810 219464
rect 667386 134544 667442 134600
rect 668030 213152 668086 213208
rect 668030 207576 668086 207632
rect 668030 204040 668086 204096
rect 667938 199144 667994 199200
rect 667938 194112 667994 194168
rect 667938 189624 667994 189680
rect 668030 184320 668086 184376
rect 668030 179424 668086 179480
rect 667754 174936 667810 174992
rect 667570 133320 667626 133376
rect 668214 173032 668270 173088
rect 668398 169632 668454 169688
rect 668214 164872 668270 164928
rect 668214 163276 668216 163296
rect 668216 163276 668268 163296
rect 668268 163276 668270 163296
rect 668214 163240 668270 163276
rect 668214 160012 668216 160032
rect 668216 160012 668268 160032
rect 668268 160012 668270 160032
rect 668214 159976 668270 160012
rect 668582 158344 668638 158400
rect 668306 155116 668308 155136
rect 668308 155116 668360 155136
rect 668360 155116 668362 155136
rect 668306 155080 668362 155116
rect 668214 148552 668270 148608
rect 668214 135496 668270 135552
rect 669042 223760 669098 223816
rect 669042 222536 669098 222592
rect 670606 392264 670662 392320
rect 669962 345616 670018 345672
rect 669410 174664 669466 174720
rect 669410 171944 669466 172000
rect 669778 234232 669834 234288
rect 669410 148960 669466 149016
rect 669226 143656 669282 143712
rect 668950 138760 669006 138816
rect 670422 261296 670478 261352
rect 670238 259664 670294 259720
rect 670422 247152 670478 247208
rect 670238 245520 670294 245576
rect 670422 233960 670478 234016
rect 671986 372544 672042 372600
rect 673182 401240 673238 401296
rect 672998 394712 673054 394768
rect 672998 380976 673054 381032
rect 672814 357448 672870 357504
rect 672354 357040 672410 357096
rect 672170 355408 672226 355464
rect 671986 350104 672042 350160
rect 671986 332288 672042 332344
rect 673366 400560 673422 400616
rect 673182 356768 673238 356824
rect 672538 356224 672594 356280
rect 672354 312432 672410 312488
rect 673918 399744 673974 399800
rect 673734 393080 673790 393136
rect 673734 376624 673790 376680
rect 673366 355816 673422 355872
rect 674378 396480 674434 396536
rect 676586 402872 676642 402928
rect 676034 402600 676090 402656
rect 674838 402192 674894 402248
rect 674838 401648 674894 401704
rect 676586 400832 676642 400888
rect 674838 399336 674894 399392
rect 676218 398384 676274 398440
rect 675022 398112 675078 398168
rect 674746 395664 674802 395720
rect 674562 395256 674618 395312
rect 674286 394440 674342 394496
rect 681002 397568 681058 397624
rect 676034 394032 676090 394088
rect 676034 393080 676090 393136
rect 683026 392672 683082 392728
rect 683026 389816 683082 389872
rect 681002 388456 681058 388512
rect 675390 386008 675446 386064
rect 675758 385328 675814 385384
rect 675758 381656 675814 381712
rect 675390 380976 675446 381032
rect 675758 378664 675814 378720
rect 675758 377304 675814 377360
rect 675114 376624 675170 376680
rect 675758 373632 675814 373688
rect 675666 372952 675722 373008
rect 675114 372544 675170 372600
rect 675574 358264 675630 358320
rect 673918 355000 673974 355056
rect 674102 354592 674158 354648
rect 673734 352552 673790 352608
rect 672998 351328 673054 351384
rect 672722 348472 672778 348528
rect 672538 311616 672594 311672
rect 672170 310800 672226 310856
rect 672538 304272 672594 304328
rect 671526 302232 671582 302288
rect 671342 258440 671398 258496
rect 670790 256400 670846 256456
rect 670974 250824 671030 250880
rect 670974 247968 671030 248024
rect 673366 349696 673422 349752
rect 672998 337184 673054 337240
rect 673550 349288 673606 349344
rect 673366 335552 673422 335608
rect 673918 348880 673974 348936
rect 673734 333920 673790 333976
rect 673550 332696 673606 332752
rect 673918 331200 673974 331256
rect 674746 354184 674802 354240
rect 674286 350920 674342 350976
rect 674562 350512 674618 350568
rect 675942 357856 675998 357912
rect 675942 356496 675998 356552
rect 675850 353776 675906 353832
rect 675574 352824 675630 352880
rect 675850 351872 675906 351928
rect 676034 351736 676090 351792
rect 683118 347656 683174 347712
rect 676034 347248 676090 347304
rect 676494 346568 676550 346624
rect 683118 346432 683174 346488
rect 676034 345616 676090 345672
rect 675574 340720 675630 340776
rect 675758 340176 675814 340232
rect 675114 338680 675170 338736
rect 675666 337728 675722 337784
rect 675114 337184 675170 337240
rect 675114 335552 675170 335608
rect 675114 333920 675170 333976
rect 675114 332696 675170 332752
rect 675114 332288 675170 332344
rect 675114 331200 675170 331256
rect 675758 328344 675814 328400
rect 673366 312704 673422 312760
rect 673182 311208 673238 311264
rect 672998 305496 673054 305552
rect 672538 287816 672594 287872
rect 671894 262112 671950 262168
rect 671710 260888 671766 260944
rect 671710 246880 671766 246936
rect 671158 224712 671214 224768
rect 671250 224168 671306 224224
rect 671250 223796 671252 223816
rect 671252 223796 671304 223816
rect 671304 223796 671306 223816
rect 671250 223760 671306 223796
rect 672078 246200 672134 246256
rect 672998 285504 673054 285560
rect 672814 283872 672870 283928
rect 674194 310392 674250 310448
rect 674010 303864 674066 303920
rect 673642 303456 673698 303512
rect 673366 267416 673422 267472
rect 673182 266600 673238 266656
rect 673366 260480 673422 260536
rect 673182 258848 673238 258904
rect 671894 232484 671950 232520
rect 671894 232464 671896 232484
rect 671896 232464 671948 232484
rect 671948 232464 671950 232484
rect 671894 231532 671950 231568
rect 671894 231512 671896 231532
rect 671896 231512 671948 231532
rect 671948 231512 671950 231532
rect 672262 226072 672318 226128
rect 672262 225684 672318 225720
rect 672262 225664 672264 225684
rect 672264 225664 672316 225684
rect 672316 225664 672318 225684
rect 672078 225392 672134 225448
rect 672262 225256 672318 225312
rect 672032 225140 672088 225176
rect 672032 225120 672034 225140
rect 672034 225120 672086 225140
rect 672086 225120 672088 225140
rect 673182 241032 673238 241088
rect 674010 286456 674066 286512
rect 673918 267008 673974 267064
rect 673366 240216 673422 240272
rect 673090 236680 673146 236736
rect 672722 226380 672724 226400
rect 672724 226380 672776 226400
rect 672776 226380 672778 226400
rect 672722 226344 672778 226380
rect 672630 225800 672686 225856
rect 671818 224440 671874 224496
rect 671020 223388 671022 223408
rect 671022 223388 671074 223408
rect 671074 223388 671076 223408
rect 671020 223352 671076 223388
rect 671158 223080 671214 223136
rect 670790 210432 670846 210488
rect 670790 209888 670846 209944
rect 670790 193160 670846 193216
rect 670606 170992 670662 171048
rect 670606 170312 670662 170368
rect 671342 219680 671398 219736
rect 671158 177928 671214 177984
rect 670606 147600 670662 147656
rect 672078 223760 672134 223816
rect 672078 219000 672134 219056
rect 671894 216552 671950 216608
rect 671894 204448 671950 204504
rect 672722 224712 672778 224768
rect 672446 223352 672502 223408
rect 672722 222808 672778 222864
rect 672630 220224 672686 220280
rect 672446 217232 672502 217288
rect 672538 213696 672594 213752
rect 672722 213288 672778 213344
rect 672538 196288 672594 196344
rect 672262 180240 672318 180296
rect 672354 176024 672410 176080
rect 671986 170720 672042 170776
rect 672170 169088 672226 169144
rect 671986 154400 672042 154456
rect 672170 153040 672226 153096
rect 671710 150184 671766 150240
rect 671526 145288 671582 145344
rect 669226 133728 669282 133784
rect 669226 132640 669282 132696
rect 668950 131144 669006 131200
rect 668766 130600 668822 130656
rect 668582 128968 668638 129024
rect 668582 127744 668638 127800
rect 668030 125296 668086 125352
rect 667202 116048 667258 116104
rect 590290 114960 590346 115016
rect 589462 111696 589518 111752
rect 589462 110064 589518 110120
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589830 105168 589886 105224
rect 668214 111016 668270 111072
rect 666650 109316 666706 109372
rect 667938 107752 667994 107808
rect 668122 106120 668178 106176
rect 589462 101904 589518 101960
rect 591302 54440 591358 54496
rect 625434 94424 625490 94480
rect 635554 96872 635610 96928
rect 635738 95920 635794 95976
rect 637026 96872 637082 96928
rect 641994 96464 642050 96520
rect 645582 96076 645638 96112
rect 645582 96056 645584 96076
rect 645584 96056 645636 96076
rect 645636 96056 645638 96076
rect 645766 95512 645822 95568
rect 647514 96076 647570 96112
rect 647514 96056 647516 96076
rect 647516 96056 647568 96076
rect 647568 96056 647570 96076
rect 647514 95512 647570 95568
rect 647330 94968 647386 95024
rect 626354 93608 626410 93664
rect 626170 92792 626226 92848
rect 625802 91976 625858 92032
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 647698 89800 647754 89856
rect 626262 89528 626318 89584
rect 626446 88712 626502 88768
rect 624974 88304 625030 88360
rect 626262 88304 626318 88360
rect 626446 87896 626502 87952
rect 626262 87080 626318 87136
rect 648802 91976 648858 92032
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 626446 85484 626448 85504
rect 626448 85484 626500 85504
rect 626500 85484 626502 85504
rect 626446 85448 626502 85484
rect 625250 84632 625306 84688
rect 648618 84632 648674 84688
rect 626446 83816 626502 83872
rect 628746 83272 628802 83328
rect 650550 87080 650606 87136
rect 654322 94152 654378 94208
rect 654690 93336 654746 93392
rect 655426 91432 655482 91488
rect 655426 90616 655482 90672
rect 655794 89800 655850 89856
rect 663798 93064 663854 93120
rect 663982 91704 664038 91760
rect 664350 90616 664406 90672
rect 664534 89800 664590 89856
rect 665362 93336 665418 93392
rect 665178 88984 665234 89040
rect 650274 82184 650330 82240
rect 629206 81640 629262 81696
rect 623042 77288 623098 77344
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 77560 639658 77616
rect 646502 74160 646558 74216
rect 646686 71712 646742 71768
rect 646318 69128 646374 69184
rect 646134 67088 646190 67144
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 129094 44276 129096 44296
rect 129096 44276 129148 44296
rect 129148 44276 129150 44296
rect 129094 44240 129150 44276
rect 470322 53644 470378 53680
rect 470322 53624 470324 53644
rect 470324 53624 470376 53644
rect 470376 53624 470378 53644
rect 471978 53644 472034 53680
rect 471978 53624 471980 53644
rect 471980 53624 472032 53644
rect 472032 53624 472034 53644
rect 463882 53080 463938 53136
rect 470966 53352 471022 53408
rect 471150 53080 471206 53136
rect 476762 53352 476818 53408
rect 308034 50224 308090 50280
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 131946 44240 132002 44296
rect 458362 46688 458418 46744
rect 458178 44376 458234 44432
rect 142618 44240 142674 44296
rect 307298 44104 307354 44160
rect 194322 42064 194378 42120
rect 419722 43560 419778 43616
rect 440238 43596 440240 43616
rect 440240 43596 440292 43616
rect 440292 43596 440294 43616
rect 440238 43560 440294 43596
rect 441066 43596 441068 43616
rect 441068 43596 441120 43616
rect 441120 43596 441122 43616
rect 441066 43560 441122 43596
rect 416594 42336 416650 42392
rect 404634 42064 404690 42120
rect 405186 42064 405242 42120
rect 415582 42064 415638 42120
rect 310426 41792 310482 41848
rect 311070 41792 311126 41848
rect 361946 41792 362002 41848
rect 365166 41792 365222 41848
rect 461030 44376 461086 44432
rect 460846 43832 460902 43888
rect 461766 42880 461822 42936
rect 462870 43560 462926 43616
rect 462686 43152 462742 43208
rect 463698 44376 463754 44432
rect 549994 48864 550050 48920
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 465078 46688 465134 46744
rect 647514 78104 647570 78160
rect 647330 64368 647386 64424
rect 648986 62056 649042 62112
rect 648618 59200 648674 59256
rect 647514 57296 647570 57352
rect 661590 48454 661646 48510
rect 661774 47733 661830 47789
rect 667938 102720 667994 102776
rect 668306 104760 668362 104816
rect 668306 104352 668362 104408
rect 668766 119992 668822 120048
rect 669962 130872 670018 130928
rect 669226 125976 669282 126032
rect 669226 124072 669282 124128
rect 668950 119176 669006 119232
rect 669226 117000 669282 117056
rect 669226 114280 669282 114336
rect 672170 131688 672226 131744
rect 672538 175616 672594 175672
rect 672538 168272 672594 168328
rect 672354 131416 672410 131472
rect 672538 131144 672594 131200
rect 671986 126792 672042 126848
rect 671526 122712 671582 122768
rect 670698 121352 670754 121408
rect 671526 112648 671582 112704
rect 668766 104760 668822 104816
rect 668582 102720 668638 102776
rect 673274 234912 673330 234968
rect 675298 325488 675354 325544
rect 675114 325216 675170 325272
rect 676218 313928 676274 313984
rect 674654 312976 674710 313032
rect 674838 312704 674894 312760
rect 674838 312024 674894 312080
rect 674654 311888 674710 311944
rect 674378 309984 674434 310040
rect 674562 309576 674618 309632
rect 674378 305088 674434 305144
rect 674378 283464 674434 283520
rect 674378 267824 674434 267880
rect 674378 266192 674434 266248
rect 674194 265784 674250 265840
rect 674102 265376 674158 265432
rect 675850 309304 675906 309360
rect 676034 308352 676090 308408
rect 675114 307944 675170 308000
rect 674930 301824 674986 301880
rect 676034 307536 676090 307592
rect 676034 304680 676090 304736
rect 675850 301824 675906 301880
rect 676494 305904 676550 305960
rect 676494 301552 676550 301608
rect 676034 300600 676090 300656
rect 679622 306720 679678 306776
rect 677598 306312 677654 306368
rect 683026 302640 683082 302696
rect 683026 299376 683082 299432
rect 676126 296792 676182 296848
rect 675942 296520 675998 296576
rect 675574 295296 675630 295352
rect 675758 294480 675814 294536
rect 675206 293800 675262 293856
rect 675574 292168 675630 292224
rect 675758 291488 675814 291544
rect 675758 290808 675814 290864
rect 675114 287816 675170 287872
rect 675390 286456 675446 286512
rect 675114 285504 675170 285560
rect 675666 283600 675722 283656
rect 675666 282784 675722 282840
rect 675758 281152 675814 281208
rect 683118 271088 683174 271144
rect 683118 268504 683174 268560
rect 674562 264968 674618 265024
rect 674654 264560 674710 264616
rect 674286 262520 674342 262576
rect 674286 243616 674342 243672
rect 674102 241848 674158 241904
rect 674378 241576 674434 241632
rect 673918 236680 673974 236736
rect 673458 229064 673514 229120
rect 673458 227024 673514 227080
rect 673458 226788 673460 226808
rect 673460 226788 673512 226808
rect 673512 226788 673514 226808
rect 673458 226752 673514 226788
rect 673366 224712 673422 224768
rect 673458 224168 673514 224224
rect 673458 216008 673514 216064
rect 673182 215736 673238 215792
rect 681002 263200 681058 263256
rect 676218 262792 676274 262848
rect 674746 259256 674802 259312
rect 675298 254904 675354 254960
rect 675022 254632 675078 254688
rect 675022 249192 675078 249248
rect 676218 257080 676274 257136
rect 676218 256400 676274 256456
rect 683026 257488 683082 257544
rect 681002 254904 681058 254960
rect 676034 254632 676090 254688
rect 675482 250824 675538 250880
rect 675758 250144 675814 250200
rect 675390 249464 675446 249520
rect 675298 247152 675354 247208
rect 675206 246880 675262 246936
rect 675206 245520 675262 245576
rect 675206 243616 675262 243672
rect 675758 242256 675814 242312
rect 675390 241032 675446 241088
rect 675390 240216 675446 240272
rect 674562 235184 674618 235240
rect 674838 234640 674894 234696
rect 674102 233844 674158 233880
rect 674102 233824 674104 233844
rect 674104 233824 674156 233844
rect 674156 233824 674158 233844
rect 673642 215192 673698 215248
rect 673642 214920 673698 214976
rect 673090 201320 673146 201376
rect 673642 200504 673698 200560
rect 674102 228520 674158 228576
rect 674102 226752 674158 226808
rect 675850 235184 675906 235240
rect 674674 230444 674730 230480
rect 674674 230424 674676 230444
rect 674676 230424 674728 230444
rect 674728 230424 674730 230444
rect 674838 230424 674894 230480
rect 674470 229336 674526 229392
rect 674838 226072 674894 226128
rect 674378 222264 674434 222320
rect 675022 225800 675078 225856
rect 674838 221448 674894 221504
rect 675206 225256 675262 225312
rect 675022 220496 675078 220552
rect 676034 233844 676090 233880
rect 676034 233824 676036 233844
rect 676036 233824 676088 233844
rect 676088 233824 676090 233844
rect 675850 232500 675852 232520
rect 675852 232500 675904 232520
rect 675904 232500 675906 232520
rect 675850 232464 675906 232500
rect 675850 231532 675906 231568
rect 675850 231512 675852 231532
rect 675852 231512 675904 231532
rect 675904 231512 675906 231532
rect 676678 230424 676734 230480
rect 676034 230152 676090 230208
rect 675114 218592 675170 218648
rect 675022 217776 675078 217832
rect 674654 216960 674710 217016
rect 674378 216280 674434 216336
rect 674378 215464 674434 215520
rect 674102 213968 674158 214024
rect 674010 212744 674066 212800
rect 672906 177656 672962 177712
rect 673366 176840 673422 176896
rect 673182 167864 673238 167920
rect 673090 166912 673146 166968
rect 672906 165552 672962 165608
rect 672722 125976 672778 126032
rect 672722 123936 672778 123992
rect 674102 209616 674158 209672
rect 673918 177248 673974 177304
rect 673918 168680 673974 168736
rect 673734 153312 673790 153368
rect 673918 151000 673974 151056
rect 673366 132096 673422 132152
rect 673734 123528 673790 123584
rect 673550 123120 673606 123176
rect 673366 120672 673422 120728
rect 673090 117544 673146 117600
rect 672906 115776 672962 115832
rect 672722 106528 672778 106584
rect 672354 106120 672410 106176
rect 673550 117000 673606 117056
rect 674838 216144 674894 216200
rect 674470 214104 674526 214160
rect 674470 200776 674526 200832
rect 676402 228520 676458 228576
rect 676034 221448 676090 221504
rect 676034 219000 676090 219056
rect 675574 217504 675630 217560
rect 675942 215500 675944 215520
rect 675944 215500 675996 215520
rect 675996 215500 675998 215520
rect 675942 215464 675998 215500
rect 677046 227024 677102 227080
rect 675942 214648 675998 214704
rect 675850 212064 675906 212120
rect 675850 209616 675906 209672
rect 678242 223760 678298 223816
rect 683210 222672 683266 222728
rect 683578 223080 683634 223136
rect 683394 219816 683450 219872
rect 683302 218592 683358 218648
rect 683118 212880 683174 212936
rect 678978 211384 679034 211440
rect 680358 210568 680414 210624
rect 683302 210296 683358 210352
rect 678978 207576 679034 207632
rect 676862 206896 676918 206952
rect 675758 205536 675814 205592
rect 675114 204448 675170 204504
rect 675758 204176 675814 204232
rect 675114 201320 675170 201376
rect 675298 200776 675354 200832
rect 675114 200504 675170 200560
rect 675758 200640 675814 200696
rect 675758 198328 675814 198384
rect 675114 196288 675170 196344
rect 675298 195744 675354 195800
rect 675114 193160 675170 193216
rect 675666 192616 675722 192672
rect 676862 189624 676918 189680
rect 674286 178064 674342 178120
rect 674654 175208 674710 175264
rect 674378 174392 674434 174448
rect 675206 173984 675262 174040
rect 674838 169360 674894 169416
rect 676034 173168 676090 173224
rect 675390 171128 675446 171184
rect 675942 169360 675998 169416
rect 676586 169904 676642 169960
rect 675850 167864 675906 167920
rect 676034 167048 676090 167104
rect 674838 160520 674894 160576
rect 675850 166912 675906 166968
rect 678242 171536 678298 171592
rect 676586 166368 676642 166424
rect 676862 166368 676918 166424
rect 676034 165552 676090 165608
rect 675482 161336 675538 161392
rect 675482 160520 675538 160576
rect 675022 159432 675078 159488
rect 675482 159432 675538 159488
rect 675758 156984 675814 157040
rect 675758 155624 675814 155680
rect 675114 154400 675170 154456
rect 675114 153040 675170 153096
rect 675666 153040 675722 153096
rect 675758 151408 675814 151464
rect 675114 151000 675170 151056
rect 675298 148960 675354 149016
rect 675114 147600 675170 147656
rect 675758 148416 675814 148472
rect 675666 147600 675722 147656
rect 676034 134544 676090 134600
rect 676034 132504 676090 132560
rect 674654 130464 674710 130520
rect 676218 130192 676274 130248
rect 674378 129648 674434 129704
rect 674286 129240 674342 129296
rect 674102 120400 674158 120456
rect 675206 128832 675262 128888
rect 674470 125568 674526 125624
rect 674286 119992 674342 120048
rect 674654 124752 674710 124808
rect 674470 111288 674526 111344
rect 676678 128152 676734 128208
rect 676218 127744 676274 127800
rect 676402 127744 676458 127800
rect 675942 125316 675998 125352
rect 675942 125296 675944 125316
rect 675944 125296 675996 125316
rect 675996 125296 675998 125316
rect 676126 125296 676182 125352
rect 676678 126112 676734 126168
rect 683118 126112 683174 126168
rect 676862 125704 676918 125760
rect 676586 125316 676642 125352
rect 676586 125296 676588 125316
rect 676588 125296 676640 125316
rect 676640 125296 676642 125316
rect 676126 120672 676182 120728
rect 675298 118496 675354 118552
rect 675850 118496 675906 118552
rect 675022 116320 675078 116376
rect 674838 114280 674894 114336
rect 678978 125296 679034 125352
rect 677598 122032 677654 122088
rect 675850 116320 675906 116376
rect 683118 122848 683174 122904
rect 678978 121624 679034 121680
rect 675482 116048 675538 116104
rect 677598 116048 677654 116104
rect 675390 114280 675446 114336
rect 675758 114280 675814 114336
rect 675758 112376 675814 112432
rect 675390 111288 675446 111344
rect 675758 110336 675814 110392
rect 675666 108024 675722 108080
rect 675114 106528 675170 106584
rect 673366 104488 673422 104544
rect 675114 104488 675170 104544
rect 675758 103128 675814 103184
rect 675666 102584 675722 102640
rect 671986 99320 672042 99376
rect 675298 99320 675354 99376
rect 662418 47368 662474 47424
rect 464710 44512 464766 44568
rect 463882 44104 463938 44160
rect 471058 43832 471114 43888
rect 465814 43152 465870 43208
rect 463974 42880 464030 42936
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 461950 41792 462006 41848
rect 458178 41112 458234 41168
rect 141698 40296 141754 40352
<< metal3 >>
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 675845 896746 675911 896749
rect 675845 896744 676292 896746
rect 675845 896688 675850 896744
rect 675906 896688 676292 896744
rect 675845 896686 676292 896688
rect 675845 896683 675911 896686
rect 676029 896338 676095 896341
rect 676029 896336 676292 896338
rect 676029 896280 676034 896336
rect 676090 896280 676292 896336
rect 676029 896278 676292 896280
rect 676029 896275 676095 896278
rect 675845 895522 675911 895525
rect 675845 895520 676292 895522
rect 675845 895464 675850 895520
rect 675906 895464 676292 895520
rect 675845 895462 676292 895464
rect 675845 895459 675911 895462
rect 676029 894706 676095 894709
rect 676029 894704 676292 894706
rect 676029 894648 676034 894704
rect 676090 894648 676292 894704
rect 676029 894646 676292 894648
rect 676029 894643 676095 894646
rect 675845 893890 675911 893893
rect 675845 893888 676292 893890
rect 675845 893832 675850 893888
rect 675906 893832 676292 893888
rect 675845 893830 676292 893832
rect 675845 893827 675911 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 676029 892666 676095 892669
rect 676029 892664 676292 892666
rect 676029 892608 676034 892664
rect 676090 892608 676292 892664
rect 676029 892606 676292 892608
rect 676029 892603 676095 892606
rect 675886 892196 675892 892260
rect 675956 892258 675962 892260
rect 675956 892198 676292 892258
rect 675956 892196 675962 892198
rect 679617 891850 679683 891853
rect 679604 891848 679683 891850
rect 679604 891792 679622 891848
rect 679678 891792 679683 891848
rect 679604 891790 679683 891792
rect 679617 891787 679683 891790
rect 676029 891442 676095 891445
rect 676029 891440 676292 891442
rect 676029 891384 676034 891440
rect 676090 891384 676292 891440
rect 676029 891382 676292 891384
rect 676029 891379 676095 891382
rect 675201 891034 675267 891037
rect 675201 891032 676292 891034
rect 675201 890976 675206 891032
rect 675262 890976 676292 891032
rect 675201 890974 676292 890976
rect 675201 890971 675267 890974
rect 680997 890626 681063 890629
rect 680997 890624 681076 890626
rect 680997 890568 681002 890624
rect 681058 890568 681076 890624
rect 680997 890566 681076 890568
rect 680997 890563 681063 890566
rect 676029 890218 676095 890221
rect 676029 890216 676292 890218
rect 676029 890160 676034 890216
rect 676090 890160 676292 890216
rect 676029 890158 676292 890160
rect 676029 890155 676095 890158
rect 678237 889810 678303 889813
rect 678237 889808 678316 889810
rect 678237 889752 678242 889808
rect 678298 889752 678316 889808
rect 678237 889750 678316 889752
rect 678237 889747 678303 889750
rect 676029 889402 676095 889405
rect 676029 889400 676292 889402
rect 676029 889344 676034 889400
rect 676090 889344 676292 889400
rect 676029 889342 676292 889344
rect 676029 889339 676095 889342
rect 676029 888994 676095 888997
rect 676029 888992 676292 888994
rect 676029 888936 676034 888992
rect 676090 888936 676292 888992
rect 676029 888934 676292 888936
rect 676029 888931 676095 888934
rect 674741 888586 674807 888589
rect 674741 888584 676292 888586
rect 674741 888528 674746 888584
rect 674802 888528 676292 888584
rect 674741 888526 676292 888528
rect 674741 888523 674807 888526
rect 683113 888178 683179 888181
rect 683100 888176 683179 888178
rect 683100 888120 683118 888176
rect 683174 888120 683179 888176
rect 683100 888118 683179 888120
rect 683113 888115 683179 888118
rect 675886 887708 675892 887772
rect 675956 887770 675962 887772
rect 675956 887710 676292 887770
rect 675956 887708 675962 887710
rect 676029 887362 676095 887365
rect 676029 887360 676292 887362
rect 676029 887304 676034 887360
rect 676090 887304 676292 887360
rect 676029 887302 676292 887304
rect 676029 887299 676095 887302
rect 676029 886954 676095 886957
rect 676029 886952 676292 886954
rect 676029 886896 676034 886952
rect 676090 886896 676292 886952
rect 676029 886894 676292 886896
rect 676029 886891 676095 886894
rect 683070 886138 683130 886516
rect 675894 886108 683130 886138
rect 675894 886078 683100 886108
rect 675702 885804 675708 885868
rect 675772 885866 675778 885868
rect 675894 885866 675954 886078
rect 675772 885806 675954 885866
rect 675772 885804 675778 885806
rect 676029 885730 676095 885733
rect 676029 885728 676292 885730
rect 676029 885672 676034 885728
rect 676090 885672 676292 885728
rect 676029 885670 676292 885672
rect 676029 885667 676095 885670
rect 675518 880636 675524 880700
rect 675588 880698 675594 880700
rect 680997 880698 681063 880701
rect 675588 880696 681063 880698
rect 675588 880640 681002 880696
rect 681058 880640 681063 880696
rect 675588 880638 681063 880640
rect 675588 880636 675594 880638
rect 680997 880635 681063 880638
rect 676254 880364 676260 880428
rect 676324 880426 676330 880428
rect 683113 880426 683179 880429
rect 676324 880424 683179 880426
rect 676324 880368 683118 880424
rect 683174 880368 683179 880424
rect 676324 880366 683179 880368
rect 676324 880364 676330 880366
rect 683113 880363 683179 880366
rect 675334 878460 675340 878524
rect 675404 878522 675410 878524
rect 675753 878522 675819 878525
rect 675404 878520 675819 878522
rect 675404 878464 675758 878520
rect 675814 878464 675819 878520
rect 675404 878462 675819 878464
rect 675404 878460 675410 878462
rect 675753 878459 675819 878462
rect 675334 874108 675340 874172
rect 675404 874170 675410 874172
rect 675569 874170 675635 874173
rect 675404 874168 675635 874170
rect 675404 874112 675574 874168
rect 675630 874112 675635 874168
rect 675404 874110 675635 874112
rect 675404 874108 675410 874110
rect 675569 874107 675635 874110
rect 675017 873082 675083 873085
rect 676438 873082 676444 873084
rect 675017 873080 676444 873082
rect 675017 873024 675022 873080
rect 675078 873024 676444 873080
rect 675017 873022 676444 873024
rect 675017 873019 675083 873022
rect 676438 873020 676444 873022
rect 676508 873020 676514 873084
rect 675753 872810 675819 872813
rect 676254 872810 676260 872812
rect 675753 872808 676260 872810
rect 675753 872752 675758 872808
rect 675814 872752 676260 872808
rect 675753 872750 676260 872752
rect 675753 872747 675819 872750
rect 676254 872748 676260 872750
rect 676324 872748 676330 872812
rect 675017 869410 675083 869413
rect 674974 869408 675083 869410
rect 674974 869352 675022 869408
rect 675078 869352 675083 869408
rect 674974 869347 675083 869352
rect 674974 869005 675034 869347
rect 674974 869000 675083 869005
rect 674974 868944 675022 869000
rect 675078 868944 675083 869000
rect 674974 868942 675083 868944
rect 675017 868939 675083 868942
rect 651465 868594 651531 868597
rect 649950 868592 651531 868594
rect 649950 868536 651470 868592
rect 651526 868536 651531 868592
rect 649950 868534 651531 868536
rect 649950 868246 650010 868534
rect 651465 868531 651531 868534
rect 674281 868594 674347 868597
rect 675385 868594 675451 868597
rect 674281 868592 675451 868594
rect 674281 868536 674286 868592
rect 674342 868536 675390 868592
rect 675446 868536 675451 868592
rect 674281 868534 675451 868536
rect 674281 868531 674347 868534
rect 675385 868531 675451 868534
rect 652017 867642 652083 867645
rect 649950 867640 652083 867642
rect 649950 867584 652022 867640
rect 652078 867584 652083 867640
rect 649950 867582 652083 867584
rect 649950 867064 650010 867582
rect 652017 867579 652083 867582
rect 651465 866282 651531 866285
rect 649950 866280 651531 866282
rect 649950 866224 651470 866280
rect 651526 866224 651531 866280
rect 649950 866222 651531 866224
rect 649950 865882 650010 866222
rect 651465 866219 651531 866222
rect 675293 865738 675359 865741
rect 675702 865738 675708 865740
rect 675293 865736 675708 865738
rect 675293 865680 675298 865736
rect 675354 865680 675708 865736
rect 675293 865678 675708 865680
rect 675293 865675 675359 865678
rect 675702 865676 675708 865678
rect 675772 865676 675778 865740
rect 675753 865466 675819 865469
rect 676070 865466 676076 865468
rect 675753 865464 676076 865466
rect 675753 865408 675758 865464
rect 675814 865408 676076 865464
rect 675753 865406 676076 865408
rect 675753 865403 675819 865406
rect 676070 865404 676076 865406
rect 676140 865404 676146 865468
rect 651373 865194 651439 865197
rect 649950 865192 651439 865194
rect 649950 865136 651378 865192
rect 651434 865136 651439 865192
rect 649950 865134 651439 865136
rect 649950 864700 650010 865134
rect 651373 865131 651439 865134
rect 675661 865058 675727 865061
rect 675886 865058 675892 865060
rect 675661 865056 675892 865058
rect 675661 865000 675666 865056
rect 675722 865000 675892 865056
rect 675661 864998 675892 865000
rect 675661 864995 675727 864998
rect 675886 864996 675892 864998
rect 675956 864996 675962 865060
rect 651465 863834 651531 863837
rect 649766 863832 651531 863834
rect 649766 863776 651470 863832
rect 651526 863776 651531 863832
rect 649766 863774 651531 863776
rect 649766 863518 649826 863774
rect 651465 863771 651531 863774
rect 651465 862338 651531 862341
rect 649766 862336 651531 862338
rect 649766 862280 651470 862336
rect 651526 862280 651531 862336
rect 649766 862278 651531 862280
rect 651465 862275 651531 862278
rect 35617 818002 35683 818005
rect 35574 818000 35683 818002
rect 35574 817944 35622 818000
rect 35678 817944 35683 818000
rect 35574 817939 35683 817944
rect 35574 817700 35634 817939
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 35617 816914 35683 816917
rect 35604 816912 35683 816914
rect 35604 816856 35622 816912
rect 35678 816856 35683 816912
rect 35604 816854 35683 816856
rect 35617 816851 35683 816854
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815282 35683 815285
rect 35604 815280 35683 815282
rect 35604 815224 35622 815280
rect 35678 815224 35683 815280
rect 35604 815222 35683 815224
rect 35617 815219 35683 815222
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41321 813650 41387 813653
rect 41308 813648 41387 813650
rect 41308 813592 41326 813648
rect 41382 813592 41387 813648
rect 41308 813590 41387 813592
rect 41321 813587 41387 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 41137 812834 41203 812837
rect 41124 812832 41203 812834
rect 41124 812776 41142 812832
rect 41198 812776 41203 812832
rect 41124 812774 41203 812776
rect 41137 812771 41203 812774
rect 40493 812426 40559 812429
rect 40493 812424 40572 812426
rect 40493 812368 40498 812424
rect 40554 812368 40572 812424
rect 40493 812366 40572 812368
rect 40493 812363 40559 812366
rect 41822 812018 41828 812020
rect 41492 811958 41828 812018
rect 41822 811956 41828 811958
rect 41892 811956 41898 812020
rect 39297 811610 39363 811613
rect 39284 811608 39363 811610
rect 39284 811552 39302 811608
rect 39358 811552 39363 811608
rect 39284 811550 39363 811552
rect 39297 811547 39363 811550
rect 33041 811202 33107 811205
rect 33028 811200 33107 811202
rect 33028 811144 33046 811200
rect 33102 811144 33107 811200
rect 33028 811142 33107 811144
rect 33041 811139 33107 811142
rect 41781 810794 41847 810797
rect 41492 810792 41847 810794
rect 41492 810736 41786 810792
rect 41842 810736 41847 810792
rect 41492 810734 41847 810736
rect 41781 810731 41847 810734
rect 41965 810386 42031 810389
rect 41492 810384 42031 810386
rect 41492 810328 41970 810384
rect 42026 810328 42031 810384
rect 41492 810326 42031 810328
rect 41965 810323 42031 810326
rect 31017 809978 31083 809981
rect 31004 809976 31083 809978
rect 31004 809920 31022 809976
rect 31078 809920 31083 809976
rect 31004 809918 31083 809920
rect 31017 809915 31083 809918
rect 33777 809570 33843 809573
rect 33764 809568 33843 809570
rect 33764 809512 33782 809568
rect 33838 809512 33843 809568
rect 33764 809510 33843 809512
rect 33777 809507 33843 809510
rect 40677 809162 40743 809165
rect 40677 809160 40756 809162
rect 40677 809104 40682 809160
rect 40738 809104 40756 809160
rect 40677 809102 40756 809104
rect 40677 809099 40743 809102
rect 41781 808754 41847 808757
rect 41492 808752 41847 808754
rect 41492 808696 41786 808752
rect 41842 808696 41847 808752
rect 41492 808694 41847 808696
rect 41781 808691 41847 808694
rect 40953 808346 41019 808349
rect 40940 808344 41019 808346
rect 40940 808288 40958 808344
rect 41014 808288 41019 808344
rect 40940 808286 41019 808288
rect 40953 808283 41019 808286
rect 41137 807938 41203 807941
rect 41124 807936 41203 807938
rect 41124 807880 41142 807936
rect 41198 807880 41203 807936
rect 41124 807878 41203 807880
rect 41137 807875 41203 807878
rect 42885 807530 42951 807533
rect 41492 807528 42951 807530
rect 41492 807472 42890 807528
rect 42946 807472 42951 807528
rect 41492 807470 42951 807472
rect 42885 807467 42951 807470
rect 31710 806717 31770 807092
rect 31710 806712 31819 806717
rect 31710 806684 31758 806712
rect 31740 806656 31758 806684
rect 31814 806656 31819 806712
rect 31740 806654 31819 806656
rect 31753 806651 31819 806654
rect 41321 806306 41387 806309
rect 41308 806304 41387 806306
rect 41308 806248 41326 806304
rect 41382 806248 41387 806304
rect 41308 806246 41387 806248
rect 41321 806243 41387 806246
rect 40493 805626 40559 805629
rect 41638 805626 41644 805628
rect 40493 805624 41644 805626
rect 40493 805568 40498 805624
rect 40554 805568 41644 805624
rect 40493 805566 41644 805568
rect 40493 805563 40559 805566
rect 41638 805564 41644 805566
rect 41708 805564 41714 805628
rect 40902 805156 40908 805220
rect 40972 805218 40978 805220
rect 41781 805218 41847 805221
rect 40972 805216 41847 805218
rect 40972 805160 41786 805216
rect 41842 805160 41847 805216
rect 40972 805158 41847 805160
rect 40972 805156 40978 805158
rect 41781 805155 41847 805158
rect 40718 804884 40724 804948
rect 40788 804946 40794 804948
rect 41965 804946 42031 804949
rect 40788 804944 42031 804946
rect 40788 804888 41970 804944
rect 42026 804888 42031 804944
rect 40788 804886 42031 804888
rect 40788 804884 40794 804886
rect 41965 804883 42031 804886
rect 40534 804612 40540 804676
rect 40604 804674 40610 804676
rect 41597 804674 41663 804677
rect 40604 804672 41663 804674
rect 40604 804616 41602 804672
rect 41658 804616 41663 804672
rect 40604 804614 41663 804616
rect 40604 804612 40610 804614
rect 41597 804611 41663 804614
rect 40125 800866 40191 800869
rect 40350 800866 40356 800868
rect 40125 800864 40356 800866
rect 40125 800808 40130 800864
rect 40186 800808 40356 800864
rect 40125 800806 40356 800808
rect 40125 800803 40191 800806
rect 40350 800804 40356 800806
rect 40420 800804 40426 800868
rect 40677 800594 40743 800597
rect 41086 800594 41092 800596
rect 40677 800592 41092 800594
rect 40677 800536 40682 800592
rect 40738 800536 41092 800592
rect 40677 800534 41092 800536
rect 40677 800531 40743 800534
rect 41086 800532 41092 800534
rect 41156 800532 41162 800596
rect 41965 800324 42031 800325
rect 41965 800322 42012 800324
rect 41920 800320 42012 800322
rect 41920 800264 41970 800320
rect 41920 800262 42012 800264
rect 41965 800260 42012 800262
rect 42076 800260 42082 800324
rect 41965 800259 42031 800260
rect 42149 797330 42215 797333
rect 43437 797330 43503 797333
rect 42149 797328 43503 797330
rect 42149 797272 42154 797328
rect 42210 797272 43442 797328
rect 43498 797272 43503 797328
rect 42149 797270 43503 797272
rect 42149 797267 42215 797270
rect 43437 797267 43503 797270
rect 40350 796180 40356 796244
rect 40420 796242 40426 796244
rect 41781 796242 41847 796245
rect 40420 796240 41847 796242
rect 40420 796184 41786 796240
rect 41842 796184 41847 796240
rect 40420 796182 41847 796184
rect 40420 796180 40426 796182
rect 41781 796179 41847 796182
rect 41086 794412 41092 794476
rect 41156 794474 41162 794476
rect 41781 794474 41847 794477
rect 41156 794472 41847 794474
rect 41156 794416 41786 794472
rect 41842 794416 41847 794472
rect 41156 794414 41847 794416
rect 41156 794412 41162 794414
rect 41781 794411 41847 794414
rect 42057 792980 42123 792981
rect 42006 792978 42012 792980
rect 41966 792918 42012 792978
rect 42076 792976 42123 792980
rect 42118 792920 42123 792976
rect 42006 792916 42012 792918
rect 42076 792916 42123 792920
rect 42057 792915 42123 792916
rect 41822 791556 41828 791620
rect 41892 791618 41898 791620
rect 42609 791618 42675 791621
rect 41892 791616 42675 791618
rect 41892 791560 42614 791616
rect 42670 791560 42675 791616
rect 41892 791558 42675 791560
rect 41892 791556 41898 791558
rect 42609 791555 42675 791558
rect 40718 791284 40724 791348
rect 40788 791346 40794 791348
rect 42241 791346 42307 791349
rect 40788 791344 42307 791346
rect 40788 791288 42246 791344
rect 42302 791288 42307 791344
rect 40788 791286 42307 791288
rect 40788 791284 40794 791286
rect 42241 791283 42307 791286
rect 40902 790604 40908 790668
rect 40972 790666 40978 790668
rect 41781 790666 41847 790669
rect 40972 790664 41847 790666
rect 40972 790608 41786 790664
rect 41842 790608 41847 790664
rect 40972 790606 41847 790608
rect 40972 790604 40978 790606
rect 41781 790603 41847 790606
rect 62205 790530 62271 790533
rect 62205 790528 64706 790530
rect 62205 790472 62210 790528
rect 62266 790472 64706 790528
rect 62205 790470 64706 790472
rect 62205 790467 62271 790470
rect 64646 790304 64706 790470
rect 62113 789170 62179 789173
rect 62113 789168 64706 789170
rect 62113 789112 62118 789168
rect 62174 789112 64706 789168
rect 62113 789110 64706 789112
rect 62113 789107 62179 789110
rect 41638 788156 41644 788220
rect 41708 788218 41714 788220
rect 42241 788218 42307 788221
rect 41708 788216 42307 788218
rect 41708 788160 42246 788216
rect 42302 788160 42307 788216
rect 41708 788158 42307 788160
rect 41708 788156 41714 788158
rect 42241 788155 42307 788158
rect 62113 787402 62179 787405
rect 64646 787402 64706 787940
rect 62113 787400 64706 787402
rect 62113 787344 62118 787400
rect 62174 787344 64706 787400
rect 62113 787342 64706 787344
rect 62113 787339 62179 787342
rect 62757 787130 62823 787133
rect 62757 787128 64706 787130
rect 62757 787072 62762 787128
rect 62818 787072 64706 787128
rect 62757 787070 64706 787072
rect 62757 787067 62823 787070
rect 41454 786796 41460 786860
rect 41524 786858 41530 786860
rect 41781 786858 41847 786861
rect 41524 786856 41847 786858
rect 41524 786800 41786 786856
rect 41842 786800 41847 786856
rect 41524 786798 41847 786800
rect 41524 786796 41530 786798
rect 41781 786795 41847 786798
rect 64646 786758 64706 787070
rect 675753 786722 675819 786725
rect 676070 786722 676076 786724
rect 675753 786720 676076 786722
rect 675753 786664 675758 786720
rect 675814 786664 676076 786720
rect 675753 786662 676076 786664
rect 675753 786659 675819 786662
rect 676070 786660 676076 786662
rect 676140 786660 676146 786724
rect 40534 786116 40540 786180
rect 40604 786178 40610 786180
rect 41781 786178 41847 786181
rect 40604 786176 41847 786178
rect 40604 786120 41786 786176
rect 41842 786120 41847 786176
rect 40604 786118 41847 786120
rect 40604 786116 40610 786118
rect 41781 786115 41847 786118
rect 61377 786178 61443 786181
rect 61377 786176 64706 786178
rect 61377 786120 61382 786176
rect 61438 786120 64706 786176
rect 61377 786118 64706 786120
rect 61377 786115 61443 786118
rect 64646 785576 64706 786118
rect 62113 784954 62179 784957
rect 62113 784952 64706 784954
rect 62113 784896 62118 784952
rect 62174 784896 64706 784952
rect 62113 784894 64706 784896
rect 62113 784891 62179 784894
rect 64646 784394 64706 784894
rect 674230 783804 674236 783868
rect 674300 783866 674306 783868
rect 675477 783866 675543 783869
rect 674300 783864 675543 783866
rect 674300 783808 675482 783864
rect 675538 783808 675543 783864
rect 674300 783806 675543 783808
rect 674300 783804 674306 783806
rect 675477 783803 675543 783806
rect 674598 782444 674604 782508
rect 674668 782506 674674 782508
rect 675109 782506 675175 782509
rect 674668 782504 675175 782506
rect 674668 782448 675114 782504
rect 675170 782448 675175 782504
rect 674668 782446 675175 782448
rect 674668 782444 674674 782446
rect 675109 782443 675175 782446
rect 671613 779378 671679 779381
rect 675477 779378 675543 779381
rect 671613 779376 675543 779378
rect 671613 779320 671618 779376
rect 671674 779320 675482 779376
rect 675538 779320 675543 779376
rect 671613 779318 675543 779320
rect 671613 779315 671679 779318
rect 675477 779315 675543 779318
rect 673729 778834 673795 778837
rect 675477 778834 675543 778837
rect 673729 778832 675543 778834
rect 649950 778426 650010 778824
rect 673729 778776 673734 778832
rect 673790 778776 675482 778832
rect 675538 778776 675543 778832
rect 673729 778774 675543 778776
rect 673729 778771 673795 778774
rect 675477 778771 675543 778774
rect 651465 778426 651531 778429
rect 649950 778424 651531 778426
rect 649950 778368 651470 778424
rect 651526 778368 651531 778424
rect 649950 778366 651531 778368
rect 651465 778363 651531 778366
rect 649950 777066 650010 777642
rect 674465 777474 674531 777477
rect 675477 777474 675543 777477
rect 674465 777472 675543 777474
rect 674465 777416 674470 777472
rect 674526 777416 675482 777472
rect 675538 777416 675543 777472
rect 674465 777414 675543 777416
rect 674465 777411 674531 777414
rect 675477 777411 675543 777414
rect 652017 777066 652083 777069
rect 649950 777064 652083 777066
rect 649950 777008 652022 777064
rect 652078 777008 652083 777064
rect 649950 777006 652083 777008
rect 652017 777003 652083 777006
rect 40493 776658 40559 776661
rect 45001 776658 45067 776661
rect 40493 776656 45067 776658
rect 40493 776600 40498 776656
rect 40554 776600 45006 776656
rect 45062 776600 45067 776656
rect 40493 776598 45067 776600
rect 40493 776595 40559 776598
rect 45001 776595 45067 776598
rect 649950 776114 650010 776460
rect 651465 776114 651531 776117
rect 649950 776112 651531 776114
rect 649950 776056 651470 776112
rect 651526 776056 651531 776112
rect 649950 776054 651531 776056
rect 651465 776051 651531 776054
rect 674097 775706 674163 775709
rect 675477 775706 675543 775709
rect 674097 775704 675543 775706
rect 674097 775648 674102 775704
rect 674158 775648 675482 775704
rect 675538 775648 675543 775704
rect 674097 775646 675543 775648
rect 674097 775643 674163 775646
rect 675477 775643 675543 775646
rect 651373 775298 651439 775301
rect 649950 775296 651439 775298
rect 649950 775240 651378 775296
rect 651434 775240 651439 775296
rect 649950 775238 651439 775240
rect 651373 775235 651439 775238
rect 35801 774754 35867 774757
rect 35758 774752 35867 774754
rect 35758 774696 35806 774752
rect 35862 774696 35867 774752
rect 35758 774691 35867 774696
rect 35758 774452 35818 774691
rect 651465 774210 651531 774213
rect 649950 774208 651531 774210
rect 649950 774152 651470 774208
rect 651526 774152 651531 774208
rect 649950 774150 651531 774152
rect 649950 774096 650010 774150
rect 651465 774147 651531 774150
rect 35206 773941 35266 774044
rect 35157 773936 35266 773941
rect 35157 773880 35162 773936
rect 35218 773880 35266 773936
rect 35157 773878 35266 773880
rect 35157 773875 35223 773878
rect 35390 773533 35450 773636
rect 35341 773528 35450 773533
rect 35341 773472 35346 773528
rect 35402 773472 35450 773528
rect 35341 773470 35450 773472
rect 35341 773467 35407 773470
rect 651465 773394 651531 773397
rect 649950 773392 651531 773394
rect 649950 773336 651470 773392
rect 651526 773336 651531 773392
rect 649950 773334 651531 773336
rect 35758 773125 35818 773228
rect 35525 773122 35591 773125
rect 35525 773120 35634 773122
rect 35525 773064 35530 773120
rect 35586 773064 35634 773120
rect 35525 773059 35634 773064
rect 35758 773120 35867 773125
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773062 35867 773064
rect 35801 773059 35867 773062
rect 40493 773122 40559 773125
rect 44909 773122 44975 773125
rect 40493 773120 44975 773122
rect 40493 773064 40498 773120
rect 40554 773064 44914 773120
rect 44970 773064 44975 773120
rect 40493 773062 44975 773064
rect 40493 773059 40559 773062
rect 44909 773059 44975 773062
rect 35574 772820 35634 773059
rect 649950 772914 650010 773334
rect 651465 773331 651531 773334
rect 35574 772309 35634 772412
rect 35574 772304 35683 772309
rect 35574 772248 35622 772304
rect 35678 772248 35683 772304
rect 35574 772246 35683 772248
rect 35617 772243 35683 772246
rect 41321 772306 41387 772309
rect 44265 772306 44331 772309
rect 41321 772304 44331 772306
rect 41321 772248 41326 772304
rect 41382 772248 44270 772304
rect 44326 772248 44331 772304
rect 41321 772246 44331 772248
rect 41321 772243 41387 772246
rect 44265 772243 44331 772246
rect 35758 771901 35818 772004
rect 35758 771896 35867 771901
rect 35758 771840 35806 771896
rect 35862 771840 35867 771896
rect 35758 771838 35867 771840
rect 35801 771835 35867 771838
rect 35758 771493 35818 771596
rect 35758 771488 35867 771493
rect 35758 771432 35806 771488
rect 35862 771432 35867 771488
rect 35758 771430 35867 771432
rect 35801 771427 35867 771430
rect 39573 771490 39639 771493
rect 43069 771490 43135 771493
rect 39573 771488 43135 771490
rect 39573 771432 39578 771488
rect 39634 771432 43074 771488
rect 43130 771432 43135 771488
rect 39573 771430 43135 771432
rect 39573 771427 39639 771430
rect 43069 771427 43135 771430
rect 35574 771085 35634 771188
rect 35574 771080 35683 771085
rect 35574 771024 35622 771080
rect 35678 771024 35683 771080
rect 35574 771022 35683 771024
rect 35617 771019 35683 771022
rect 35758 770677 35818 770780
rect 35758 770672 35867 770677
rect 35758 770616 35806 770672
rect 35862 770616 35867 770672
rect 35758 770614 35867 770616
rect 35801 770611 35867 770614
rect 40033 770674 40099 770677
rect 43253 770674 43319 770677
rect 40033 770672 43319 770674
rect 40033 770616 40038 770672
rect 40094 770616 43258 770672
rect 43314 770616 43319 770672
rect 40033 770614 43319 770616
rect 40033 770611 40099 770614
rect 43253 770611 43319 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35390 769453 35450 769556
rect 35341 769448 35450 769453
rect 35341 769392 35346 769448
rect 35402 769392 35450 769448
rect 35341 769390 35450 769392
rect 35341 769387 35407 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 39757 768634 39823 768637
rect 42701 768634 42767 768637
rect 39757 768632 42767 768634
rect 39757 768576 39762 768632
rect 39818 768576 42706 768632
rect 42762 768576 42767 768632
rect 39757 768574 42767 768576
rect 39757 768571 39823 768574
rect 42701 768571 42767 768574
rect 35574 768229 35634 768332
rect 35574 768224 35683 768229
rect 35574 768168 35622 768224
rect 35678 768168 35683 768224
rect 35574 768166 35683 768168
rect 35617 768163 35683 768166
rect 32998 767821 33058 767924
rect 32998 767816 33107 767821
rect 35801 767818 35867 767821
rect 32998 767760 33046 767816
rect 33102 767760 33107 767816
rect 32998 767758 33107 767760
rect 33041 767755 33107 767758
rect 35758 767816 35867 767818
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35758 767755 35867 767760
rect 35758 767516 35818 767755
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 40309 767002 40375 767005
rect 44541 767002 44607 767005
rect 40309 767000 44607 767002
rect 40309 766944 40314 767000
rect 40370 766944 44546 767000
rect 44602 766944 44607 767000
rect 40309 766942 44607 766944
rect 35157 766939 35223 766942
rect 40309 766939 40375 766942
rect 44541 766939 44607 766942
rect 35801 766594 35867 766597
rect 40726 766596 40786 766700
rect 35758 766592 35867 766594
rect 35758 766536 35806 766592
rect 35862 766536 35867 766592
rect 35758 766531 35867 766536
rect 40718 766532 40724 766596
rect 40788 766532 40794 766596
rect 35758 766292 35818 766531
rect 35758 765781 35818 765884
rect 35758 765776 35867 765781
rect 35758 765720 35806 765776
rect 35862 765720 35867 765776
rect 35758 765718 35867 765720
rect 35801 765715 35867 765718
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40910 764964 40970 765068
rect 40902 764900 40908 764964
rect 40972 764900 40978 764964
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 39297 764554 39363 764557
rect 45093 764554 45159 764557
rect 39297 764552 45159 764554
rect 39297 764496 39302 764552
rect 39358 764496 45098 764552
rect 45154 764496 45159 764552
rect 39297 764494 45159 764496
rect 39297 764491 39363 764494
rect 45093 764491 45159 764494
rect 35758 764149 35818 764252
rect 35758 764144 35867 764149
rect 35758 764088 35806 764144
rect 35862 764088 35867 764144
rect 35758 764086 35867 764088
rect 35801 764083 35867 764086
rect 40401 764146 40467 764149
rect 43621 764146 43687 764149
rect 40401 764144 43687 764146
rect 40401 764088 40406 764144
rect 40462 764088 43626 764144
rect 43682 764088 43687 764144
rect 40401 764086 43687 764088
rect 40401 764083 40467 764086
rect 43621 764083 43687 764086
rect 37046 763741 37106 763844
rect 37046 763738 37155 763741
rect 41689 763738 41755 763741
rect 45277 763738 45343 763741
rect 37046 763736 37236 763738
rect 37046 763680 37094 763736
rect 37150 763680 37236 763736
rect 37046 763678 37236 763680
rect 41689 763736 45343 763738
rect 41689 763680 41694 763736
rect 41750 763680 45282 763736
rect 45338 763680 45343 763736
rect 41689 763678 45343 763680
rect 37046 763675 37155 763678
rect 41689 763675 41755 763678
rect 45277 763675 45343 763678
rect 37046 763436 37106 763675
rect 41689 763330 41755 763333
rect 45553 763330 45619 763333
rect 41689 763328 45619 763330
rect 41689 763272 41694 763328
rect 41750 763272 45558 763328
rect 45614 763272 45619 763328
rect 41689 763270 45619 763272
rect 41689 763267 41755 763270
rect 45553 763267 45619 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 40493 759522 40559 759525
rect 42425 759522 42491 759525
rect 40493 759520 42491 759522
rect 40493 759464 40498 759520
rect 40554 759464 42430 759520
rect 42486 759464 42491 759520
rect 40493 759462 42491 759464
rect 40493 759459 40559 759462
rect 42425 759459 42491 759462
rect 36537 759114 36603 759117
rect 42006 759114 42012 759116
rect 36537 759112 42012 759114
rect 36537 759056 36542 759112
rect 36598 759056 42012 759112
rect 36537 759054 42012 759056
rect 36537 759051 36603 759054
rect 42006 759052 42012 759054
rect 42076 759052 42082 759116
rect 42149 758980 42215 758981
rect 42149 758976 42196 758980
rect 42260 758978 42266 758980
rect 42149 758920 42154 758976
rect 42149 758916 42196 758920
rect 42260 758918 42306 758978
rect 42260 758916 42266 758918
rect 42149 758915 42215 758916
rect 40677 757754 40743 757757
rect 41638 757754 41644 757756
rect 40677 757752 41644 757754
rect 40677 757696 40682 757752
rect 40738 757696 41644 757752
rect 40677 757694 41644 757696
rect 40677 757691 40743 757694
rect 41638 757692 41644 757694
rect 41708 757692 41714 757756
rect 39941 757482 40007 757485
rect 43253 757482 43319 757485
rect 39941 757480 43319 757482
rect 39941 757424 39946 757480
rect 40002 757424 43258 757480
rect 43314 757424 43319 757480
rect 39941 757422 43319 757424
rect 39941 757419 40007 757422
rect 43253 757419 43319 757422
rect 41781 757076 41847 757077
rect 41781 757074 41828 757076
rect 41736 757072 41828 757074
rect 41736 757016 41786 757072
rect 41736 757014 41828 757016
rect 41781 757012 41828 757014
rect 41892 757012 41898 757076
rect 41781 757011 41847 757012
rect 41873 755444 41939 755445
rect 41822 755442 41828 755444
rect 41782 755382 41828 755442
rect 41892 755440 41939 755444
rect 41934 755384 41939 755440
rect 41822 755380 41828 755382
rect 41892 755380 41939 755384
rect 41873 755379 41939 755380
rect 42149 754900 42215 754901
rect 40902 754836 40908 754900
rect 40972 754898 40978 754900
rect 41822 754898 41828 754900
rect 40972 754838 41828 754898
rect 40972 754836 40978 754838
rect 41822 754836 41828 754838
rect 41892 754836 41898 754900
rect 42149 754896 42196 754900
rect 42260 754898 42266 754900
rect 42149 754840 42154 754896
rect 42149 754836 42196 754840
rect 42260 754838 42306 754898
rect 42260 754836 42266 754838
rect 42149 754835 42215 754836
rect 42057 754082 42123 754085
rect 44725 754082 44791 754085
rect 42057 754080 44791 754082
rect 42057 754024 42062 754080
rect 42118 754024 44730 754080
rect 44786 754024 44791 754080
rect 42057 754022 44791 754024
rect 42057 754019 42123 754022
rect 44725 754019 44791 754022
rect 42057 752994 42123 752997
rect 43437 752994 43503 752997
rect 42057 752992 43503 752994
rect 42057 752936 42062 752992
rect 42118 752936 43442 752992
rect 43498 752936 43503 752992
rect 42057 752934 43503 752936
rect 42057 752931 42123 752934
rect 43437 752931 43503 752934
rect 42057 751770 42123 751773
rect 45093 751770 45159 751773
rect 42057 751768 45159 751770
rect 42057 751712 42062 751768
rect 42118 751712 45098 751768
rect 45154 751712 45159 751768
rect 42057 751710 45159 751712
rect 42057 751707 42123 751710
rect 45093 751707 45159 751710
rect 41781 750412 41847 750413
rect 41781 750408 41828 750412
rect 41892 750410 41898 750412
rect 41781 750352 41786 750408
rect 41781 750348 41828 750352
rect 41892 750350 41938 750410
rect 41892 750348 41898 750350
rect 41781 750347 41847 750348
rect 40534 749532 40540 749596
rect 40604 749594 40610 749596
rect 42333 749594 42399 749597
rect 40604 749592 42399 749594
rect 40604 749536 42338 749592
rect 42394 749536 42399 749592
rect 40604 749534 42399 749536
rect 40604 749532 40610 749534
rect 42333 749531 42399 749534
rect 62757 747690 62823 747693
rect 62757 747688 64706 747690
rect 62757 747632 62762 747688
rect 62818 747632 64706 747688
rect 62757 747630 64706 747632
rect 62757 747627 62823 747630
rect 64646 747082 64706 747630
rect 40718 746676 40724 746740
rect 40788 746738 40794 746740
rect 41781 746738 41847 746741
rect 40788 746736 41847 746738
rect 40788 746680 41786 746736
rect 41842 746680 41847 746736
rect 40788 746678 41847 746680
rect 40788 746676 40794 746678
rect 41781 746675 41847 746678
rect 62113 746194 62179 746197
rect 62113 746192 64706 746194
rect 62113 746136 62118 746192
rect 62174 746136 64706 746192
rect 62113 746134 64706 746136
rect 62113 746131 62179 746134
rect 64646 745900 64706 746134
rect 41638 745044 41644 745108
rect 41708 745106 41714 745108
rect 42517 745106 42583 745109
rect 41708 745104 42583 745106
rect 41708 745048 42522 745104
rect 42578 745048 42583 745104
rect 41708 745046 42583 745048
rect 41708 745044 41714 745046
rect 42517 745043 42583 745046
rect 42057 744836 42123 744837
rect 42006 744834 42012 744836
rect 41966 744774 42012 744834
rect 42076 744832 42123 744836
rect 42118 744776 42123 744832
rect 42006 744772 42012 744774
rect 42076 744772 42123 744776
rect 42057 744771 42123 744772
rect 62113 744154 62179 744157
rect 64646 744154 64706 744718
rect 62113 744152 64706 744154
rect 62113 744096 62118 744152
rect 62174 744096 64706 744152
rect 62113 744094 64706 744096
rect 62113 744091 62179 744094
rect 41454 743684 41460 743748
rect 41524 743746 41530 743748
rect 41781 743746 41847 743749
rect 41524 743744 41847 743746
rect 41524 743688 41786 743744
rect 41842 743688 41847 743744
rect 41524 743686 41847 743688
rect 41524 743684 41530 743686
rect 41781 743683 41847 743686
rect 62113 743746 62179 743749
rect 62113 743744 64706 743746
rect 62113 743688 62118 743744
rect 62174 743688 64706 743744
rect 62113 743686 64706 743688
rect 62113 743683 62179 743686
rect 64646 743536 64706 743686
rect 62113 742386 62179 742389
rect 62113 742384 64706 742386
rect 62113 742328 62118 742384
rect 62174 742328 64706 742384
rect 62113 742326 64706 742328
rect 62113 742323 62179 742326
rect 62389 741842 62455 741845
rect 62389 741840 64706 741842
rect 62389 741784 62394 741840
rect 62450 741784 64706 741840
rect 62389 741782 64706 741784
rect 62389 741779 62455 741782
rect 64646 741172 64706 741782
rect 675753 739802 675819 739805
rect 676806 739802 676812 739804
rect 675753 739800 676812 739802
rect 675753 739744 675758 739800
rect 675814 739744 676812 739800
rect 675753 739742 676812 739744
rect 675753 739739 675819 739742
rect 676806 739740 676812 739742
rect 676876 739740 676882 739804
rect 674414 738108 674420 738172
rect 674484 738170 674490 738172
rect 675293 738170 675359 738173
rect 674484 738168 675359 738170
rect 674484 738112 675298 738168
rect 675354 738112 675359 738168
rect 674484 738110 675359 738112
rect 674484 738108 674490 738110
rect 675293 738107 675359 738110
rect 673821 735722 673887 735725
rect 675477 735722 675543 735725
rect 673821 735720 675543 735722
rect 673821 735664 673826 735720
rect 673882 735664 675482 735720
rect 675538 735664 675543 735720
rect 673821 735662 675543 735664
rect 673821 735659 673887 735662
rect 675477 735659 675543 735662
rect 674097 735042 674163 735045
rect 675477 735042 675543 735045
rect 674097 735040 675543 735042
rect 674097 734984 674102 735040
rect 674158 734984 675482 735040
rect 675538 734984 675543 735040
rect 674097 734982 675543 734984
rect 674097 734979 674163 734982
rect 675477 734979 675543 734982
rect 649950 734226 650010 734402
rect 651465 734226 651531 734229
rect 649950 734224 651531 734226
rect 649950 734168 651470 734224
rect 651526 734168 651531 734224
rect 649950 734166 651531 734168
rect 651465 734163 651531 734166
rect 669037 733818 669103 733821
rect 675569 733818 675635 733821
rect 669037 733816 675635 733818
rect 669037 733760 669042 733816
rect 669098 733760 675574 733816
rect 675630 733760 675635 733816
rect 669037 733758 675635 733760
rect 669037 733755 669103 733758
rect 675569 733755 675635 733758
rect 649950 733002 650010 733220
rect 651465 733002 651531 733005
rect 649950 733000 651531 733002
rect 649950 732944 651470 733000
rect 651526 732944 651531 733000
rect 649950 732942 651531 732944
rect 651465 732939 651531 732942
rect 39573 732322 39639 732325
rect 43069 732322 43135 732325
rect 39573 732320 43135 732322
rect 39573 732264 39578 732320
rect 39634 732264 43074 732320
rect 43130 732264 43135 732320
rect 39573 732262 43135 732264
rect 39573 732259 39639 732262
rect 43069 732259 43135 732262
rect 39941 732050 40007 732053
rect 44909 732050 44975 732053
rect 39941 732048 44975 732050
rect 39941 731992 39946 732048
rect 40002 731992 44914 732048
rect 44970 731992 44975 732048
rect 39941 731990 44975 731992
rect 39941 731987 40007 731990
rect 44909 731987 44975 731990
rect 649950 731778 650010 732038
rect 651465 731778 651531 731781
rect 649950 731776 651531 731778
rect 649950 731720 651470 731776
rect 651526 731720 651531 731776
rect 649950 731718 651531 731720
rect 651465 731715 651531 731718
rect 40401 731642 40467 731645
rect 44541 731642 44607 731645
rect 40401 731640 44607 731642
rect 40401 731584 40406 731640
rect 40462 731584 44546 731640
rect 44602 731584 44607 731640
rect 40401 731582 44607 731584
rect 40401 731579 40467 731582
rect 44541 731579 44607 731582
rect 35801 731370 35867 731373
rect 35788 731368 35867 731370
rect 35788 731312 35806 731368
rect 35862 731312 35867 731368
rect 35788 731310 35867 731312
rect 35801 731307 35867 731310
rect 651465 731098 651531 731101
rect 649950 731096 651531 731098
rect 649950 731040 651470 731096
rect 651526 731040 651531 731096
rect 649950 731038 651531 731040
rect 35617 730962 35683 730965
rect 35604 730960 35683 730962
rect 35604 730904 35622 730960
rect 35678 730904 35683 730960
rect 35604 730902 35683 730904
rect 35617 730899 35683 730902
rect 649950 730856 650010 731038
rect 651465 731035 651531 731038
rect 35433 730554 35499 730557
rect 35420 730552 35499 730554
rect 35420 730496 35438 730552
rect 35494 730496 35499 730552
rect 35420 730494 35499 730496
rect 35433 730491 35499 730494
rect 41689 730282 41755 730285
rect 46197 730282 46263 730285
rect 41689 730280 46263 730282
rect 41689 730224 41694 730280
rect 41750 730224 46202 730280
rect 46258 730224 46263 730280
rect 41689 730222 46263 730224
rect 41689 730219 41755 730222
rect 46197 730219 46263 730222
rect 35801 730146 35867 730149
rect 35788 730144 35867 730146
rect 35788 730088 35806 730144
rect 35862 730088 35867 730144
rect 35788 730086 35867 730088
rect 35801 730083 35867 730086
rect 651465 729874 651531 729877
rect 649950 729872 651531 729874
rect 649950 729816 651470 729872
rect 651526 729816 651531 729872
rect 649950 729814 651531 729816
rect 35249 729738 35315 729741
rect 35236 729736 35315 729738
rect 35236 729680 35254 729736
rect 35310 729680 35315 729736
rect 35236 729678 35315 729680
rect 35249 729675 35315 729678
rect 649950 729674 650010 729814
rect 651465 729811 651531 729814
rect 35617 729330 35683 729333
rect 35604 729328 35683 729330
rect 35604 729272 35622 729328
rect 35678 729272 35683 729328
rect 35604 729270 35683 729272
rect 35617 729267 35683 729270
rect 35801 728922 35867 728925
rect 35788 728920 35867 728922
rect 35788 728864 35806 728920
rect 35862 728864 35867 728920
rect 35788 728862 35867 728864
rect 35801 728859 35867 728862
rect 41689 728650 41755 728653
rect 45185 728650 45251 728653
rect 41689 728648 45251 728650
rect 41689 728592 41694 728648
rect 41750 728592 45190 728648
rect 45246 728592 45251 728648
rect 41689 728590 45251 728592
rect 41689 728587 41755 728590
rect 45185 728587 45251 728590
rect 35617 728514 35683 728517
rect 651465 728514 651531 728517
rect 35604 728512 35683 728514
rect 35604 728456 35622 728512
rect 35678 728456 35683 728512
rect 35604 728454 35683 728456
rect 649950 728512 651531 728514
rect 649950 728456 651470 728512
rect 651526 728456 651531 728512
rect 649950 728454 651531 728456
rect 35617 728451 35683 728454
rect 651465 728451 651531 728454
rect 35801 728106 35867 728109
rect 35788 728104 35867 728106
rect 35788 728048 35806 728104
rect 35862 728048 35867 728104
rect 35788 728046 35867 728048
rect 35801 728043 35867 728046
rect 674281 728106 674347 728109
rect 675845 728106 675911 728109
rect 674281 728104 675911 728106
rect 674281 728048 674286 728104
rect 674342 728048 675850 728104
rect 675906 728048 675911 728104
rect 674281 728046 675911 728048
rect 674281 728043 674347 728046
rect 675845 728043 675911 728046
rect 674649 727834 674715 727837
rect 676029 727834 676095 727837
rect 674649 727832 676095 727834
rect 674649 727776 674654 727832
rect 674710 727776 676034 727832
rect 676090 727776 676095 727832
rect 674649 727774 676095 727776
rect 674649 727771 674715 727774
rect 676029 727771 676095 727774
rect 35801 727698 35867 727701
rect 35788 727696 35867 727698
rect 35788 727640 35806 727696
rect 35862 727640 35867 727696
rect 35788 727638 35867 727640
rect 35801 727635 35867 727638
rect 35801 727290 35867 727293
rect 35788 727288 35867 727290
rect 35788 727232 35806 727288
rect 35862 727232 35867 727288
rect 35788 727230 35867 727232
rect 35801 727227 35867 727230
rect 673913 727290 673979 727293
rect 674465 727290 674531 727293
rect 673913 727288 674531 727290
rect 673913 727232 673918 727288
rect 673974 727232 674470 727288
rect 674526 727232 674531 727288
rect 673913 727230 674531 727232
rect 673913 727227 673979 727230
rect 674465 727227 674531 727230
rect 41689 727018 41755 727021
rect 44265 727018 44331 727021
rect 41689 727016 44331 727018
rect 41689 726960 41694 727016
rect 41750 726960 44270 727016
rect 44326 726960 44331 727016
rect 41689 726958 44331 726960
rect 41689 726955 41755 726958
rect 44265 726955 44331 726958
rect 41137 726882 41203 726885
rect 41124 726880 41203 726882
rect 41124 726824 41142 726880
rect 41198 726824 41203 726880
rect 41124 726822 41203 726824
rect 41137 726819 41203 726822
rect 676070 726820 676076 726884
rect 676140 726882 676146 726884
rect 680997 726882 681063 726885
rect 676140 726880 681063 726882
rect 676140 726824 681002 726880
rect 681058 726824 681063 726880
rect 676140 726822 681063 726824
rect 676140 726820 676146 726822
rect 680997 726819 681063 726822
rect 41278 726239 41338 726444
rect 674230 726412 674236 726476
rect 674300 726474 674306 726476
rect 683113 726474 683179 726477
rect 674300 726472 683179 726474
rect 674300 726416 683118 726472
rect 683174 726416 683179 726472
rect 674300 726414 683179 726416
rect 674300 726412 674306 726414
rect 683113 726411 683179 726414
rect 39297 726236 39363 726239
rect 39254 726234 39363 726236
rect 39254 726178 39302 726234
rect 39358 726178 39363 726234
rect 39254 726173 39363 726178
rect 41278 726234 41387 726239
rect 41278 726178 41326 726234
rect 41382 726178 41387 726234
rect 41278 726176 41387 726178
rect 41321 726173 41387 726176
rect 39254 726036 39314 726173
rect 41781 725796 41847 725797
rect 41781 725794 41828 725796
rect 41736 725792 41828 725794
rect 41736 725736 41786 725792
rect 41736 725734 41828 725736
rect 41781 725732 41828 725734
rect 41892 725732 41898 725796
rect 41781 725731 41847 725732
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 41137 725250 41203 725253
rect 41124 725248 41203 725250
rect 41124 725192 41142 725248
rect 41198 725192 41203 725248
rect 41124 725190 41203 725192
rect 41137 725187 41203 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 31661 724434 31727 724437
rect 31661 724432 31740 724434
rect 31661 724376 31666 724432
rect 31722 724376 31740 724432
rect 31661 724374 31740 724376
rect 31661 724371 31727 724374
rect 33041 724026 33107 724029
rect 33028 724024 33107 724026
rect 33028 723968 33046 724024
rect 33102 723968 33107 724024
rect 33028 723966 33107 723968
rect 33041 723963 33107 723966
rect 43437 723618 43503 723621
rect 41492 723616 43503 723618
rect 41492 723560 43442 723616
rect 43498 723560 43503 723616
rect 41492 723558 43503 723560
rect 43437 723555 43503 723558
rect 33777 723210 33843 723213
rect 33764 723208 33843 723210
rect 33764 723152 33782 723208
rect 33838 723152 33843 723208
rect 33764 723150 33843 723152
rect 33777 723147 33843 723150
rect 44449 722802 44515 722805
rect 41492 722800 44515 722802
rect 41492 722744 44454 722800
rect 44510 722744 44515 722800
rect 41492 722742 44515 722744
rect 44449 722739 44515 722742
rect 41965 722394 42031 722397
rect 41492 722392 42031 722394
rect 41492 722336 41970 722392
rect 42026 722336 42031 722392
rect 41492 722334 42031 722336
rect 41965 722331 42031 722334
rect 674833 722260 674899 722261
rect 674782 722258 674788 722260
rect 674742 722198 674788 722258
rect 674852 722256 674899 722260
rect 674894 722200 674899 722256
rect 674782 722196 674788 722198
rect 674852 722196 674899 722200
rect 674833 722195 674899 722196
rect 41781 721986 41847 721989
rect 41492 721984 41847 721986
rect 41492 721928 41786 721984
rect 41842 721928 41847 721984
rect 41492 721926 41847 721928
rect 41781 721923 41847 721926
rect 674649 721986 674715 721989
rect 674649 721984 675034 721986
rect 674649 721928 674654 721984
rect 674710 721928 675034 721984
rect 674649 721926 675034 721928
rect 674649 721923 674715 721926
rect 674974 721714 675034 721926
rect 674974 721654 675218 721714
rect 44633 721578 44699 721581
rect 41492 721576 44699 721578
rect 41492 721520 44638 721576
rect 44694 721520 44699 721576
rect 41492 721518 44699 721520
rect 675158 721578 675218 721654
rect 676070 721578 676076 721580
rect 675158 721518 676076 721578
rect 44633 721515 44699 721518
rect 676070 721516 676076 721518
rect 676140 721516 676146 721580
rect 47209 721170 47275 721173
rect 41492 721168 47275 721170
rect 41492 721112 47214 721168
rect 47270 721112 47275 721168
rect 41492 721110 47275 721112
rect 47209 721107 47275 721110
rect 41278 720357 41338 720732
rect 41278 720352 41387 720357
rect 41278 720324 41326 720352
rect 41308 720296 41326 720324
rect 41382 720296 41387 720352
rect 41308 720294 41387 720296
rect 41321 720291 41387 720294
rect 47025 719946 47091 719949
rect 41492 719944 47091 719946
rect 41492 719888 47030 719944
rect 47086 719888 47091 719944
rect 41492 719886 47091 719888
rect 47025 719883 47091 719886
rect 41137 719266 41203 719269
rect 42609 719266 42675 719269
rect 41137 719264 42675 719266
rect 41137 719208 41142 719264
rect 41198 719208 42614 719264
rect 42670 719208 42675 719264
rect 41137 719206 42675 719208
rect 41137 719203 41203 719206
rect 42609 719203 42675 719206
rect 41505 718994 41571 718997
rect 42609 718994 42675 718997
rect 41505 718992 42675 718994
rect 41505 718936 41510 718992
rect 41566 718936 42614 718992
rect 42670 718936 42675 718992
rect 41505 718934 42675 718936
rect 41505 718931 41571 718934
rect 42609 718931 42675 718934
rect 40718 718524 40724 718588
rect 40788 718586 40794 718588
rect 41781 718586 41847 718589
rect 40788 718584 41847 718586
rect 40788 718528 41786 718584
rect 41842 718528 41847 718584
rect 40788 718526 41847 718528
rect 40788 718524 40794 718526
rect 41781 718523 41847 718526
rect 31661 718314 31727 718317
rect 41638 718314 41644 718316
rect 31661 718312 41644 718314
rect 31661 718256 31666 718312
rect 31722 718256 41644 718312
rect 31661 718254 41644 718256
rect 31661 718251 31727 718254
rect 41638 718252 41644 718254
rect 41708 718252 41714 718316
rect 40534 717980 40540 718044
rect 40604 718042 40610 718044
rect 41965 718042 42031 718045
rect 40604 718040 42031 718042
rect 40604 717984 41970 718040
rect 42026 717984 42031 718040
rect 40604 717982 42031 717984
rect 40604 717980 40610 717982
rect 41965 717979 42031 717982
rect 674005 716546 674071 716549
rect 674005 716544 676292 716546
rect 674005 716488 674010 716544
rect 674066 716488 676292 716544
rect 674005 716486 676292 716488
rect 674005 716483 674071 716486
rect 39297 716138 39363 716141
rect 41822 716138 41828 716140
rect 39297 716136 41828 716138
rect 39297 716080 39302 716136
rect 39358 716080 41828 716136
rect 39297 716078 41828 716080
rect 39297 716075 39363 716078
rect 41822 716076 41828 716078
rect 41892 716076 41898 716140
rect 674005 716138 674071 716141
rect 674005 716136 676292 716138
rect 674005 716080 674010 716136
rect 674066 716080 676292 716136
rect 674005 716078 676292 716080
rect 674005 716075 674071 716078
rect 673269 715730 673335 715733
rect 673269 715728 676292 715730
rect 673269 715672 673274 715728
rect 673330 715672 676292 715728
rect 673269 715670 676292 715672
rect 673269 715667 673335 715670
rect 39849 715594 39915 715597
rect 42425 715594 42491 715597
rect 39849 715592 42491 715594
rect 39849 715536 39854 715592
rect 39910 715536 42430 715592
rect 42486 715536 42491 715592
rect 39849 715534 42491 715536
rect 39849 715531 39915 715534
rect 42425 715531 42491 715534
rect 672533 715322 672599 715325
rect 672533 715320 676292 715322
rect 672533 715264 672538 715320
rect 672594 715264 676292 715320
rect 672533 715262 676292 715264
rect 672533 715259 672599 715262
rect 671797 714914 671863 714917
rect 671797 714912 676292 714914
rect 671797 714856 671802 714912
rect 671858 714856 676292 714912
rect 671797 714854 676292 714856
rect 671797 714851 671863 714854
rect 37733 714506 37799 714509
rect 42057 714506 42123 714509
rect 37733 714504 42123 714506
rect 37733 714448 37738 714504
rect 37794 714448 42062 714504
rect 42118 714448 42123 714504
rect 37733 714446 42123 714448
rect 37733 714443 37799 714446
rect 42057 714443 42123 714446
rect 673085 714506 673151 714509
rect 673085 714504 676292 714506
rect 673085 714448 673090 714504
rect 673146 714448 676292 714504
rect 673085 714446 676292 714448
rect 673085 714443 673151 714446
rect 41229 714236 41295 714237
rect 41229 714234 41276 714236
rect 41184 714232 41276 714234
rect 41184 714176 41234 714232
rect 41184 714174 41276 714176
rect 41229 714172 41276 714174
rect 41340 714172 41346 714236
rect 41229 714171 41295 714172
rect 673269 714098 673335 714101
rect 673269 714096 676292 714098
rect 673269 714040 673274 714096
rect 673330 714040 676292 714096
rect 673269 714038 676292 714040
rect 673269 714035 673335 714038
rect 674005 713690 674071 713693
rect 674005 713688 676292 713690
rect 674005 713632 674010 713688
rect 674066 713632 676292 713688
rect 674005 713630 676292 713632
rect 674005 713627 674071 713630
rect 674005 713282 674071 713285
rect 674005 713280 676292 713282
rect 674005 713224 674010 713280
rect 674066 713224 676292 713280
rect 674005 713222 676292 713224
rect 674005 713219 674071 713222
rect 673453 713010 673519 713013
rect 674741 713010 674807 713013
rect 673453 713008 674807 713010
rect 673453 712952 673458 713008
rect 673514 712952 674746 713008
rect 674802 712952 674807 713008
rect 673453 712950 674807 712952
rect 673453 712947 673519 712950
rect 674741 712947 674807 712950
rect 674925 712874 674991 712877
rect 674925 712872 676292 712874
rect 674925 712816 674930 712872
rect 674986 712816 676292 712872
rect 674925 712814 676292 712816
rect 674925 712811 674991 712814
rect 673545 712738 673611 712741
rect 674373 712738 674439 712741
rect 673545 712736 674439 712738
rect 673545 712680 673550 712736
rect 673606 712680 674378 712736
rect 674434 712680 674439 712736
rect 673545 712678 674439 712680
rect 673545 712675 673611 712678
rect 674373 712675 674439 712678
rect 674005 712466 674071 712469
rect 674005 712464 676292 712466
rect 674005 712408 674010 712464
rect 674066 712408 676292 712464
rect 674005 712406 676292 712408
rect 674005 712403 674071 712406
rect 41270 712132 41276 712196
rect 41340 712194 41346 712196
rect 41781 712194 41847 712197
rect 41340 712192 41847 712194
rect 41340 712136 41786 712192
rect 41842 712136 41847 712192
rect 41340 712134 41847 712136
rect 41340 712132 41346 712134
rect 41781 712131 41847 712134
rect 672165 712194 672231 712197
rect 674925 712194 674991 712197
rect 672165 712192 674991 712194
rect 672165 712136 672170 712192
rect 672226 712136 674930 712192
rect 674986 712136 674991 712192
rect 672165 712134 674991 712136
rect 672165 712131 672231 712134
rect 674925 712131 674991 712134
rect 680997 712058 681063 712061
rect 680997 712056 681076 712058
rect 680997 712000 681002 712056
rect 681058 712000 681076 712056
rect 680997 711998 681076 712000
rect 680997 711995 681063 711998
rect 683297 711650 683363 711653
rect 683284 711648 683363 711650
rect 683284 711592 683302 711648
rect 683358 711592 683363 711648
rect 683284 711590 683363 711592
rect 683297 711587 683363 711590
rect 674005 711242 674071 711245
rect 674005 711240 676292 711242
rect 674005 711184 674010 711240
rect 674066 711184 676292 711240
rect 674005 711182 676292 711184
rect 674005 711179 674071 711182
rect 42149 710834 42215 710837
rect 43621 710834 43687 710837
rect 42149 710832 43687 710834
rect 42149 710776 42154 710832
rect 42210 710776 43626 710832
rect 43682 710776 43687 710832
rect 42149 710774 43687 710776
rect 42149 710771 42215 710774
rect 43621 710771 43687 710774
rect 675385 710834 675451 710837
rect 675385 710832 676292 710834
rect 675385 710776 675390 710832
rect 675446 710776 676292 710832
rect 675385 710774 676292 710776
rect 675385 710771 675451 710774
rect 674005 710426 674071 710429
rect 674005 710424 676292 710426
rect 674005 710368 674010 710424
rect 674066 710368 676292 710424
rect 674005 710366 676292 710368
rect 674005 710363 674071 710366
rect 674005 710018 674071 710021
rect 674005 710016 676292 710018
rect 674005 709960 674010 710016
rect 674066 709960 676292 710016
rect 674005 709958 676292 709960
rect 674005 709955 674071 709958
rect 674005 709610 674071 709613
rect 674005 709608 676292 709610
rect 674005 709552 674010 709608
rect 674066 709552 676292 709608
rect 674005 709550 676292 709552
rect 674005 709547 674071 709550
rect 672901 709202 672967 709205
rect 672901 709200 676292 709202
rect 672901 709144 672906 709200
rect 672962 709144 676292 709200
rect 672901 709142 676292 709144
rect 672901 709139 672967 709142
rect 683113 708794 683179 708797
rect 683100 708792 683179 708794
rect 683100 708736 683118 708792
rect 683174 708736 683179 708792
rect 683100 708734 683179 708736
rect 683113 708731 683179 708734
rect 42057 708522 42123 708525
rect 44449 708522 44515 708525
rect 42057 708520 44515 708522
rect 42057 708464 42062 708520
rect 42118 708464 44454 708520
rect 44510 708464 44515 708520
rect 42057 708462 44515 708464
rect 42057 708459 42123 708462
rect 44449 708459 44515 708462
rect 683481 708386 683547 708389
rect 683468 708384 683547 708386
rect 683468 708328 683486 708384
rect 683542 708328 683547 708384
rect 683468 708326 683547 708328
rect 683481 708323 683547 708326
rect 674005 707978 674071 707981
rect 674005 707976 676292 707978
rect 674005 707920 674010 707976
rect 674066 707920 676292 707976
rect 674005 707918 676292 707920
rect 674005 707915 674071 707918
rect 42057 707706 42123 707709
rect 43621 707706 43687 707709
rect 42057 707704 43687 707706
rect 42057 707648 42062 707704
rect 42118 707648 43626 707704
rect 43682 707648 43687 707704
rect 42057 707646 43687 707648
rect 42057 707643 42123 707646
rect 43621 707643 43687 707646
rect 674598 707508 674604 707572
rect 674668 707570 674674 707572
rect 674668 707510 676292 707570
rect 674668 707508 674674 707510
rect 40718 707372 40724 707436
rect 40788 707434 40794 707436
rect 41781 707434 41847 707437
rect 40788 707432 41847 707434
rect 40788 707376 41786 707432
rect 41842 707376 41847 707432
rect 40788 707374 41847 707376
rect 40788 707372 40794 707374
rect 41781 707371 41847 707374
rect 674741 707162 674807 707165
rect 674741 707160 676292 707162
rect 674741 707104 674746 707160
rect 674802 707104 676292 707160
rect 674741 707102 676292 707104
rect 674741 707099 674807 707102
rect 674373 706754 674439 706757
rect 674373 706752 676292 706754
rect 674373 706696 674378 706752
rect 674434 706696 676292 706752
rect 674373 706694 676292 706696
rect 674373 706691 674439 706694
rect 674598 706284 674604 706348
rect 674668 706346 674674 706348
rect 674668 706286 676292 706346
rect 674668 706284 674674 706286
rect 40534 706148 40540 706212
rect 40604 706210 40610 706212
rect 42241 706210 42307 706213
rect 40604 706208 42307 706210
rect 40604 706152 42246 706208
rect 42302 706152 42307 706208
rect 40604 706150 42307 706152
rect 40604 706148 40610 706150
rect 42241 706147 42307 706150
rect 678470 705530 678530 705908
rect 683113 705530 683179 705533
rect 678470 705528 683179 705530
rect 678470 705500 683118 705528
rect 678500 705472 683118 705500
rect 683174 705472 683179 705528
rect 678500 705470 683179 705472
rect 683113 705467 683179 705470
rect 674005 705394 674071 705397
rect 675845 705394 675911 705397
rect 674005 705392 675911 705394
rect 674005 705336 674010 705392
rect 674066 705336 675850 705392
rect 675906 705336 675911 705392
rect 674005 705334 675911 705336
rect 674005 705331 674071 705334
rect 675845 705331 675911 705334
rect 674005 705122 674071 705125
rect 674005 705120 676292 705122
rect 674005 705064 674010 705120
rect 674066 705064 676292 705120
rect 674005 705062 676292 705064
rect 674005 705059 674071 705062
rect 62113 704442 62179 704445
rect 62113 704440 64706 704442
rect 62113 704384 62118 704440
rect 62174 704384 64706 704440
rect 62113 704382 64706 704384
rect 62113 704379 62179 704382
rect 64646 703860 64706 704382
rect 42057 703490 42123 703493
rect 43437 703490 43503 703493
rect 42057 703488 43503 703490
rect 42057 703432 42062 703488
rect 42118 703432 43442 703488
rect 43498 703432 43503 703488
rect 42057 703430 43503 703432
rect 42057 703427 42123 703430
rect 43437 703427 43503 703430
rect 62113 703354 62179 703357
rect 62113 703352 64706 703354
rect 62113 703296 62118 703352
rect 62174 703296 64706 703352
rect 62113 703294 64706 703296
rect 62113 703291 62179 703294
rect 64646 702678 64706 703294
rect 41822 702068 41828 702132
rect 41892 702130 41898 702132
rect 42701 702130 42767 702133
rect 41892 702128 42767 702130
rect 41892 702072 42706 702128
rect 42762 702072 42767 702128
rect 41892 702070 42767 702072
rect 41892 702068 41898 702070
rect 42701 702067 42767 702070
rect 41638 701796 41644 701860
rect 41708 701858 41714 701860
rect 42333 701858 42399 701861
rect 41708 701856 42399 701858
rect 41708 701800 42338 701856
rect 42394 701800 42399 701856
rect 41708 701798 42399 701800
rect 41708 701796 41714 701798
rect 42333 701795 42399 701798
rect 62205 701314 62271 701317
rect 64646 701314 64706 701496
rect 62205 701312 64706 701314
rect 62205 701256 62210 701312
rect 62266 701256 64706 701312
rect 62205 701254 64706 701256
rect 62205 701251 62271 701254
rect 673545 701042 673611 701045
rect 675109 701042 675175 701045
rect 673545 701040 675175 701042
rect 673545 700984 673550 701040
rect 673606 700984 675114 701040
rect 675170 700984 675175 701040
rect 673545 700982 675175 700984
rect 673545 700979 673611 700982
rect 675109 700979 675175 700982
rect 62757 700906 62823 700909
rect 62757 700904 64706 700906
rect 62757 700848 62762 700904
rect 62818 700848 64706 700904
rect 62757 700846 64706 700848
rect 62757 700843 62823 700846
rect 41454 700436 41460 700500
rect 41524 700498 41530 700500
rect 41781 700498 41847 700501
rect 41524 700496 41847 700498
rect 41524 700440 41786 700496
rect 41842 700440 41847 700496
rect 41524 700438 41847 700440
rect 41524 700436 41530 700438
rect 41781 700435 41847 700438
rect 64646 700314 64706 700846
rect 61377 699682 61443 699685
rect 61377 699680 64706 699682
rect 61377 699624 61382 699680
rect 61438 699624 64706 699680
rect 61377 699622 64706 699624
rect 61377 699619 61443 699622
rect 64646 699132 64706 699622
rect 669405 698322 669471 698325
rect 675109 698322 675175 698325
rect 669405 698320 675175 698322
rect 669405 698264 669410 698320
rect 669466 698264 675114 698320
rect 675170 698264 675175 698320
rect 669405 698262 675175 698264
rect 669405 698259 669471 698262
rect 675109 698259 675175 698262
rect 62113 698186 62179 698189
rect 62113 698184 64706 698186
rect 62113 698128 62118 698184
rect 62174 698128 64706 698184
rect 62113 698126 64706 698128
rect 62113 698123 62179 698126
rect 64646 697950 64706 698126
rect 669221 697370 669287 697373
rect 675109 697370 675175 697373
rect 669221 697368 675175 697370
rect 669221 697312 669226 697368
rect 669282 697312 675114 697368
rect 675170 697312 675175 697368
rect 669221 697310 675175 697312
rect 669221 697307 669287 697310
rect 675109 697307 675175 697310
rect 673545 697098 673611 697101
rect 675109 697098 675175 697101
rect 673545 697096 675175 697098
rect 673545 697040 673550 697096
rect 673606 697040 675114 697096
rect 675170 697040 675175 697096
rect 673545 697038 675175 697040
rect 673545 697035 673611 697038
rect 675109 697035 675175 697038
rect 675385 696828 675451 696829
rect 675334 696826 675340 696828
rect 675294 696766 675340 696826
rect 675404 696824 675451 696828
rect 675446 696768 675451 696824
rect 675334 696764 675340 696766
rect 675404 696764 675451 696768
rect 675385 696763 675451 696764
rect 672993 695602 673059 695605
rect 674925 695602 674991 695605
rect 672993 695600 674991 695602
rect 672993 695544 672998 695600
rect 673054 695544 674930 695600
rect 674986 695544 674991 695600
rect 672993 695542 674991 695544
rect 672993 695539 673059 695542
rect 674925 695539 674991 695542
rect 672533 694650 672599 694653
rect 675109 694650 675175 694653
rect 672533 694648 675175 694650
rect 672533 694592 672538 694648
rect 672594 694592 675114 694648
rect 675170 694592 675175 694648
rect 672533 694590 675175 694592
rect 672533 694587 672599 694590
rect 675109 694587 675175 694590
rect 672165 690570 672231 690573
rect 675109 690570 675175 690573
rect 672165 690568 675175 690570
rect 672165 690512 672170 690568
rect 672226 690512 675114 690568
rect 675170 690512 675175 690568
rect 672165 690510 675175 690512
rect 672165 690507 672231 690510
rect 675109 690507 675175 690510
rect 673545 690026 673611 690029
rect 674925 690026 674991 690029
rect 673545 690024 674991 690026
rect 649950 689482 650010 689980
rect 673545 689968 673550 690024
rect 673606 689968 674930 690024
rect 674986 689968 674991 690024
rect 673545 689966 674991 689968
rect 673545 689963 673611 689966
rect 674925 689963 674991 689966
rect 651649 689482 651715 689485
rect 649950 689480 651715 689482
rect 649950 689424 651654 689480
rect 651710 689424 651715 689480
rect 649950 689422 651715 689424
rect 651649 689419 651715 689422
rect 674097 689210 674163 689213
rect 675109 689210 675175 689213
rect 674097 689208 675175 689210
rect 674097 689152 674102 689208
rect 674158 689152 675114 689208
rect 675170 689152 675175 689208
rect 674097 689150 675175 689152
rect 674097 689147 674163 689150
rect 675109 689147 675175 689150
rect 649980 688802 650562 688828
rect 651465 688802 651531 688805
rect 649980 688800 651531 688802
rect 649980 688768 651470 688800
rect 650502 688744 651470 688768
rect 651526 688744 651531 688800
rect 650502 688742 651531 688744
rect 651465 688739 651531 688742
rect 670785 688530 670851 688533
rect 675109 688530 675175 688533
rect 670785 688528 675175 688530
rect 670785 688472 670790 688528
rect 670846 688472 675114 688528
rect 675170 688472 675175 688528
rect 670785 688470 675175 688472
rect 670785 688467 670851 688470
rect 675109 688467 675175 688470
rect 42701 688122 42767 688125
rect 41492 688120 42767 688122
rect 41492 688064 42706 688120
rect 42762 688064 42767 688120
rect 41492 688062 42767 688064
rect 42701 688059 42767 688062
rect 44817 687714 44883 687717
rect 41492 687712 44883 687714
rect 41492 687656 44822 687712
rect 44878 687656 44883 687712
rect 41492 687654 44883 687656
rect 44817 687651 44883 687654
rect 673545 687714 673611 687717
rect 675293 687714 675359 687717
rect 673545 687712 675359 687714
rect 673545 687656 673550 687712
rect 673606 687656 675298 687712
rect 675354 687656 675359 687712
rect 673545 687654 675359 687656
rect 673545 687651 673611 687654
rect 675293 687651 675359 687654
rect 43437 687306 43503 687309
rect 41492 687304 43503 687306
rect 41492 687248 43442 687304
rect 43498 687248 43503 687304
rect 41492 687246 43503 687248
rect 649950 687306 650010 687616
rect 652017 687306 652083 687309
rect 649950 687304 652083 687306
rect 649950 687248 652022 687304
rect 652078 687248 652083 687304
rect 649950 687246 652083 687248
rect 43437 687243 43503 687246
rect 652017 687243 652083 687246
rect 674925 687170 674991 687173
rect 675334 687170 675340 687172
rect 674925 687168 675340 687170
rect 674925 687112 674930 687168
rect 674986 687112 675340 687168
rect 674925 687110 675340 687112
rect 674925 687107 674991 687110
rect 675334 687108 675340 687110
rect 675404 687108 675410 687172
rect 40861 686898 40927 686901
rect 651465 686898 651531 686901
rect 40861 686896 40940 686898
rect 40861 686840 40866 686896
rect 40922 686840 40940 686896
rect 40861 686838 40940 686840
rect 649950 686896 651531 686898
rect 649950 686840 651470 686896
rect 651526 686840 651531 686896
rect 649950 686838 651531 686840
rect 40861 686835 40927 686838
rect 41137 686490 41203 686493
rect 41124 686488 41203 686490
rect 41124 686432 41142 686488
rect 41198 686432 41203 686488
rect 649950 686434 650010 686838
rect 651465 686835 651531 686838
rect 41124 686430 41203 686432
rect 41137 686427 41203 686430
rect 675753 686218 675819 686221
rect 676990 686218 676996 686220
rect 675753 686216 676996 686218
rect 675753 686160 675758 686216
rect 675814 686160 676996 686216
rect 675753 686158 676996 686160
rect 675753 686155 675819 686158
rect 676990 686156 676996 686158
rect 677060 686156 677066 686220
rect 43069 686082 43135 686085
rect 41492 686080 43135 686082
rect 41492 686024 43074 686080
rect 43130 686024 43135 686080
rect 41492 686022 43135 686024
rect 43069 686019 43135 686022
rect 41045 685912 41111 685915
rect 41045 685910 41154 685912
rect 41045 685854 41050 685910
rect 41106 685854 41154 685910
rect 41045 685849 41154 685854
rect 41094 685644 41154 685849
rect 673177 685810 673243 685813
rect 675109 685810 675175 685813
rect 673177 685808 675175 685810
rect 673177 685752 673182 685808
rect 673238 685752 675114 685808
rect 675170 685752 675175 685808
rect 673177 685750 675175 685752
rect 673177 685747 673243 685750
rect 675109 685747 675175 685750
rect 668393 685538 668459 685541
rect 675477 685538 675543 685541
rect 668393 685536 675543 685538
rect 668393 685480 668398 685536
rect 668454 685480 675482 685536
rect 675538 685480 675543 685536
rect 668393 685478 675543 685480
rect 668393 685475 668459 685478
rect 675477 685475 675543 685478
rect 44265 685266 44331 685269
rect 651465 685266 651531 685269
rect 41492 685264 44331 685266
rect 41492 685208 44270 685264
rect 44326 685208 44331 685264
rect 41492 685206 44331 685208
rect 649950 685264 651531 685266
rect 649950 685208 651470 685264
rect 651526 685208 651531 685264
rect 649950 685206 651531 685208
rect 44265 685203 44331 685206
rect 651465 685203 651531 685206
rect 40861 684858 40927 684861
rect 40861 684856 40940 684858
rect 40861 684800 40866 684856
rect 40922 684800 40940 684856
rect 40861 684798 40940 684800
rect 40861 684795 40927 684798
rect 41689 684722 41755 684725
rect 44449 684722 44515 684725
rect 41689 684720 44515 684722
rect 41689 684664 41694 684720
rect 41750 684664 44454 684720
rect 44510 684664 44515 684720
rect 41689 684662 44515 684664
rect 41689 684659 41755 684662
rect 44449 684659 44515 684662
rect 45001 684450 45067 684453
rect 652569 684450 652635 684453
rect 41492 684448 45067 684450
rect 41492 684392 45006 684448
rect 45062 684392 45067 684448
rect 41492 684390 45067 684392
rect 45001 684387 45067 684390
rect 649950 684448 652635 684450
rect 649950 684392 652574 684448
rect 652630 684392 652635 684448
rect 649950 684390 652635 684392
rect 649950 684070 650010 684390
rect 652569 684387 652635 684390
rect 44265 684042 44331 684045
rect 41492 684040 44331 684042
rect 41492 683984 44270 684040
rect 44326 683984 44331 684040
rect 41492 683982 44331 683984
rect 44265 683979 44331 683982
rect 41822 683634 41828 683636
rect 41492 683574 41828 683634
rect 41822 683572 41828 683574
rect 41892 683572 41898 683636
rect 41321 683464 41387 683467
rect 41278 683462 41387 683464
rect 41278 683406 41326 683462
rect 41382 683406 41387 683462
rect 41278 683401 41387 683406
rect 41278 683196 41338 683401
rect 40953 682818 41019 682821
rect 40940 682816 41019 682818
rect 40940 682760 40958 682816
rect 41014 682760 41019 682816
rect 40940 682758 41019 682760
rect 40953 682755 41019 682758
rect 673637 682546 673703 682549
rect 675845 682546 675911 682549
rect 673637 682544 675911 682546
rect 673637 682488 673642 682544
rect 673698 682488 675850 682544
rect 675906 682488 675911 682544
rect 673637 682486 675911 682488
rect 673637 682483 673703 682486
rect 675845 682483 675911 682486
rect 42517 682410 42583 682413
rect 41492 682408 42583 682410
rect 41492 682352 42522 682408
rect 42578 682352 42583 682408
rect 41492 682350 42583 682352
rect 42517 682347 42583 682350
rect 673637 682274 673703 682277
rect 675661 682274 675727 682277
rect 673637 682272 675727 682274
rect 673637 682216 673642 682272
rect 673698 682216 675666 682272
rect 675722 682216 675727 682272
rect 673637 682214 675727 682216
rect 673637 682211 673703 682214
rect 675661 682211 675727 682214
rect 675886 682076 675892 682140
rect 675956 682138 675962 682140
rect 682377 682138 682443 682141
rect 675956 682136 682443 682138
rect 675956 682080 682382 682136
rect 682438 682080 682443 682136
rect 675956 682078 682443 682080
rect 675956 682076 675962 682078
rect 682377 682075 682443 682078
rect 35157 682002 35223 682005
rect 35157 682000 35236 682002
rect 35157 681944 35162 682000
rect 35218 681944 35236 682000
rect 35157 681942 35236 681944
rect 35157 681939 35223 681942
rect 676070 681804 676076 681868
rect 676140 681866 676146 681868
rect 678237 681866 678303 681869
rect 676140 681864 678303 681866
rect 676140 681808 678242 681864
rect 678298 681808 678303 681864
rect 676140 681806 678303 681808
rect 676140 681804 676146 681806
rect 678237 681803 678303 681806
rect 42241 681594 42307 681597
rect 41492 681592 42307 681594
rect 41492 681536 42246 681592
rect 42302 681536 42307 681592
rect 41492 681534 42307 681536
rect 42241 681531 42307 681534
rect 32397 681186 32463 681189
rect 32397 681184 32476 681186
rect 32397 681128 32402 681184
rect 32458 681128 32476 681184
rect 32397 681126 32476 681128
rect 32397 681123 32463 681126
rect 33777 680778 33843 680781
rect 33764 680776 33843 680778
rect 33764 680720 33782 680776
rect 33838 680720 33843 680776
rect 33764 680718 33843 680720
rect 33777 680715 33843 680718
rect 43621 680370 43687 680373
rect 41492 680368 43687 680370
rect 41492 680312 43626 680368
rect 43682 680312 43687 680368
rect 41492 680310 43687 680312
rect 43621 680307 43687 680310
rect 41137 679962 41203 679965
rect 41124 679960 41203 679962
rect 41124 679904 41142 679960
rect 41198 679904 41203 679960
rect 41124 679902 41203 679904
rect 41137 679899 41203 679902
rect 43989 679554 44055 679557
rect 41492 679552 44055 679554
rect 41492 679496 43994 679552
rect 44050 679496 44055 679552
rect 41492 679494 44055 679496
rect 43989 679491 44055 679494
rect 40542 678992 40602 679116
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678928 40794 678992
rect 40726 678708 40786 678928
rect 41781 678876 41847 678877
rect 41781 678872 41828 678876
rect 41892 678874 41898 678876
rect 41781 678816 41786 678872
rect 41781 678812 41828 678816
rect 41892 678814 41938 678874
rect 41892 678812 41898 678814
rect 41781 678811 41847 678812
rect 41781 678330 41847 678333
rect 41492 678328 41847 678330
rect 41492 678272 41786 678328
rect 41842 678272 41847 678328
rect 41492 678270 41847 678272
rect 41781 678267 41847 678270
rect 43069 677922 43135 677925
rect 41492 677920 43135 677922
rect 41492 677864 43074 677920
rect 43130 677864 43135 677920
rect 41492 677862 43135 677864
rect 43069 677859 43135 677862
rect 40953 677754 41019 677755
rect 40902 677752 40908 677754
rect 40862 677692 40908 677752
rect 40972 677750 41019 677754
rect 41014 677694 41019 677750
rect 40902 677690 40908 677692
rect 40972 677690 41019 677694
rect 40953 677689 41019 677690
rect 39990 677109 40050 677484
rect 39941 677104 40050 677109
rect 39941 677048 39946 677104
rect 40002 677076 40050 677104
rect 40002 677048 40020 677076
rect 39941 677046 40020 677048
rect 39941 677043 40007 677046
rect 43437 676698 43503 676701
rect 41492 676696 43503 676698
rect 41492 676640 43442 676696
rect 43498 676640 43503 676696
rect 41492 676638 43503 676640
rect 43437 676635 43503 676638
rect 675293 676426 675359 676429
rect 676070 676426 676076 676428
rect 675293 676424 676076 676426
rect 675293 676368 675298 676424
rect 675354 676368 676076 676424
rect 675293 676366 676076 676368
rect 675293 676363 675359 676366
rect 676070 676364 676076 676366
rect 676140 676364 676146 676428
rect 39941 673026 40007 673029
rect 41086 673026 41092 673028
rect 39941 673024 41092 673026
rect 39941 672968 39946 673024
rect 40002 672968 41092 673024
rect 39941 672966 41092 672968
rect 39941 672963 40007 672966
rect 41086 672964 41092 672966
rect 41156 672964 41162 673028
rect 32397 672754 32463 672757
rect 41822 672754 41828 672756
rect 32397 672752 41828 672754
rect 32397 672696 32402 672752
rect 32458 672696 41828 672752
rect 32397 672694 41828 672696
rect 32397 672691 32463 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 43253 671940 43319 671941
rect 43253 671936 43300 671940
rect 43364 671938 43370 671940
rect 43253 671880 43258 671936
rect 43253 671876 43300 671880
rect 43364 671878 43410 671938
rect 43364 671876 43370 671878
rect 43253 671875 43319 671876
rect 673637 671394 673703 671397
rect 673637 671392 676292 671394
rect 673637 671336 673642 671392
rect 673698 671336 676292 671392
rect 673637 671334 676292 671336
rect 673637 671331 673703 671334
rect 38929 671258 38995 671261
rect 42793 671258 42859 671261
rect 38929 671256 42859 671258
rect 38929 671200 38934 671256
rect 38990 671200 42798 671256
rect 42854 671200 42859 671256
rect 38929 671198 42859 671200
rect 38929 671195 38995 671198
rect 42793 671195 42859 671198
rect 38193 670986 38259 670989
rect 40350 670986 40356 670988
rect 38193 670984 40356 670986
rect 38193 670928 38198 670984
rect 38254 670928 40356 670984
rect 38193 670926 40356 670928
rect 38193 670923 38259 670926
rect 40350 670924 40356 670926
rect 40420 670924 40426 670988
rect 674005 670986 674071 670989
rect 674005 670984 676292 670986
rect 674005 670928 674010 670984
rect 674066 670928 676292 670984
rect 674005 670926 676292 670928
rect 674005 670923 674071 670926
rect 673637 670578 673703 670581
rect 673637 670576 676292 670578
rect 673637 670520 673642 670576
rect 673698 670520 676292 670576
rect 673637 670518 676292 670520
rect 673637 670515 673703 670518
rect 674005 670170 674071 670173
rect 674005 670168 676292 670170
rect 674005 670112 674010 670168
rect 674066 670112 676292 670168
rect 674005 670110 676292 670112
rect 674005 670107 674071 670110
rect 674005 669762 674071 669765
rect 674005 669760 676292 669762
rect 674005 669704 674010 669760
rect 674066 669704 676292 669760
rect 674005 669702 676292 669704
rect 674005 669699 674071 669702
rect 673361 669490 673427 669493
rect 673361 669488 676322 669490
rect 673361 669432 673366 669488
rect 673422 669432 676322 669488
rect 673361 669430 676322 669432
rect 673361 669427 673427 669430
rect 676262 669324 676322 669430
rect 41086 669020 41092 669084
rect 41156 669082 41162 669084
rect 41781 669082 41847 669085
rect 41156 669080 41847 669082
rect 41156 669024 41786 669080
rect 41842 669024 41847 669080
rect 41156 669022 41847 669024
rect 41156 669020 41162 669022
rect 41781 669019 41847 669022
rect 673637 668946 673703 668949
rect 673637 668944 676292 668946
rect 673637 668888 673642 668944
rect 673698 668888 676292 668944
rect 673637 668886 676292 668888
rect 673637 668883 673703 668886
rect 674005 668538 674071 668541
rect 674005 668536 676292 668538
rect 674005 668480 674010 668536
rect 674066 668480 676292 668536
rect 674005 668478 676292 668480
rect 674005 668475 674071 668478
rect 674005 668130 674071 668133
rect 674005 668128 676292 668130
rect 674005 668072 674010 668128
rect 674066 668072 676292 668128
rect 674005 668070 676292 668072
rect 674005 668067 674071 668070
rect 674005 667722 674071 667725
rect 674005 667720 676292 667722
rect 674005 667664 674010 667720
rect 674066 667664 676292 667720
rect 674005 667662 676292 667664
rect 674005 667659 674071 667662
rect 42190 667388 42196 667452
rect 42260 667450 42266 667452
rect 45001 667450 45067 667453
rect 42260 667448 45067 667450
rect 42260 667392 45006 667448
rect 45062 667392 45067 667448
rect 42260 667390 45067 667392
rect 42260 667388 42266 667390
rect 45001 667387 45067 667390
rect 673637 667314 673703 667317
rect 673637 667312 676292 667314
rect 673637 667256 673642 667312
rect 673698 667256 676292 667312
rect 673637 667254 676292 667256
rect 673637 667251 673703 667254
rect 678237 667042 678303 667045
rect 678237 667040 678346 667042
rect 678237 666984 678242 667040
rect 678298 666984 678346 667040
rect 678237 666979 678346 666984
rect 43294 666844 43300 666908
rect 43364 666844 43370 666908
rect 678286 666876 678346 666979
rect 42149 666636 42215 666637
rect 42149 666634 42196 666636
rect 42104 666632 42196 666634
rect 42104 666576 42154 666632
rect 42104 666574 42196 666576
rect 42149 666572 42196 666574
rect 42260 666572 42266 666636
rect 43302 666573 43362 666844
rect 682377 666634 682443 666637
rect 42149 666571 42215 666572
rect 43253 666568 43362 666573
rect 43253 666512 43258 666568
rect 43314 666512 43362 666568
rect 43253 666510 43362 666512
rect 682334 666632 682443 666634
rect 682334 666576 682382 666632
rect 682438 666576 682443 666632
rect 682334 666571 682443 666576
rect 43253 666507 43319 666510
rect 682334 666468 682394 666571
rect 673637 666090 673703 666093
rect 673637 666088 676292 666090
rect 673637 666032 673642 666088
rect 673698 666032 676292 666088
rect 673637 666030 676292 666032
rect 673637 666027 673703 666030
rect 42057 665954 42123 665957
rect 45737 665954 45803 665957
rect 42057 665952 45803 665954
rect 42057 665896 42062 665952
rect 42118 665896 45742 665952
rect 45798 665896 45803 665952
rect 42057 665894 45803 665896
rect 42057 665891 42123 665894
rect 45737 665891 45803 665894
rect 674005 665682 674071 665685
rect 674005 665680 676292 665682
rect 674005 665624 674010 665680
rect 674066 665624 676292 665680
rect 674005 665622 676292 665624
rect 674005 665619 674071 665622
rect 40350 665484 40356 665548
rect 40420 665546 40426 665548
rect 42425 665546 42491 665549
rect 40420 665544 42491 665546
rect 40420 665488 42430 665544
rect 42486 665488 42491 665544
rect 40420 665486 42491 665488
rect 40420 665484 40426 665486
rect 42425 665483 42491 665486
rect 683205 665410 683271 665413
rect 683205 665408 683314 665410
rect 683205 665352 683210 665408
rect 683266 665352 683314 665408
rect 683205 665347 683314 665352
rect 40902 665212 40908 665276
rect 40972 665274 40978 665276
rect 42241 665274 42307 665277
rect 40972 665272 42307 665274
rect 40972 665216 42246 665272
rect 42302 665216 42307 665272
rect 683254 665244 683314 665347
rect 40972 665214 42307 665216
rect 40972 665212 40978 665214
rect 42241 665211 42307 665214
rect 673637 664866 673703 664869
rect 673637 664864 676292 664866
rect 673637 664808 673642 664864
rect 673698 664808 676292 664864
rect 673637 664806 676292 664808
rect 673637 664803 673703 664806
rect 673361 664186 673427 664189
rect 676262 664186 676322 664428
rect 673361 664184 676322 664186
rect 673361 664128 673366 664184
rect 673422 664128 676322 664184
rect 673361 664126 676322 664128
rect 673361 664123 673427 664126
rect 676806 664124 676812 664188
rect 676876 664124 676882 664188
rect 40718 663988 40724 664052
rect 40788 664050 40794 664052
rect 41781 664050 41847 664053
rect 40788 664048 41847 664050
rect 40788 663992 41786 664048
rect 41842 663992 41847 664048
rect 676814 664020 676874 664124
rect 40788 663990 41847 663992
rect 40788 663988 40794 663990
rect 41781 663987 41847 663990
rect 672717 663914 672783 663917
rect 673637 663914 673703 663917
rect 672717 663912 673703 663914
rect 672717 663856 672722 663912
rect 672778 663856 673642 663912
rect 673698 663856 673703 663912
rect 672717 663854 673703 663856
rect 672717 663851 672783 663854
rect 673637 663851 673703 663854
rect 674005 663642 674071 663645
rect 674005 663640 676292 663642
rect 674005 663584 674010 663640
rect 674066 663584 676292 663640
rect 674005 663582 676292 663584
rect 674005 663579 674071 663582
rect 683389 663370 683455 663373
rect 683389 663368 683498 663370
rect 683389 663312 683394 663368
rect 683450 663312 683498 663368
rect 683389 663307 683498 663312
rect 683438 663204 683498 663307
rect 42057 662826 42123 662829
rect 41370 662824 42123 662826
rect 41370 662768 42062 662824
rect 42118 662768 42123 662824
rect 41370 662766 42123 662768
rect 40534 662628 40540 662692
rect 40604 662690 40610 662692
rect 41370 662690 41430 662766
rect 42057 662763 42123 662766
rect 674005 662826 674071 662829
rect 674005 662824 676292 662826
rect 674005 662768 674010 662824
rect 674066 662768 676292 662824
rect 674005 662766 676292 662768
rect 674005 662763 674071 662766
rect 40604 662630 41430 662690
rect 40604 662628 40610 662630
rect 674414 662356 674420 662420
rect 674484 662418 674490 662420
rect 674484 662358 676292 662418
rect 674484 662356 674490 662358
rect 673821 662010 673887 662013
rect 673821 662008 676292 662010
rect 673821 661952 673826 662008
rect 673882 661952 676292 662008
rect 673821 661950 676292 661952
rect 673821 661947 673887 661950
rect 674005 661602 674071 661605
rect 674005 661600 676292 661602
rect 674005 661544 674010 661600
rect 674066 661544 676292 661600
rect 674005 661542 676292 661544
rect 674005 661539 674071 661542
rect 674005 661194 674071 661197
rect 674005 661192 676292 661194
rect 674005 661136 674010 661192
rect 674066 661136 676292 661192
rect 674005 661134 676292 661136
rect 674005 661131 674071 661134
rect 41454 660860 41460 660924
rect 41524 660922 41530 660924
rect 42701 660922 42767 660925
rect 41524 660920 42767 660922
rect 41524 660864 42706 660920
rect 42762 660864 42767 660920
rect 41524 660862 42767 660864
rect 41524 660860 41530 660862
rect 42701 660859 42767 660862
rect 62113 660922 62179 660925
rect 62113 660920 64706 660922
rect 62113 660864 62118 660920
rect 62174 660864 64706 660920
rect 62113 660862 64706 660864
rect 62113 660859 62179 660862
rect 64646 660638 64706 660862
rect 683070 660109 683130 660756
rect 674005 660106 674071 660109
rect 675845 660106 675911 660109
rect 674005 660104 675911 660106
rect 674005 660048 674010 660104
rect 674066 660048 675850 660104
rect 675906 660048 675911 660104
rect 674005 660046 675911 660048
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 674005 660043 674071 660046
rect 675845 660043 675911 660046
rect 683113 660043 683179 660046
rect 673269 659698 673335 659701
rect 676262 659698 676322 659940
rect 673269 659696 676322 659698
rect 673269 659640 673274 659696
rect 673330 659640 676322 659696
rect 673269 659638 676322 659640
rect 673269 659635 673335 659638
rect 62113 659562 62179 659565
rect 62113 659560 64706 659562
rect 62113 659504 62118 659560
rect 62174 659504 64706 659560
rect 62113 659502 64706 659504
rect 62113 659499 62179 659502
rect 64646 659456 64706 659502
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42517 658610 42583 658613
rect 41708 658608 42583 658610
rect 41708 658552 42522 658608
rect 42578 658552 42583 658608
rect 41708 658550 42583 658552
rect 41708 658548 41714 658550
rect 42517 658547 42583 658550
rect 41781 658340 41847 658341
rect 41781 658336 41828 658340
rect 41892 658338 41898 658340
rect 62113 658338 62179 658341
rect 41781 658280 41786 658336
rect 41781 658276 41828 658280
rect 41892 658278 41938 658338
rect 62113 658336 64706 658338
rect 62113 658280 62118 658336
rect 62174 658280 64706 658336
rect 62113 658278 64706 658280
rect 41892 658276 41898 658278
rect 41781 658275 41847 658276
rect 62113 658275 62179 658278
rect 64646 658274 64706 658278
rect 62757 657658 62823 657661
rect 62757 657656 64706 657658
rect 62757 657600 62762 657656
rect 62818 657600 64706 657656
rect 62757 657598 64706 657600
rect 62757 657595 62823 657598
rect 64646 657092 64706 657598
rect 61377 656570 61443 656573
rect 61377 656568 64706 656570
rect 61377 656512 61382 656568
rect 61438 656512 64706 656568
rect 61377 656510 64706 656512
rect 61377 656507 61443 656510
rect 64646 655910 64706 656510
rect 674005 655618 674071 655621
rect 675109 655618 675175 655621
rect 674005 655616 675175 655618
rect 674005 655560 674010 655616
rect 674066 655560 675114 655616
rect 675170 655560 675175 655616
rect 674005 655558 675175 655560
rect 674005 655555 674071 655558
rect 675109 655555 675175 655558
rect 62113 655346 62179 655349
rect 62113 655344 64706 655346
rect 62113 655288 62118 655344
rect 62174 655288 64706 655344
rect 62113 655286 64706 655288
rect 62113 655283 62179 655286
rect 64646 654728 64706 655286
rect 674005 654122 674071 654125
rect 674925 654122 674991 654125
rect 674005 654120 674991 654122
rect 674005 654064 674010 654120
rect 674066 654064 674930 654120
rect 674986 654064 674991 654120
rect 674005 654062 674991 654064
rect 674005 654059 674071 654062
rect 674925 654059 674991 654062
rect 671981 652898 672047 652901
rect 675385 652898 675451 652901
rect 671981 652896 675451 652898
rect 671981 652840 671986 652896
rect 672042 652840 675390 652896
rect 675446 652840 675451 652896
rect 671981 652838 675451 652840
rect 671981 652835 672047 652838
rect 675385 652835 675451 652838
rect 672717 651402 672783 651405
rect 675109 651402 675175 651405
rect 672717 651400 675175 651402
rect 672717 651344 672722 651400
rect 672778 651344 675114 651400
rect 675170 651344 675175 651400
rect 672717 651342 675175 651344
rect 672717 651339 672783 651342
rect 675109 651339 675175 651342
rect 674230 649708 674236 649772
rect 674300 649770 674306 649772
rect 675385 649770 675451 649773
rect 674300 649768 675451 649770
rect 674300 649712 675390 649768
rect 675446 649712 675451 649768
rect 674300 649710 675451 649712
rect 674300 649708 674306 649710
rect 675385 649707 675451 649710
rect 673637 649226 673703 649229
rect 675385 649226 675451 649229
rect 673637 649224 675451 649226
rect 673637 649168 673642 649224
rect 673698 649168 675390 649224
rect 675446 649168 675451 649224
rect 673637 649166 675451 649168
rect 673637 649163 673703 649166
rect 675385 649163 675451 649166
rect 675753 648682 675819 648685
rect 676806 648682 676812 648684
rect 675753 648680 676812 648682
rect 675753 648624 675758 648680
rect 675814 648624 676812 648680
rect 675753 648622 676812 648624
rect 675753 648619 675819 648622
rect 676806 648620 676812 648622
rect 676876 648620 676882 648684
rect 669037 647866 669103 647869
rect 675385 647866 675451 647869
rect 669037 647864 675451 647866
rect 669037 647808 669042 647864
rect 669098 647808 675390 647864
rect 675446 647808 675451 647864
rect 669037 647806 675451 647808
rect 669037 647803 669103 647806
rect 675385 647803 675451 647806
rect 674005 647322 674071 647325
rect 675109 647322 675175 647325
rect 674005 647320 675175 647322
rect 674005 647264 674010 647320
rect 674066 647264 675114 647320
rect 675170 647264 675175 647320
rect 674005 647262 675175 647264
rect 674005 647259 674071 647262
rect 675109 647259 675175 647262
rect 35758 644741 35818 644912
rect 35758 644736 35867 644741
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644678 35867 644680
rect 35801 644675 35867 644678
rect 40125 644738 40191 644741
rect 44449 644738 44515 644741
rect 40125 644736 44515 644738
rect 40125 644680 40130 644736
rect 40186 644680 44454 644736
rect 44510 644680 44515 644736
rect 40125 644678 44515 644680
rect 40125 644675 40191 644678
rect 44449 644675 44515 644678
rect 673821 644738 673887 644741
rect 675293 644738 675359 644741
rect 673821 644736 675359 644738
rect 673821 644680 673826 644736
rect 673882 644680 675298 644736
rect 675354 644680 675359 644736
rect 673821 644678 675359 644680
rect 673821 644675 673887 644678
rect 675293 644675 675359 644678
rect 38518 644333 38578 644504
rect 38518 644328 38627 644333
rect 38518 644272 38566 644328
rect 38622 644272 38627 644328
rect 38518 644270 38627 644272
rect 38561 644267 38627 644270
rect 35390 643925 35450 644096
rect 674557 644058 674623 644061
rect 674782 644058 674788 644060
rect 674557 644056 674788 644058
rect 674557 644000 674562 644056
rect 674618 644000 674788 644056
rect 674557 643998 674788 644000
rect 674557 643995 674623 643998
rect 674782 643996 674788 643998
rect 674852 643996 674858 644060
rect 35341 643920 35450 643925
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 35341 643859 35407 643862
rect 35574 643517 35634 643688
rect 671153 643650 671219 643653
rect 675385 643650 675451 643653
rect 671153 643648 675451 643650
rect 671153 643592 671158 643648
rect 671214 643592 675390 643648
rect 675446 643592 675451 643648
rect 671153 643590 675451 643592
rect 671153 643587 671219 643590
rect 675385 643587 675451 643590
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 35758 643280 35818 643451
rect 649950 643242 650010 643558
rect 651465 643242 651531 643245
rect 649950 643240 651531 643242
rect 649950 643184 651470 643240
rect 651526 643184 651531 643240
rect 649950 643182 651531 643184
rect 651465 643179 651531 643182
rect 39941 643106 40007 643109
rect 44725 643106 44791 643109
rect 39941 643104 44791 643106
rect 39941 643048 39946 643104
rect 40002 643048 44730 643104
rect 44786 643048 44791 643104
rect 39941 643046 44791 643048
rect 39941 643043 40007 643046
rect 44725 643043 44791 643046
rect 674005 643106 674071 643109
rect 675109 643106 675175 643109
rect 674005 643104 675175 643106
rect 674005 643048 674010 643104
rect 674066 643048 675114 643104
rect 675170 643048 675175 643104
rect 674005 643046 675175 643048
rect 674005 643043 674071 643046
rect 675109 643043 675175 643046
rect 35574 642701 35634 642872
rect 35574 642696 35683 642701
rect 35574 642640 35622 642696
rect 35678 642640 35683 642696
rect 35574 642638 35683 642640
rect 35617 642635 35683 642638
rect 35801 642290 35867 642293
rect 35758 642288 35867 642290
rect 35758 642232 35806 642288
rect 35862 642232 35867 642288
rect 35758 642227 35867 642232
rect 41462 642290 41522 642464
rect 44214 642290 44220 642292
rect 41462 642230 44220 642290
rect 44214 642228 44220 642230
rect 44284 642228 44290 642292
rect 35758 642056 35818 642227
rect 649950 641882 650010 642376
rect 652017 641882 652083 641885
rect 649950 641880 652083 641882
rect 649950 641824 652022 641880
rect 652078 641824 652083 641880
rect 649950 641822 652083 641824
rect 652017 641819 652083 641822
rect 671797 641746 671863 641749
rect 675293 641746 675359 641749
rect 671797 641744 675359 641746
rect 671797 641688 671802 641744
rect 671858 641688 675298 641744
rect 675354 641688 675359 641744
rect 671797 641686 675359 641688
rect 671797 641683 671863 641686
rect 675293 641683 675359 641686
rect 35390 641477 35450 641648
rect 35390 641472 35499 641477
rect 35390 641416 35438 641472
rect 35494 641416 35499 641472
rect 35390 641414 35499 641416
rect 35433 641411 35499 641414
rect 35758 641069 35818 641240
rect 35758 641064 35867 641069
rect 35758 641008 35806 641064
rect 35862 641008 35867 641064
rect 35758 641006 35867 641008
rect 35801 641003 35867 641006
rect 39757 641066 39823 641069
rect 44265 641066 44331 641069
rect 39757 641064 44331 641066
rect 39757 641008 39762 641064
rect 39818 641008 44270 641064
rect 44326 641008 44331 641064
rect 39757 641006 44331 641008
rect 39757 641003 39823 641006
rect 44265 641003 44331 641006
rect 35574 640661 35634 640832
rect 649950 640794 650010 641194
rect 651465 640794 651531 640797
rect 649950 640792 651531 640794
rect 649950 640736 651470 640792
rect 651526 640736 651531 640792
rect 649950 640734 651531 640736
rect 651465 640731 651531 640734
rect 35574 640656 35683 640661
rect 41638 640658 41644 640660
rect 35574 640600 35622 640656
rect 35678 640600 35683 640656
rect 35574 640598 35683 640600
rect 35617 640595 35683 640598
rect 41462 640598 41644 640658
rect 41462 640424 41522 640598
rect 41638 640596 41644 640598
rect 41708 640596 41714 640660
rect 40033 640250 40099 640253
rect 45093 640250 45159 640253
rect 40033 640248 45159 640250
rect 40033 640192 40038 640248
rect 40094 640192 45098 640248
rect 45154 640192 45159 640248
rect 40033 640190 45159 640192
rect 40033 640187 40099 640190
rect 45093 640187 45159 640190
rect 674465 640250 674531 640253
rect 674782 640250 674788 640252
rect 674465 640248 674788 640250
rect 674465 640192 674470 640248
rect 674526 640192 674788 640248
rect 674465 640190 674788 640192
rect 674465 640187 674531 640190
rect 674782 640188 674788 640190
rect 674852 640188 674858 640252
rect 651373 640114 651439 640117
rect 649950 640112 651439 640114
rect 649950 640056 651378 640112
rect 651434 640056 651439 640112
rect 649950 640054 651439 640056
rect 35758 639845 35818 640016
rect 649950 640012 650010 640054
rect 651373 640051 651439 640054
rect 35758 639840 35867 639845
rect 35758 639784 35806 639840
rect 35862 639784 35867 639840
rect 35758 639782 35867 639784
rect 35801 639779 35867 639782
rect 41462 639436 41522 639608
rect 41454 639372 41460 639436
rect 41524 639372 41530 639436
rect 35758 639029 35818 639200
rect 35758 639024 35867 639029
rect 35758 638968 35806 639024
rect 35862 638968 35867 639024
rect 35758 638966 35867 638968
rect 35801 638963 35867 638966
rect 35574 638621 35634 638792
rect 35574 638616 35683 638621
rect 35574 638560 35622 638616
rect 35678 638560 35683 638616
rect 35574 638558 35683 638560
rect 649766 638618 649826 638830
rect 668853 638754 668919 638757
rect 675477 638754 675543 638757
rect 668853 638752 675543 638754
rect 668853 638696 668858 638752
rect 668914 638696 675482 638752
rect 675538 638696 675543 638752
rect 668853 638694 675543 638696
rect 668853 638691 668919 638694
rect 675477 638691 675543 638694
rect 651465 638618 651531 638621
rect 649766 638616 651531 638618
rect 649766 638560 651470 638616
rect 651526 638560 651531 638616
rect 649766 638558 651531 638560
rect 35617 638555 35683 638558
rect 651465 638555 651531 638558
rect 35758 638213 35818 638384
rect 35758 638208 35867 638213
rect 651649 638210 651715 638213
rect 35758 638152 35806 638208
rect 35862 638152 35867 638208
rect 35758 638150 35867 638152
rect 35801 638147 35867 638150
rect 649950 638208 651715 638210
rect 649950 638152 651654 638208
rect 651710 638152 651715 638208
rect 649950 638150 651715 638152
rect 35206 637805 35266 637976
rect 35157 637800 35266 637805
rect 35157 637744 35162 637800
rect 35218 637744 35266 637800
rect 35157 637742 35266 637744
rect 35157 637739 35223 637742
rect 649950 637648 650010 638150
rect 651649 638147 651715 638150
rect 40542 637396 40602 637568
rect 40534 637332 40540 637396
rect 40604 637332 40610 637396
rect 31894 636989 31954 637160
rect 31894 636984 32003 636989
rect 31894 636928 31942 636984
rect 31998 636928 32003 636984
rect 31894 636926 32003 636928
rect 31937 636923 32003 636926
rect 674097 636850 674163 636853
rect 675845 636850 675911 636853
rect 674097 636848 675911 636850
rect 674097 636792 674102 636848
rect 674158 636792 675850 636848
rect 675906 636792 675911 636848
rect 674097 636790 675911 636792
rect 674097 636787 674163 636790
rect 675845 636787 675911 636790
rect 35574 636581 35634 636752
rect 35525 636576 35634 636581
rect 35801 636578 35867 636581
rect 35525 636520 35530 636576
rect 35586 636520 35634 636576
rect 35525 636518 35634 636520
rect 35758 636576 35867 636578
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35525 636515 35591 636518
rect 35758 636515 35867 636520
rect 40677 636578 40743 636581
rect 42701 636578 42767 636581
rect 40677 636576 42767 636578
rect 40677 636520 40682 636576
rect 40738 636520 42706 636576
rect 42762 636520 42767 636576
rect 40677 636518 42767 636520
rect 40677 636515 40743 636518
rect 42701 636515 42767 636518
rect 675477 636578 675543 636581
rect 683205 636578 683271 636581
rect 675477 636576 683271 636578
rect 675477 636520 675482 636576
rect 675538 636520 683210 636576
rect 683266 636520 683271 636576
rect 675477 636518 683271 636520
rect 675477 636515 675543 636518
rect 683205 636515 683271 636518
rect 35758 636344 35818 636515
rect 39849 636170 39915 636173
rect 43989 636170 44055 636173
rect 39849 636168 44055 636170
rect 39849 636112 39854 636168
rect 39910 636112 43994 636168
rect 44050 636112 44055 636168
rect 39849 636110 44055 636112
rect 39849 636107 39915 636110
rect 43989 636107 44055 636110
rect 676070 636108 676076 636172
rect 676140 636170 676146 636172
rect 680997 636170 681063 636173
rect 676140 636168 681063 636170
rect 676140 636112 681002 636168
rect 681058 636112 681063 636168
rect 676140 636110 681063 636112
rect 676140 636108 676146 636110
rect 680997 636107 681063 636110
rect 35758 635765 35818 635936
rect 35758 635760 35867 635765
rect 35758 635704 35806 635760
rect 35862 635704 35867 635760
rect 35758 635702 35867 635704
rect 35801 635699 35867 635702
rect 40726 635356 40786 635528
rect 40718 635292 40724 635356
rect 40788 635292 40794 635356
rect 40910 634948 40970 635120
rect 40902 634884 40908 634948
rect 40972 634884 40978 634948
rect 41597 634946 41663 634949
rect 44357 634946 44423 634949
rect 41597 634944 44423 634946
rect 41597 634888 41602 634944
rect 41658 634888 44362 634944
rect 44418 634888 44423 634944
rect 41597 634886 44423 634888
rect 41597 634883 41663 634886
rect 44357 634883 44423 634886
rect 35574 634541 35634 634712
rect 35574 634536 35683 634541
rect 35574 634480 35622 634536
rect 35678 634480 35683 634536
rect 35574 634478 35683 634480
rect 35617 634475 35683 634478
rect 38518 633725 38578 634304
rect 35801 633722 35867 633725
rect 35758 633720 35867 633722
rect 35758 633664 35806 633720
rect 35862 633664 35867 633720
rect 35758 633659 35867 633664
rect 38518 633720 38627 633725
rect 38518 633664 38566 633720
rect 38622 633664 38627 633720
rect 38518 633662 38627 633664
rect 38561 633659 38627 633662
rect 35758 633488 35818 633659
rect 41413 632906 41479 632909
rect 42374 632906 42380 632908
rect 41413 632904 42380 632906
rect 41413 632848 41418 632904
rect 41474 632848 42380 632904
rect 41413 632846 42380 632848
rect 41413 632843 41479 632846
rect 42374 632844 42380 632846
rect 42444 632844 42450 632908
rect 40125 631954 40191 631957
rect 43621 631954 43687 631957
rect 40125 631952 43687 631954
rect 40125 631896 40130 631952
rect 40186 631896 43626 631952
rect 43682 631896 43687 631952
rect 40125 631894 43687 631896
rect 40125 631891 40191 631894
rect 43621 631891 43687 631894
rect 37917 631410 37983 631413
rect 42609 631410 42675 631413
rect 37917 631408 42675 631410
rect 37917 631352 37922 631408
rect 37978 631352 42614 631408
rect 42670 631352 42675 631408
rect 37917 631350 42675 631352
rect 37917 631347 37983 631350
rect 42609 631347 42675 631350
rect 39573 630730 39639 630733
rect 44909 630730 44975 630733
rect 39573 630728 44975 630730
rect 39573 630672 39578 630728
rect 39634 630672 44914 630728
rect 44970 630672 44975 630728
rect 39573 630670 44975 630672
rect 39573 630667 39639 630670
rect 44909 630667 44975 630670
rect 35157 629914 35223 629917
rect 41822 629914 41828 629916
rect 35157 629912 41828 629914
rect 35157 629856 35162 629912
rect 35218 629856 41828 629912
rect 35157 629854 41828 629856
rect 35157 629851 35223 629854
rect 41822 629852 41828 629854
rect 41892 629852 41898 629916
rect 40217 629234 40283 629237
rect 42149 629234 42215 629237
rect 40217 629232 42215 629234
rect 40217 629176 40222 629232
rect 40278 629176 42154 629232
rect 42210 629176 42215 629232
rect 40217 629174 42215 629176
rect 40217 629171 40283 629174
rect 42149 629171 42215 629174
rect 42333 628316 42399 628319
rect 42333 628314 42442 628316
rect 40493 628282 40559 628285
rect 42333 628282 42338 628314
rect 40493 628280 42338 628282
rect 40493 628224 40498 628280
rect 40554 628258 42338 628280
rect 42394 628258 42442 628314
rect 40554 628224 42442 628258
rect 40493 628222 42442 628224
rect 40493 628219 40559 628222
rect 674741 626650 674807 626653
rect 675845 626650 675911 626653
rect 674741 626648 675911 626650
rect 674741 626592 674746 626648
rect 674802 626592 675850 626648
rect 675906 626592 675911 626648
rect 674741 626590 675911 626592
rect 674741 626587 674807 626590
rect 675845 626587 675911 626590
rect 674005 626378 674071 626381
rect 674005 626376 676292 626378
rect 674005 626320 674010 626376
rect 674066 626320 676292 626376
rect 674005 626318 676292 626320
rect 674005 626315 674071 626318
rect 673453 625970 673519 625973
rect 673453 625968 676292 625970
rect 673453 625912 673458 625968
rect 673514 625912 676292 625968
rect 673453 625910 676292 625912
rect 673453 625907 673519 625910
rect 42241 625700 42307 625701
rect 42190 625636 42196 625700
rect 42260 625698 42307 625700
rect 42260 625696 42352 625698
rect 42302 625640 42352 625696
rect 42260 625638 42352 625640
rect 42260 625636 42307 625638
rect 42241 625635 42307 625636
rect 674005 625562 674071 625565
rect 674005 625560 676292 625562
rect 674005 625504 674010 625560
rect 674066 625504 676292 625560
rect 674005 625502 676292 625504
rect 674005 625499 674071 625502
rect 674005 625154 674071 625157
rect 674005 625152 676292 625154
rect 674005 625096 674010 625152
rect 674066 625096 676292 625152
rect 674005 625094 676292 625096
rect 674005 625091 674071 625094
rect 674005 624746 674071 624749
rect 674005 624744 676292 624746
rect 674005 624688 674010 624744
rect 674066 624688 676292 624744
rect 674005 624686 676292 624688
rect 674005 624683 674071 624686
rect 42374 624548 42380 624612
rect 42444 624610 42450 624612
rect 42701 624610 42767 624613
rect 42444 624608 42767 624610
rect 42444 624552 42706 624608
rect 42762 624552 42767 624608
rect 42444 624550 42767 624552
rect 42444 624548 42450 624550
rect 42701 624547 42767 624550
rect 674005 624338 674071 624341
rect 674005 624336 676292 624338
rect 674005 624280 674010 624336
rect 674066 624280 676292 624336
rect 674005 624278 676292 624280
rect 674005 624275 674071 624278
rect 674005 623930 674071 623933
rect 674005 623928 676292 623930
rect 674005 623872 674010 623928
rect 674066 623872 676292 623928
rect 674005 623870 676292 623872
rect 674005 623867 674071 623870
rect 40902 623732 40908 623796
rect 40972 623794 40978 623796
rect 42057 623794 42123 623797
rect 40972 623792 42123 623794
rect 40972 623736 42062 623792
rect 42118 623736 42123 623792
rect 40972 623734 42123 623736
rect 40972 623732 40978 623734
rect 42057 623731 42123 623734
rect 674005 623522 674071 623525
rect 674005 623520 676292 623522
rect 674005 623464 674010 623520
rect 674066 623464 676292 623520
rect 674005 623462 676292 623464
rect 674005 623459 674071 623462
rect 42057 623386 42123 623389
rect 43989 623386 44055 623389
rect 42057 623384 44055 623386
rect 42057 623328 42062 623384
rect 42118 623328 43994 623384
rect 44050 623328 44055 623384
rect 42057 623326 44055 623328
rect 42057 623323 42123 623326
rect 43989 623323 44055 623326
rect 674005 623114 674071 623117
rect 674005 623112 676292 623114
rect 674005 623056 674010 623112
rect 674066 623056 676292 623112
rect 674005 623054 676292 623056
rect 674005 623051 674071 623054
rect 674005 622706 674071 622709
rect 674005 622704 676292 622706
rect 674005 622648 674010 622704
rect 674066 622648 676292 622704
rect 674005 622646 676292 622648
rect 674005 622643 674071 622646
rect 674005 622298 674071 622301
rect 674005 622296 676292 622298
rect 674005 622240 674010 622296
rect 674066 622240 676292 622296
rect 674005 622238 676292 622240
rect 674005 622235 674071 622238
rect 42057 622162 42123 622165
rect 44173 622162 44239 622165
rect 42057 622160 44239 622162
rect 42057 622104 42062 622160
rect 42118 622104 44178 622160
rect 44234 622104 44239 622160
rect 42057 622102 44239 622104
rect 42057 622099 42123 622102
rect 44173 622099 44239 622102
rect 680997 622026 681063 622029
rect 680997 622024 681106 622026
rect 680997 621968 681002 622024
rect 681058 621968 681106 622024
rect 680997 621963 681106 621968
rect 681046 621860 681106 621963
rect 676990 621556 676996 621620
rect 677060 621556 677066 621620
rect 676998 621452 677058 621556
rect 674005 621210 674071 621213
rect 674005 621208 676322 621210
rect 674005 621152 674010 621208
rect 674066 621152 676322 621208
rect 674005 621150 676322 621152
rect 674005 621147 674071 621150
rect 676262 621044 676322 621150
rect 40718 620876 40724 620940
rect 40788 620938 40794 620940
rect 41781 620938 41847 620941
rect 40788 620936 41847 620938
rect 40788 620880 41786 620936
rect 41842 620880 41847 620936
rect 40788 620878 41847 620880
rect 40788 620876 40794 620878
rect 41781 620875 41847 620878
rect 673453 620666 673519 620669
rect 673453 620664 676292 620666
rect 673453 620608 673458 620664
rect 673514 620608 676292 620664
rect 673453 620606 676292 620608
rect 673453 620603 673519 620606
rect 673085 620258 673151 620261
rect 673085 620256 676292 620258
rect 673085 620200 673090 620256
rect 673146 620200 676292 620256
rect 673085 620198 676292 620200
rect 673085 620195 673151 620198
rect 42190 619788 42196 619852
rect 42260 619850 42266 619852
rect 42517 619850 42583 619853
rect 42260 619848 42583 619850
rect 42260 619792 42522 619848
rect 42578 619792 42583 619848
rect 42260 619790 42583 619792
rect 42260 619788 42266 619790
rect 42517 619787 42583 619790
rect 673085 619850 673151 619853
rect 673085 619848 676292 619850
rect 673085 619792 673090 619848
rect 673146 619792 676292 619848
rect 673085 619790 676292 619792
rect 673085 619787 673151 619790
rect 673453 619442 673519 619445
rect 673453 619440 676292 619442
rect 673453 619384 673458 619440
rect 673514 619384 676292 619440
rect 673453 619382 676292 619384
rect 673453 619379 673519 619382
rect 672533 619034 672599 619037
rect 672533 619032 676292 619034
rect 672533 618976 672538 619032
rect 672594 618976 676292 619032
rect 672533 618974 676292 618976
rect 672533 618971 672599 618974
rect 672901 618626 672967 618629
rect 672901 618624 676292 618626
rect 672901 618568 672906 618624
rect 672962 618568 676292 618624
rect 672901 618566 676292 618568
rect 672901 618563 672967 618566
rect 674465 618218 674531 618221
rect 674465 618216 676292 618218
rect 674465 618160 674470 618216
rect 674526 618160 676292 618216
rect 674465 618158 676292 618160
rect 674465 618155 674531 618158
rect 62941 618082 63007 618085
rect 62941 618080 64706 618082
rect 62941 618024 62946 618080
rect 63002 618024 64706 618080
rect 62941 618022 64706 618024
rect 62941 618019 63007 618022
rect 64646 617416 64706 618022
rect 683389 617946 683455 617949
rect 683389 617944 683498 617946
rect 683389 617888 683394 617944
rect 683450 617888 683498 617944
rect 683389 617883 683498 617888
rect 683438 617780 683498 617883
rect 683113 617538 683179 617541
rect 683070 617536 683179 617538
rect 683070 617480 683118 617536
rect 683174 617480 683179 617536
rect 683070 617475 683179 617480
rect 683070 617372 683130 617475
rect 683297 617130 683363 617133
rect 683254 617128 683363 617130
rect 683254 617072 683302 617128
rect 683358 617072 683363 617128
rect 683254 617067 683363 617072
rect 683254 616964 683314 617067
rect 668393 616858 668459 616861
rect 675845 616858 675911 616861
rect 668393 616856 675911 616858
rect 668393 616800 668398 616856
rect 668454 616800 675850 616856
rect 675906 616800 675911 616856
rect 668393 616798 675911 616800
rect 668393 616795 668459 616798
rect 675845 616795 675911 616798
rect 62113 616586 62179 616589
rect 673453 616586 673519 616589
rect 62113 616584 64706 616586
rect 62113 616528 62118 616584
rect 62174 616528 64706 616584
rect 62113 616526 64706 616528
rect 62113 616523 62179 616526
rect 40534 616388 40540 616452
rect 40604 616450 40610 616452
rect 41781 616450 41847 616453
rect 40604 616448 41847 616450
rect 40604 616392 41786 616448
rect 41842 616392 41847 616448
rect 40604 616390 41847 616392
rect 40604 616388 40610 616390
rect 41781 616387 41847 616390
rect 64646 616234 64706 616526
rect 673453 616584 676292 616586
rect 673453 616528 673458 616584
rect 673514 616528 676292 616584
rect 673453 616526 676292 616528
rect 673453 616523 673519 616526
rect 41822 616116 41828 616180
rect 41892 616178 41898 616180
rect 42609 616178 42675 616181
rect 41892 616176 42675 616178
rect 41892 616120 42614 616176
rect 42670 616120 42675 616176
rect 41892 616118 42675 616120
rect 41892 616116 41898 616118
rect 42609 616115 42675 616118
rect 674414 616116 674420 616180
rect 674484 616178 674490 616180
rect 674484 616118 676292 616178
rect 674484 616116 674490 616118
rect 41638 615708 41644 615772
rect 41708 615770 41714 615772
rect 42333 615770 42399 615773
rect 41708 615768 42399 615770
rect 41708 615712 42338 615768
rect 42394 615712 42399 615768
rect 41708 615710 42399 615712
rect 41708 615708 41714 615710
rect 42333 615707 42399 615710
rect 683070 615501 683130 615740
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 41454 615164 41460 615228
rect 41524 615226 41530 615228
rect 42609 615226 42675 615229
rect 41524 615224 42675 615226
rect 41524 615168 42614 615224
rect 42670 615168 42675 615224
rect 41524 615166 42675 615168
rect 41524 615164 41530 615166
rect 42609 615163 42675 615166
rect 62113 614682 62179 614685
rect 64646 614682 64706 615052
rect 673453 614954 673519 614957
rect 673453 614952 676292 614954
rect 673453 614896 673458 614952
rect 673514 614896 676292 614952
rect 673453 614894 676292 614896
rect 673453 614891 673519 614894
rect 62113 614680 64706 614682
rect 62113 614624 62118 614680
rect 62174 614624 64706 614680
rect 62113 614622 64706 614624
rect 62113 614619 62179 614622
rect 42885 613866 42951 613869
rect 44081 613866 44147 613869
rect 42885 613864 44147 613866
rect 42885 613808 42890 613864
rect 42946 613808 44086 613864
rect 44142 613808 44147 613864
rect 42885 613806 44147 613808
rect 42885 613803 42951 613806
rect 44081 613803 44147 613806
rect 61377 613866 61443 613869
rect 64646 613866 64706 613870
rect 61377 613864 64706 613866
rect 61377 613808 61382 613864
rect 61438 613808 64706 613864
rect 61377 613806 64706 613808
rect 61377 613803 61443 613806
rect 62113 612642 62179 612645
rect 64646 612642 64706 612688
rect 62113 612640 64706 612642
rect 62113 612584 62118 612640
rect 62174 612584 64706 612640
rect 62113 612582 64706 612584
rect 62113 612579 62179 612582
rect 43253 612234 43319 612237
rect 43759 612234 43825 612237
rect 43253 612232 43825 612234
rect 43253 612176 43258 612232
rect 43314 612176 43764 612232
rect 43820 612176 43825 612232
rect 43253 612174 43825 612176
rect 43253 612171 43319 612174
rect 43759 612171 43825 612174
rect 44081 612098 44147 612101
rect 45553 612098 45619 612101
rect 44081 612096 45619 612098
rect 44081 612040 44086 612096
rect 44142 612040 45558 612096
rect 45614 612040 45619 612096
rect 44081 612038 45619 612040
rect 44081 612035 44147 612038
rect 45553 612035 45619 612038
rect 62757 612098 62823 612101
rect 62757 612096 64706 612098
rect 62757 612040 62762 612096
rect 62818 612040 64706 612096
rect 62757 612038 64706 612040
rect 62757 612035 62823 612038
rect 43989 611826 44055 611829
rect 47025 611826 47091 611829
rect 43989 611824 47091 611826
rect 43989 611768 43994 611824
rect 44050 611768 47030 611824
rect 47086 611768 47091 611824
rect 43989 611766 47091 611768
rect 43989 611763 44055 611766
rect 47025 611763 47091 611766
rect 44081 611554 44147 611557
rect 47209 611554 47275 611557
rect 44081 611552 47275 611554
rect 44081 611496 44086 611552
rect 44142 611496 47214 611552
rect 47270 611496 47275 611552
rect 64646 611506 64706 612038
rect 44081 611494 47275 611496
rect 44081 611491 44147 611494
rect 47209 611491 47275 611494
rect 673453 611418 673519 611421
rect 675385 611418 675451 611421
rect 673453 611416 675451 611418
rect 673453 611360 673458 611416
rect 673514 611360 675390 611416
rect 675446 611360 675451 611416
rect 673453 611358 675451 611360
rect 673453 611355 673519 611358
rect 675385 611355 675451 611358
rect 675385 608292 675451 608293
rect 675334 608290 675340 608292
rect 675294 608230 675340 608290
rect 675404 608288 675451 608292
rect 675446 608232 675451 608288
rect 675334 608228 675340 608230
rect 675404 608228 675451 608232
rect 675385 608227 675451 608228
rect 669221 608018 669287 608021
rect 675385 608018 675451 608021
rect 669221 608016 675451 608018
rect 669221 607960 669226 608016
rect 669282 607960 675390 608016
rect 675446 607960 675451 608016
rect 669221 607958 675451 607960
rect 669221 607955 669287 607958
rect 675385 607955 675451 607958
rect 672533 606522 672599 606525
rect 675385 606522 675451 606525
rect 672533 606520 675451 606522
rect 672533 606464 672538 606520
rect 672594 606464 675390 606520
rect 675446 606464 675451 606520
rect 672533 606462 675451 606464
rect 672533 606459 672599 606462
rect 675385 606459 675451 606462
rect 675477 604620 675543 604621
rect 675477 604616 675524 604620
rect 675588 604618 675594 604620
rect 675477 604560 675482 604616
rect 675477 604556 675524 604560
rect 675588 604558 675634 604618
rect 675588 604556 675594 604558
rect 675477 604555 675543 604556
rect 673085 604346 673151 604349
rect 675385 604346 675451 604349
rect 673085 604344 675451 604346
rect 673085 604288 673090 604344
rect 673146 604288 675390 604344
rect 675446 604288 675451 604344
rect 673085 604286 675451 604288
rect 673085 604283 673151 604286
rect 675385 604283 675451 604286
rect 672257 603530 672323 603533
rect 675477 603530 675543 603533
rect 672257 603528 675543 603530
rect 672257 603472 672262 603528
rect 672318 603472 675482 603528
rect 675538 603472 675543 603528
rect 672257 603470 675543 603472
rect 672257 603467 672323 603470
rect 675477 603467 675543 603470
rect 673913 602986 673979 602989
rect 675385 602986 675451 602989
rect 673913 602984 675451 602986
rect 673913 602928 673918 602984
rect 673974 602928 675390 602984
rect 675446 602928 675451 602984
rect 673913 602926 675451 602928
rect 673913 602923 673979 602926
rect 675385 602923 675451 602926
rect 35801 601762 35867 601765
rect 35788 601760 35867 601762
rect 35788 601704 35806 601760
rect 35862 601704 35867 601760
rect 35788 601702 35867 601704
rect 35801 601699 35867 601702
rect 38561 601354 38627 601357
rect 38548 601352 38627 601354
rect 38548 601296 38566 601352
rect 38622 601296 38627 601352
rect 38548 601294 38627 601296
rect 38561 601291 38627 601294
rect 39941 600946 40007 600949
rect 39941 600944 40020 600946
rect 39941 600888 39946 600944
rect 40002 600888 40020 600944
rect 39941 600886 40020 600888
rect 39941 600883 40007 600886
rect 44633 600538 44699 600541
rect 41492 600536 44699 600538
rect 41492 600480 44638 600536
rect 44694 600480 44699 600536
rect 41492 600478 44699 600480
rect 44633 600475 44699 600478
rect 670417 600402 670483 600405
rect 675477 600402 675543 600405
rect 670417 600400 675543 600402
rect 670417 600344 670422 600400
rect 670478 600344 675482 600400
rect 675538 600344 675543 600400
rect 670417 600342 675543 600344
rect 670417 600339 670483 600342
rect 675477 600339 675543 600342
rect 44909 600130 44975 600133
rect 41492 600128 44975 600130
rect 41492 600072 44914 600128
rect 44970 600072 44975 600128
rect 41492 600070 44975 600072
rect 44909 600067 44975 600070
rect 673453 600130 673519 600133
rect 674833 600130 674899 600133
rect 673453 600128 674899 600130
rect 673453 600072 673458 600128
rect 673514 600072 674838 600128
rect 674894 600072 674899 600128
rect 673453 600070 674899 600072
rect 673453 600067 673519 600070
rect 674833 600067 674899 600070
rect 675753 599858 675819 599861
rect 675710 599856 675819 599858
rect 675710 599800 675758 599856
rect 675814 599800 675819 599856
rect 675710 599795 675819 599800
rect 44214 599722 44220 599724
rect 41492 599662 44220 599722
rect 44214 599660 44220 599662
rect 44284 599660 44290 599724
rect 672901 599722 672967 599725
rect 675477 599722 675543 599725
rect 672901 599720 675543 599722
rect 672901 599664 672906 599720
rect 672962 599664 675482 599720
rect 675538 599664 675543 599720
rect 672901 599662 675543 599664
rect 672901 599659 672967 599662
rect 675477 599659 675543 599662
rect 674557 599450 674623 599453
rect 675710 599450 675770 599795
rect 674557 599448 675770 599450
rect 674557 599392 674562 599448
rect 674618 599392 675770 599448
rect 674557 599390 675770 599392
rect 674557 599387 674623 599390
rect 43110 599314 43116 599316
rect 41492 599254 43116 599314
rect 43110 599252 43116 599254
rect 43180 599252 43186 599316
rect 675477 599178 675543 599181
rect 675477 599176 675586 599178
rect 675477 599120 675482 599176
rect 675538 599120 675586 599176
rect 675477 599115 675586 599120
rect 673453 599042 673519 599045
rect 675293 599042 675359 599045
rect 673453 599040 675359 599042
rect 673453 598984 673458 599040
rect 673514 598984 675298 599040
rect 675354 598984 675359 599040
rect 673453 598982 675359 598984
rect 673453 598979 673519 598982
rect 675293 598979 675359 598982
rect 45093 598906 45159 598909
rect 41492 598904 45159 598906
rect 41492 598848 45098 598904
rect 45154 598848 45159 598904
rect 41492 598846 45159 598848
rect 675526 598906 675586 599115
rect 676990 598906 676996 598908
rect 675526 598846 676996 598906
rect 45093 598843 45159 598846
rect 676990 598844 676996 598846
rect 677060 598844 677066 598908
rect 674833 598634 674899 598637
rect 675477 598634 675543 598637
rect 675753 598634 675819 598637
rect 674833 598632 675543 598634
rect 674833 598576 674838 598632
rect 674894 598576 675482 598632
rect 675538 598576 675543 598632
rect 674833 598574 675543 598576
rect 674833 598571 674899 598574
rect 675477 598571 675543 598574
rect 675710 598632 675819 598634
rect 675710 598576 675758 598632
rect 675814 598576 675819 598632
rect 675710 598571 675819 598576
rect 45093 598498 45159 598501
rect 41492 598496 45159 598498
rect 41492 598440 45098 598496
rect 45154 598440 45159 598496
rect 41492 598438 45159 598440
rect 45093 598435 45159 598438
rect 674373 598362 674439 598365
rect 675710 598362 675770 598571
rect 674373 598360 675770 598362
rect 45277 598090 45343 598093
rect 41492 598088 45343 598090
rect 41492 598032 45282 598088
rect 45338 598032 45343 598088
rect 41492 598030 45343 598032
rect 45277 598027 45343 598030
rect 649950 597954 650010 598336
rect 674373 598304 674378 598360
rect 674434 598304 675770 598360
rect 674373 598302 675770 598304
rect 674373 598299 674439 598302
rect 651465 597954 651531 597957
rect 649950 597952 651531 597954
rect 649950 597896 651470 597952
rect 651526 597896 651531 597952
rect 649950 597894 651531 597896
rect 651465 597891 651531 597894
rect 42977 597682 43043 597685
rect 41492 597680 43043 597682
rect 41492 597624 42982 597680
rect 43038 597624 43043 597680
rect 41492 597622 43043 597624
rect 42977 597619 43043 597622
rect 674189 597410 674255 597413
rect 675477 597410 675543 597413
rect 674189 597408 675543 597410
rect 674189 597352 674194 597408
rect 674250 597352 675482 597408
rect 675538 597352 675543 597408
rect 674189 597350 675543 597352
rect 674189 597347 674255 597350
rect 675477 597347 675543 597350
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 43161 597004 43227 597005
rect 43110 597002 43116 597004
rect 43070 596942 43116 597002
rect 43180 597000 43227 597004
rect 43222 596944 43227 597000
rect 43110 596940 43116 596942
rect 43180 596940 43227 596944
rect 43161 596939 43227 596940
rect 42609 596866 42675 596869
rect 41492 596864 42675 596866
rect 41492 596808 42614 596864
rect 42670 596808 42675 596864
rect 41492 596806 42675 596808
rect 42609 596803 42675 596806
rect 649950 596730 650010 597154
rect 651465 596730 651531 596733
rect 649950 596728 651531 596730
rect 649950 596672 651470 596728
rect 651526 596672 651531 596728
rect 649950 596670 651531 596672
rect 651465 596667 651531 596670
rect 42190 596458 42196 596460
rect 41492 596398 42196 596458
rect 42190 596396 42196 596398
rect 42260 596396 42266 596460
rect 675293 596322 675359 596325
rect 675518 596322 675524 596324
rect 675293 596320 675524 596322
rect 675293 596264 675298 596320
rect 675354 596264 675524 596320
rect 675293 596262 675524 596264
rect 675293 596259 675359 596262
rect 675518 596260 675524 596262
rect 675588 596260 675594 596324
rect 42333 596050 42399 596053
rect 41492 596048 42399 596050
rect 41492 595992 42338 596048
rect 42394 595992 42399 596048
rect 41492 595990 42399 595992
rect 42333 595987 42399 595990
rect 41689 595778 41755 595781
rect 62941 595778 63007 595781
rect 41689 595776 63007 595778
rect 41689 595720 41694 595776
rect 41750 595720 62946 595776
rect 63002 595720 63007 595776
rect 41689 595718 63007 595720
rect 41689 595715 41755 595718
rect 62941 595715 63007 595718
rect 35390 595407 35450 595612
rect 649950 595506 650010 595972
rect 651465 595506 651531 595509
rect 649950 595504 651531 595506
rect 649950 595448 651470 595504
rect 651526 595448 651531 595504
rect 649950 595446 651531 595448
rect 651465 595443 651531 595446
rect 667565 595506 667631 595509
rect 675385 595506 675451 595509
rect 667565 595504 675451 595506
rect 667565 595448 667570 595504
rect 667626 595448 675390 595504
rect 675446 595448 675451 595504
rect 667565 595446 675451 595448
rect 667565 595443 667631 595446
rect 675385 595443 675451 595446
rect 33041 595404 33107 595407
rect 32998 595402 33107 595404
rect 32998 595346 33046 595402
rect 33102 595346 33107 595402
rect 32998 595341 33107 595346
rect 35390 595402 35499 595407
rect 35390 595346 35438 595402
rect 35494 595346 35499 595402
rect 35390 595344 35499 595346
rect 35433 595341 35499 595344
rect 32998 595204 33058 595341
rect 651649 595234 651715 595237
rect 649950 595232 651715 595234
rect 649950 595176 651654 595232
rect 651710 595176 651715 595232
rect 649950 595174 651715 595176
rect 39297 594826 39363 594829
rect 39284 594824 39363 594826
rect 39284 594768 39302 594824
rect 39358 594768 39363 594824
rect 649950 594790 650010 595174
rect 651649 595171 651715 595174
rect 671337 594826 671403 594829
rect 675477 594826 675543 594829
rect 671337 594824 675543 594826
rect 39284 594766 39363 594768
rect 39297 594763 39363 594766
rect 671337 594768 671342 594824
rect 671398 594768 675482 594824
rect 675538 594768 675543 594824
rect 671337 594766 675543 594768
rect 671337 594763 671403 594766
rect 675477 594763 675543 594766
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 41781 594282 41847 594285
rect 41781 594280 51090 594282
rect 41781 594224 41786 594280
rect 41842 594224 51090 594280
rect 41781 594222 51090 594224
rect 41781 594219 41847 594222
rect 51030 594146 51090 594222
rect 62757 594146 62823 594149
rect 651465 594146 651531 594149
rect 51030 594144 62823 594146
rect 51030 594088 62762 594144
rect 62818 594088 62823 594144
rect 51030 594086 62823 594088
rect 62757 594083 62823 594086
rect 649950 594144 651531 594146
rect 649950 594088 651470 594144
rect 651526 594088 651531 594144
rect 649950 594086 651531 594088
rect 41822 594010 41828 594012
rect 41492 593950 41828 594010
rect 41822 593948 41828 593950
rect 41892 593948 41898 594012
rect 649950 593608 650010 594086
rect 651465 594083 651531 594086
rect 33777 593602 33843 593605
rect 33764 593600 33843 593602
rect 33764 593544 33782 593600
rect 33838 593544 33843 593600
rect 33764 593542 33843 593544
rect 33777 593539 33843 593542
rect 670969 593602 671035 593605
rect 675385 593602 675451 593605
rect 670969 593600 675451 593602
rect 670969 593544 670974 593600
rect 671030 593544 675390 593600
rect 675446 593544 675451 593600
rect 670969 593542 675451 593544
rect 670969 593539 671035 593542
rect 675385 593539 675451 593542
rect 44357 593194 44423 593197
rect 41492 593192 44423 593194
rect 41492 593136 44362 593192
rect 44418 593136 44423 593192
rect 41492 593134 44423 593136
rect 44357 593131 44423 593134
rect 40718 592894 40724 592958
rect 40788 592894 40794 592958
rect 41689 592922 41755 592925
rect 63125 592922 63191 592925
rect 41689 592920 63191 592922
rect 40726 592756 40786 592894
rect 41689 592864 41694 592920
rect 41750 592864 63130 592920
rect 63186 592864 63191 592920
rect 41689 592862 63191 592864
rect 41689 592859 41755 592862
rect 63125 592859 63191 592862
rect 674741 592922 674807 592925
rect 675845 592922 675911 592925
rect 674741 592920 675911 592922
rect 674741 592864 674746 592920
rect 674802 592864 675850 592920
rect 675906 592864 675911 592920
rect 674741 592862 675911 592864
rect 674741 592859 674807 592862
rect 675845 592859 675911 592862
rect 651465 592786 651531 592789
rect 649950 592784 651531 592786
rect 649950 592728 651470 592784
rect 651526 592728 651531 592784
rect 649950 592726 651531 592728
rect 649950 592426 650010 592726
rect 651465 592723 651531 592726
rect 674230 592588 674236 592652
rect 674300 592650 674306 592652
rect 684033 592650 684099 592653
rect 674300 592648 684099 592650
rect 674300 592592 684038 592648
rect 684094 592592 684099 592648
rect 674300 592590 684099 592592
rect 674300 592588 674306 592590
rect 684033 592587 684099 592590
rect 41462 592142 41522 592348
rect 41454 592078 41460 592142
rect 41524 592078 41530 592142
rect 675477 592108 675543 592109
rect 675477 592104 675524 592108
rect 675588 592106 675594 592108
rect 675477 592048 675482 592104
rect 675477 592044 675524 592048
rect 675588 592046 675634 592106
rect 675588 592044 675594 592046
rect 675477 592043 675543 592044
rect 44173 591970 44239 591973
rect 41492 591968 44239 591970
rect 41492 591912 44178 591968
rect 44234 591912 44239 591968
rect 41492 591910 44239 591912
rect 44173 591907 44239 591910
rect 673637 591834 673703 591837
rect 675845 591834 675911 591837
rect 673637 591832 675911 591834
rect 673637 591776 673642 591832
rect 673698 591776 675850 591832
rect 675906 591776 675911 591832
rect 673637 591774 675911 591776
rect 673637 591771 673703 591774
rect 675845 591771 675911 591774
rect 43345 591562 43411 591565
rect 41492 591560 43411 591562
rect 41492 591504 43350 591560
rect 43406 591504 43411 591560
rect 41492 591502 43411 591504
rect 43345 591499 43411 591502
rect 673453 591290 673519 591293
rect 675845 591290 675911 591293
rect 673453 591288 675911 591290
rect 673453 591232 673458 591288
rect 673514 591232 675850 591288
rect 675906 591232 675911 591288
rect 673453 591230 675911 591232
rect 673453 591227 673519 591230
rect 675845 591227 675911 591230
rect 40358 590918 40418 591124
rect 40350 590854 40356 590918
rect 40420 590854 40426 590918
rect 40358 590716 40418 590854
rect 43621 590338 43687 590341
rect 41492 590336 43687 590338
rect 41492 590280 43626 590336
rect 43682 590280 43687 590336
rect 41492 590278 43687 590280
rect 43621 590275 43687 590278
rect 40350 589596 40356 589660
rect 40420 589658 40426 589660
rect 41229 589658 41295 589661
rect 40420 589656 41295 589658
rect 40420 589600 41234 589656
rect 41290 589600 41295 589656
rect 40420 589598 41295 589600
rect 40420 589596 40426 589598
rect 41229 589595 41295 589598
rect 674925 589250 674991 589253
rect 675845 589250 675911 589253
rect 674925 589248 675911 589250
rect 674925 589192 674930 589248
rect 674986 589192 675850 589248
rect 675906 589192 675911 589248
rect 674925 589190 675911 589192
rect 674925 589187 674991 589190
rect 675845 589187 675911 589190
rect 42190 587556 42196 587620
rect 42260 587618 42266 587620
rect 42609 587618 42675 587621
rect 42260 587616 42675 587618
rect 42260 587560 42614 587616
rect 42670 587560 42675 587616
rect 42260 587558 42675 587560
rect 42260 587556 42266 587558
rect 42609 587555 42675 587558
rect 40677 587346 40743 587349
rect 42701 587346 42767 587349
rect 40677 587344 42767 587346
rect 40677 587288 40682 587344
rect 40738 587288 42706 587344
rect 42762 587288 42767 587344
rect 40677 587286 42767 587288
rect 40677 587283 40743 587286
rect 42701 587283 42767 587286
rect 675109 586260 675175 586261
rect 675109 586258 675156 586260
rect 675064 586256 675156 586258
rect 675064 586200 675114 586256
rect 675064 586198 675156 586200
rect 675109 586196 675156 586198
rect 675220 586196 675226 586260
rect 675477 586258 675543 586261
rect 676070 586258 676076 586260
rect 675477 586256 676076 586258
rect 675477 586200 675482 586256
rect 675538 586200 676076 586256
rect 675477 586198 676076 586200
rect 675109 586195 675175 586196
rect 675477 586195 675543 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 40125 585986 40191 585989
rect 40350 585986 40356 585988
rect 40125 585984 40356 585986
rect 40125 585928 40130 585984
rect 40186 585928 40356 585984
rect 40125 585926 40356 585928
rect 40125 585923 40191 585926
rect 40350 585924 40356 585926
rect 40420 585924 40426 585988
rect 41229 585850 41295 585853
rect 42149 585850 42215 585853
rect 41229 585848 42215 585850
rect 41229 585792 41234 585848
rect 41290 585792 42154 585848
rect 42210 585792 42215 585848
rect 41229 585790 42215 585792
rect 41229 585787 41295 585790
rect 42149 585787 42215 585790
rect 39297 585170 39363 585173
rect 41822 585170 41828 585172
rect 39297 585168 41828 585170
rect 39297 585112 39302 585168
rect 39358 585112 41828 585168
rect 39297 585110 41828 585112
rect 39297 585107 39363 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 40585 584626 40651 584629
rect 42701 584626 42767 584629
rect 40585 584624 42767 584626
rect 40585 584568 40590 584624
rect 40646 584568 42706 584624
rect 42762 584568 42767 584624
rect 40585 584566 42767 584568
rect 40585 584563 40651 584566
rect 42701 584563 42767 584566
rect 42149 581908 42215 581909
rect 42149 581906 42196 581908
rect 42104 581904 42196 581906
rect 42104 581848 42154 581904
rect 42104 581846 42196 581848
rect 42149 581844 42196 581846
rect 42260 581844 42266 581908
rect 42149 581843 42215 581844
rect 674005 581634 674071 581637
rect 674649 581634 674715 581637
rect 674005 581632 674715 581634
rect 674005 581576 674010 581632
rect 674066 581576 674654 581632
rect 674710 581576 674715 581632
rect 674005 581574 674715 581576
rect 674005 581571 674071 581574
rect 674649 581571 674715 581574
rect 674005 581090 674071 581093
rect 674005 581088 676292 581090
rect 674005 581032 674010 581088
rect 674066 581032 676292 581088
rect 674005 581030 676292 581032
rect 674005 581027 674071 581030
rect 42149 580682 42215 580685
rect 44633 580682 44699 580685
rect 42149 580680 44699 580682
rect 42149 580624 42154 580680
rect 42210 580624 44638 580680
rect 44694 580624 44699 580680
rect 42149 580622 44699 580624
rect 42149 580619 42215 580622
rect 44633 580619 44699 580622
rect 673637 580682 673703 580685
rect 673637 580680 676292 580682
rect 673637 580624 673642 580680
rect 673698 580624 676292 580680
rect 673637 580622 676292 580624
rect 673637 580619 673703 580622
rect 40350 580212 40356 580276
rect 40420 580274 40426 580276
rect 41781 580274 41847 580277
rect 40420 580272 41847 580274
rect 40420 580216 41786 580272
rect 41842 580216 41847 580272
rect 40420 580214 41847 580216
rect 40420 580212 40426 580214
rect 41781 580211 41847 580214
rect 674005 580274 674071 580277
rect 674005 580272 676292 580274
rect 674005 580216 674010 580272
rect 674066 580216 676292 580272
rect 674005 580214 676292 580216
rect 674005 580211 674071 580214
rect 674005 579866 674071 579869
rect 674005 579864 676292 579866
rect 674005 579808 674010 579864
rect 674066 579808 676292 579864
rect 674005 579806 676292 579808
rect 674005 579803 674071 579806
rect 673453 579458 673519 579461
rect 673453 579456 676292 579458
rect 673453 579400 673458 579456
rect 673514 579400 676292 579456
rect 673453 579398 676292 579400
rect 673453 579395 673519 579398
rect 674005 579050 674071 579053
rect 674005 579048 676292 579050
rect 674005 578992 674010 579048
rect 674066 578992 676292 579048
rect 674005 578990 676292 578992
rect 674005 578987 674071 578990
rect 42057 578778 42123 578781
rect 44173 578778 44239 578781
rect 42057 578776 44239 578778
rect 42057 578720 42062 578776
rect 42118 578720 44178 578776
rect 44234 578720 44239 578776
rect 42057 578718 44239 578720
rect 42057 578715 42123 578718
rect 44173 578715 44239 578718
rect 674005 578642 674071 578645
rect 674005 578640 676292 578642
rect 674005 578584 674010 578640
rect 674066 578584 676292 578640
rect 674005 578582 676292 578584
rect 674005 578579 674071 578582
rect 42241 578506 42307 578509
rect 45553 578506 45619 578509
rect 42241 578504 45619 578506
rect 42241 578448 42246 578504
rect 42302 578448 45558 578504
rect 45614 578448 45619 578504
rect 42241 578446 45619 578448
rect 42241 578443 42307 578446
rect 45553 578443 45619 578446
rect 673637 578234 673703 578237
rect 673637 578232 676292 578234
rect 673637 578176 673642 578232
rect 673698 578176 676292 578232
rect 673637 578174 676292 578176
rect 673637 578171 673703 578174
rect 42057 578098 42123 578101
rect 44357 578098 44423 578101
rect 42057 578096 44423 578098
rect 42057 578040 42062 578096
rect 42118 578040 44362 578096
rect 44418 578040 44423 578096
rect 42057 578038 44423 578040
rect 42057 578035 42123 578038
rect 44357 578035 44423 578038
rect 40902 577764 40908 577828
rect 40972 577826 40978 577828
rect 41781 577826 41847 577829
rect 40972 577824 41847 577826
rect 40972 577768 41786 577824
rect 41842 577768 41847 577824
rect 40972 577766 41847 577768
rect 40972 577764 40978 577766
rect 41781 577763 41847 577766
rect 675845 577826 675911 577829
rect 675845 577824 676292 577826
rect 675845 577768 675850 577824
rect 675906 577768 676292 577824
rect 675845 577766 676292 577768
rect 675845 577763 675911 577766
rect 674005 577418 674071 577421
rect 674005 577416 676292 577418
rect 674005 577360 674010 577416
rect 674066 577360 676292 577416
rect 674005 577358 676292 577360
rect 674005 577355 674071 577358
rect 674005 577010 674071 577013
rect 674005 577008 676292 577010
rect 674005 576952 674010 577008
rect 674066 576952 676292 577008
rect 674005 576950 676292 576952
rect 674005 576947 674071 576950
rect 673453 576738 673519 576741
rect 675845 576738 675911 576741
rect 673453 576736 675911 576738
rect 673453 576680 673458 576736
rect 673514 576680 675850 576736
rect 675906 576680 675911 576736
rect 673453 576678 675911 576680
rect 673453 576675 673519 576678
rect 675845 576675 675911 576678
rect 672717 576466 672783 576469
rect 676262 576466 676322 576572
rect 672717 576464 676322 576466
rect 672717 576408 672722 576464
rect 672778 576408 676322 576464
rect 672717 576406 676322 576408
rect 678237 576466 678303 576469
rect 678237 576464 678346 576466
rect 678237 576408 678242 576464
rect 678298 576408 678346 576464
rect 672717 576403 672783 576406
rect 678237 576403 678346 576408
rect 678286 576164 678346 576403
rect 674005 575786 674071 575789
rect 674005 575784 676292 575786
rect 674005 575728 674010 575784
rect 674066 575728 676292 575784
rect 674005 575726 676292 575728
rect 674005 575723 674071 575726
rect 40534 575588 40540 575652
rect 40604 575650 40610 575652
rect 42241 575650 42307 575653
rect 684033 575650 684099 575653
rect 40604 575648 42307 575650
rect 40604 575592 42246 575648
rect 42302 575592 42307 575648
rect 40604 575590 42307 575592
rect 40604 575588 40610 575590
rect 42241 575587 42307 575590
rect 683990 575648 684099 575650
rect 683990 575592 684038 575648
rect 684094 575592 684099 575648
rect 683990 575587 684099 575592
rect 683990 575348 684050 575587
rect 676990 575180 676996 575244
rect 677060 575180 677066 575244
rect 676998 574940 677058 575180
rect 62113 574834 62179 574837
rect 62113 574832 64706 574834
rect 62113 574776 62118 574832
rect 62174 574776 64706 574832
rect 62113 574774 64706 574776
rect 62113 574771 62179 574774
rect 40718 574636 40724 574700
rect 40788 574698 40794 574700
rect 41781 574698 41847 574701
rect 40788 574696 41847 574698
rect 40788 574640 41786 574696
rect 41842 574640 41847 574696
rect 40788 574638 41847 574640
rect 40788 574636 40794 574638
rect 41781 574635 41847 574638
rect 64646 574194 64706 574774
rect 673637 574562 673703 574565
rect 673637 574560 676292 574562
rect 673637 574504 673642 574560
rect 673698 574504 676292 574560
rect 673637 574502 676292 574504
rect 673637 574499 673703 574502
rect 674005 574154 674071 574157
rect 674005 574152 676292 574154
rect 674005 574096 674010 574152
rect 674066 574096 676292 574152
rect 674005 574094 676292 574096
rect 674005 574091 674071 574094
rect 684217 574018 684283 574021
rect 684174 574016 684283 574018
rect 684174 573960 684222 574016
rect 684278 573960 684283 574016
rect 684174 573955 684283 573960
rect 684174 573716 684234 573955
rect 62113 573610 62179 573613
rect 62113 573608 64706 573610
rect 62113 573552 62118 573608
rect 62174 573552 64706 573608
rect 62113 573550 64706 573552
rect 62113 573547 62179 573550
rect 64646 573012 64706 573550
rect 676806 573548 676812 573612
rect 676876 573548 676882 573612
rect 676814 573308 676874 573548
rect 674005 572930 674071 572933
rect 674005 572928 676292 572930
rect 674005 572872 674010 572928
rect 674066 572872 676292 572928
rect 674005 572870 676292 572872
rect 674005 572867 674071 572870
rect 41454 572732 41460 572796
rect 41524 572794 41530 572796
rect 42609 572794 42675 572797
rect 41524 572792 42675 572794
rect 41524 572736 42614 572792
rect 42670 572736 42675 572792
rect 41524 572734 42675 572736
rect 41524 572732 41530 572734
rect 42609 572731 42675 572734
rect 673637 572522 673703 572525
rect 673637 572520 676292 572522
rect 673637 572464 673642 572520
rect 673698 572464 676292 572520
rect 673637 572462 676292 572464
rect 673637 572459 673703 572462
rect 674005 572114 674071 572117
rect 674005 572112 676292 572114
rect 674005 572056 674010 572112
rect 674066 572056 676292 572112
rect 674005 572054 676292 572056
rect 674005 572051 674071 572054
rect 683389 571978 683455 571981
rect 683389 571976 683498 571978
rect 683389 571920 683394 571976
rect 683450 571920 683498 571976
rect 683389 571915 683498 571920
rect 41638 571508 41644 571572
rect 41708 571570 41714 571572
rect 42057 571570 42123 571573
rect 41708 571568 42123 571570
rect 41708 571512 42062 571568
rect 42118 571512 42123 571568
rect 41708 571510 42123 571512
rect 41708 571508 41714 571510
rect 42057 571507 42123 571510
rect 42425 571434 42491 571437
rect 64646 571434 64706 571830
rect 683438 571676 683498 571915
rect 42425 571432 64706 571434
rect 42425 571376 42430 571432
rect 42486 571376 64706 571432
rect 42425 571374 64706 571376
rect 674649 571434 674715 571437
rect 674649 571432 676322 571434
rect 674649 571376 674654 571432
rect 674710 571376 676322 571432
rect 674649 571374 676322 571376
rect 42425 571371 42491 571374
rect 674649 571371 674715 571374
rect 676262 571268 676322 571374
rect 62941 571162 63007 571165
rect 62941 571160 64706 571162
rect 62941 571104 62946 571160
rect 63002 571104 64706 571160
rect 62941 571102 64706 571104
rect 62941 571099 63007 571102
rect 64646 570648 64706 571102
rect 671470 570692 671476 570756
rect 671540 570754 671546 570756
rect 676262 570754 676322 570860
rect 683113 570754 683179 570757
rect 671540 570694 676322 570754
rect 683070 570752 683179 570754
rect 683070 570696 683118 570752
rect 683174 570696 683179 570752
rect 671540 570692 671546 570694
rect 683070 570691 683179 570696
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 683070 570044 683130 570691
rect 63125 569938 63191 569941
rect 63125 569936 64706 569938
rect 63125 569880 63130 569936
rect 63186 569880 64706 569936
rect 63125 569878 64706 569880
rect 63125 569875 63191 569878
rect 64646 569466 64706 569878
rect 676262 569533 676322 569636
rect 676213 569528 676322 569533
rect 676213 569472 676218 569528
rect 676274 569472 676322 569528
rect 676213 569470 676322 569472
rect 676213 569467 676279 569470
rect 62757 568578 62823 568581
rect 62757 568576 64706 568578
rect 62757 568520 62762 568576
rect 62818 568520 64706 568576
rect 62757 568518 64706 568520
rect 62757 568515 62823 568518
rect 64646 568284 64706 568518
rect 674005 565858 674071 565861
rect 675385 565858 675451 565861
rect 674005 565856 675451 565858
rect 674005 565800 674010 565856
rect 674066 565800 675390 565856
rect 675446 565800 675451 565856
rect 674005 565798 675451 565800
rect 674005 565795 674071 565798
rect 675385 565795 675451 565798
rect 673862 565524 673868 565588
rect 673932 565586 673938 565588
rect 676213 565586 676279 565589
rect 673932 565584 676279 565586
rect 673932 565528 676218 565584
rect 676274 565528 676279 565584
rect 673932 565526 676279 565528
rect 673932 565524 673938 565526
rect 676213 565523 676279 565526
rect 675753 562730 675819 562733
rect 676438 562730 676444 562732
rect 675753 562728 676444 562730
rect 675753 562672 675758 562728
rect 675814 562672 676444 562728
rect 675753 562670 676444 562672
rect 675753 562667 675819 562670
rect 676438 562668 676444 562670
rect 676508 562668 676514 562732
rect 669037 562322 669103 562325
rect 675109 562322 675175 562325
rect 669037 562320 675175 562322
rect 669037 562264 669042 562320
rect 669098 562264 675114 562320
rect 675170 562264 675175 562320
rect 669037 562262 675175 562264
rect 669037 562259 669103 562262
rect 675109 562259 675175 562262
rect 675385 561916 675451 561917
rect 675334 561914 675340 561916
rect 675294 561854 675340 561914
rect 675404 561912 675451 561916
rect 675446 561856 675451 561912
rect 675334 561852 675340 561854
rect 675404 561852 675451 561856
rect 675385 561851 675451 561852
rect 41086 558724 41092 558788
rect 41156 558786 41162 558788
rect 44909 558786 44975 558789
rect 41156 558784 44975 558786
rect 41156 558728 44914 558784
rect 44970 558728 44975 558784
rect 41156 558726 44975 558728
rect 41156 558724 41162 558726
rect 44909 558723 44975 558726
rect 41492 558454 51090 558514
rect 42333 558106 42399 558109
rect 41492 558104 42399 558106
rect 41492 558048 42338 558104
rect 42394 558048 42399 558104
rect 41492 558046 42399 558048
rect 42333 558043 42399 558046
rect 41492 557638 48330 557698
rect 41086 557488 41092 557552
rect 41156 557488 41162 557552
rect 41094 557260 41154 557488
rect 48270 557290 48330 557638
rect 51030 557562 51090 558454
rect 673637 558106 673703 558109
rect 675385 558106 675451 558109
rect 673637 558104 675451 558106
rect 673637 558048 673642 558104
rect 673698 558048 675390 558104
rect 675446 558048 675451 558104
rect 673637 558046 675451 558048
rect 673637 558043 673703 558046
rect 675385 558043 675451 558046
rect 61377 557562 61443 557565
rect 51030 557560 61443 557562
rect 51030 557504 61382 557560
rect 61438 557504 61443 557560
rect 51030 557502 61443 557504
rect 61377 557499 61443 557502
rect 673269 557562 673335 557565
rect 675385 557562 675451 557565
rect 673269 557560 675451 557562
rect 673269 557504 673274 557560
rect 673330 557504 675390 557560
rect 675446 557504 675451 557560
rect 673269 557502 675451 557504
rect 673269 557499 673335 557502
rect 675385 557499 675451 557502
rect 48270 557230 51090 557290
rect 44541 556882 44607 556885
rect 41492 556880 44607 556882
rect 41492 556824 44546 556880
rect 44602 556824 44607 556880
rect 41492 556822 44607 556824
rect 44541 556819 44607 556822
rect 51030 556746 51090 557230
rect 63401 556746 63467 556749
rect 51030 556744 63467 556746
rect 51030 556688 63406 556744
rect 63462 556688 63467 556744
rect 51030 556686 63467 556688
rect 63401 556683 63467 556686
rect 43069 556474 43135 556477
rect 41492 556472 43135 556474
rect 41492 556416 43074 556472
rect 43130 556416 43135 556472
rect 41492 556414 43135 556416
rect 43069 556411 43135 556414
rect 44265 556066 44331 556069
rect 41492 556064 44331 556066
rect 41492 556008 44270 556064
rect 44326 556008 44331 556064
rect 41492 556006 44331 556008
rect 44265 556003 44331 556006
rect 45093 555658 45159 555661
rect 41492 555656 45159 555658
rect 41492 555600 45098 555656
rect 45154 555600 45159 555656
rect 41492 555598 45159 555600
rect 45093 555595 45159 555598
rect 673913 555522 673979 555525
rect 675109 555522 675175 555525
rect 673913 555520 675175 555522
rect 673913 555464 673918 555520
rect 673974 555464 675114 555520
rect 675170 555464 675175 555520
rect 673913 555462 675175 555464
rect 673913 555459 673979 555462
rect 675109 555459 675175 555462
rect 45645 555250 45711 555253
rect 41492 555248 45711 555250
rect 41492 555192 45650 555248
rect 45706 555192 45711 555248
rect 41492 555190 45711 555192
rect 45645 555187 45711 555190
rect 668393 555250 668459 555253
rect 675385 555250 675451 555253
rect 668393 555248 675451 555250
rect 668393 555192 668398 555248
rect 668454 555192 675390 555248
rect 675446 555192 675451 555248
rect 668393 555190 675451 555192
rect 668393 555187 668459 555190
rect 675385 555187 675451 555190
rect 42793 554842 42859 554845
rect 41492 554840 42859 554842
rect 41492 554784 42798 554840
rect 42854 554784 42859 554840
rect 41492 554782 42859 554784
rect 42793 554779 42859 554782
rect 674005 554706 674071 554709
rect 675109 554706 675175 554709
rect 674005 554704 675175 554706
rect 674005 554648 674010 554704
rect 674066 554648 675114 554704
rect 675170 554648 675175 554704
rect 674005 554646 675175 554648
rect 674005 554643 674071 554646
rect 675109 554643 675175 554646
rect 45829 554434 45895 554437
rect 41492 554432 45895 554434
rect 41492 554376 45834 554432
rect 45890 554376 45895 554432
rect 41492 554374 45895 554376
rect 45829 554371 45895 554374
rect 41822 554026 41828 554028
rect 41492 553966 41828 554026
rect 41822 553964 41828 553966
rect 41892 553964 41898 554028
rect 39990 553413 40050 553588
rect 649950 553482 650010 553914
rect 675753 553890 675819 553893
rect 676806 553890 676812 553892
rect 675753 553888 676812 553890
rect 675753 553832 675758 553888
rect 675814 553832 676812 553888
rect 675753 553830 676812 553832
rect 675753 553827 675819 553830
rect 676806 553828 676812 553830
rect 676876 553828 676882 553892
rect 651465 553482 651531 553485
rect 649950 553480 651531 553482
rect 649950 553424 651470 553480
rect 651526 553424 651531 553480
rect 649950 553422 651531 553424
rect 651465 553419 651531 553422
rect 671981 553482 672047 553485
rect 675385 553482 675451 553485
rect 671981 553480 675451 553482
rect 671981 553424 671986 553480
rect 672042 553424 675390 553480
rect 675446 553424 675451 553480
rect 671981 553422 675451 553424
rect 671981 553419 672047 553422
rect 675385 553419 675451 553422
rect 39990 553408 40099 553413
rect 40953 553410 41019 553413
rect 39990 553352 40038 553408
rect 40094 553352 40099 553408
rect 39990 553350 40099 553352
rect 40033 553347 40099 553350
rect 40910 553408 41019 553410
rect 40910 553352 40958 553408
rect 41014 553352 41019 553408
rect 40910 553347 41019 553352
rect 40910 553180 40970 553347
rect 674097 552938 674163 552941
rect 675201 552938 675267 552941
rect 674097 552936 675267 552938
rect 674097 552880 674102 552936
rect 674158 552880 675206 552936
rect 675262 552880 675267 552936
rect 674097 552878 675267 552880
rect 674097 552875 674163 552878
rect 675201 552875 675267 552878
rect 41822 552802 41828 552804
rect 41492 552742 41828 552802
rect 41822 552740 41828 552742
rect 41892 552740 41898 552804
rect 42333 552666 42399 552669
rect 62941 552666 63007 552669
rect 42333 552664 63007 552666
rect 42333 552608 42338 552664
rect 42394 552608 62946 552664
rect 63002 552608 63007 552664
rect 42333 552606 63007 552608
rect 42333 552603 42399 552606
rect 62941 552603 63007 552606
rect 42977 552394 43043 552397
rect 41492 552392 43043 552394
rect 41492 552336 42982 552392
rect 43038 552336 43043 552392
rect 41492 552334 43043 552336
rect 649950 552394 650010 552732
rect 651465 552394 651531 552397
rect 649950 552392 651531 552394
rect 649950 552336 651470 552392
rect 651526 552336 651531 552392
rect 649950 552334 651531 552336
rect 42977 552331 43043 552334
rect 651465 552331 651531 552334
rect 675753 552122 675819 552125
rect 676990 552122 676996 552124
rect 675753 552120 676996 552122
rect 675753 552064 675758 552120
rect 675814 552064 676996 552120
rect 675753 552062 676996 552064
rect 675753 552059 675819 552062
rect 676990 552060 676996 552062
rect 677060 552060 677066 552124
rect 34421 551986 34487 551989
rect 34421 551984 34500 551986
rect 34421 551928 34426 551984
rect 34482 551928 34500 551984
rect 34421 551926 34500 551928
rect 34421 551923 34487 551926
rect 45185 551578 45251 551581
rect 41492 551576 45251 551578
rect 41492 551520 45190 551576
rect 45246 551520 45251 551576
rect 41492 551518 45251 551520
rect 45185 551515 45251 551518
rect 42793 551170 42859 551173
rect 41492 551168 42859 551170
rect 41492 551112 42798 551168
rect 42854 551112 42859 551168
rect 41492 551110 42859 551112
rect 42793 551107 42859 551110
rect 649950 551034 650010 551550
rect 652017 551034 652083 551037
rect 649950 551032 652083 551034
rect 649950 550976 652022 551032
rect 652078 550976 652083 551032
rect 649950 550974 652083 550976
rect 652017 550971 652083 550974
rect 45369 550762 45435 550765
rect 41492 550760 45435 550762
rect 41492 550704 45374 550760
rect 45430 550704 45435 550760
rect 41492 550702 45435 550704
rect 45369 550699 45435 550702
rect 41873 550354 41939 550357
rect 41492 550352 41939 550354
rect 41492 550296 41878 550352
rect 41934 550296 41939 550352
rect 41492 550294 41939 550296
rect 649950 550354 650010 550368
rect 651373 550354 651439 550357
rect 649950 550352 651439 550354
rect 649950 550296 651378 550352
rect 651434 550296 651439 550352
rect 649950 550294 651439 550296
rect 41873 550291 41939 550294
rect 651373 550291 651439 550294
rect 42057 549946 42123 549949
rect 41492 549944 42123 549946
rect 41492 549888 42062 549944
rect 42118 549888 42123 549944
rect 41492 549886 42123 549888
rect 42057 549883 42123 549886
rect 674833 549810 674899 549813
rect 675385 549810 675451 549813
rect 674833 549808 675451 549810
rect 674833 549752 674838 549808
rect 674894 549752 675390 549808
rect 675446 549752 675451 549808
rect 674833 549750 675451 549752
rect 674833 549747 674899 549750
rect 675385 549747 675451 549750
rect 43161 549538 43227 549541
rect 41492 549536 43227 549538
rect 41492 549480 43166 549536
rect 43222 549480 43227 549536
rect 41492 549478 43227 549480
rect 43161 549475 43227 549478
rect 673453 549266 673519 549269
rect 675385 549266 675451 549269
rect 673453 549264 675451 549266
rect 673453 549208 673458 549264
rect 673514 549208 675390 549264
rect 675446 549208 675451 549264
rect 673453 549206 675451 549208
rect 673453 549203 673519 549206
rect 675385 549203 675451 549206
rect 45001 549130 45067 549133
rect 41492 549128 45067 549130
rect 41492 549072 45006 549128
rect 45062 549072 45067 549128
rect 41492 549070 45067 549072
rect 649950 549130 650010 549186
rect 651465 549130 651531 549133
rect 649950 549128 651531 549130
rect 649950 549072 651470 549128
rect 651526 549072 651531 549128
rect 649950 549070 651531 549072
rect 45001 549067 45067 549070
rect 651465 549067 651531 549070
rect 44725 548722 44791 548725
rect 41492 548720 44791 548722
rect 41492 548664 44730 548720
rect 44786 548664 44791 548720
rect 41492 548662 44791 548664
rect 44725 548659 44791 548662
rect 651465 548450 651531 548453
rect 649950 548448 651531 548450
rect 649950 548392 651470 548448
rect 651526 548392 651531 548448
rect 649950 548390 651531 548392
rect 43805 548314 43871 548317
rect 41492 548312 43871 548314
rect 41492 548256 43810 548312
rect 43866 548256 43871 548312
rect 41492 548254 43871 548256
rect 43805 548251 43871 548254
rect 649950 548004 650010 548390
rect 651465 548387 651531 548390
rect 28766 547498 28826 547890
rect 675477 547634 675543 547637
rect 676029 547634 676095 547637
rect 675477 547632 676095 547634
rect 675477 547576 675482 547632
rect 675538 547576 676034 547632
rect 676090 547576 676095 547632
rect 675477 547574 676095 547576
rect 675477 547571 675543 547574
rect 676029 547571 676095 547574
rect 676438 547572 676444 547636
rect 676508 547634 676514 547636
rect 677409 547634 677475 547637
rect 676508 547632 677475 547634
rect 676508 547576 677414 547632
rect 677470 547576 677475 547632
rect 676508 547574 677475 547576
rect 676508 547572 676514 547574
rect 677409 547571 677475 547574
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 675886 547300 675892 547364
rect 675956 547362 675962 547364
rect 678237 547362 678303 547365
rect 675956 547360 678303 547362
rect 675956 547304 678242 547360
rect 678298 547304 678303 547360
rect 675956 547302 678303 547304
rect 675956 547300 675962 547302
rect 678237 547299 678303 547302
rect 43989 547090 44055 547093
rect 41492 547088 44055 547090
rect 41492 547032 43994 547088
rect 44050 547032 44055 547088
rect 41492 547030 44055 547032
rect 43989 547027 44055 547030
rect 676070 547028 676076 547092
rect 676140 547090 676146 547092
rect 680997 547090 681063 547093
rect 676140 547088 681063 547090
rect 676140 547032 681002 547088
rect 681058 547032 681063 547088
rect 676140 547030 681063 547032
rect 676140 547028 676146 547030
rect 680997 547027 681063 547030
rect 41321 546410 41387 546413
rect 41638 546410 41644 546412
rect 41321 546408 41644 546410
rect 41321 546352 41326 546408
rect 41382 546352 41644 546408
rect 41321 546350 41644 546352
rect 41321 546347 41387 546350
rect 41638 546348 41644 546350
rect 41708 546348 41714 546412
rect 40718 545668 40724 545732
rect 40788 545730 40794 545732
rect 41873 545730 41939 545733
rect 40788 545728 41939 545730
rect 40788 545672 41878 545728
rect 41934 545672 41939 545728
rect 40788 545670 41939 545672
rect 40788 545668 40794 545670
rect 41873 545667 41939 545670
rect 40534 545396 40540 545460
rect 40604 545458 40610 545460
rect 42057 545458 42123 545461
rect 40604 545456 42123 545458
rect 40604 545400 42062 545456
rect 42118 545400 42123 545456
rect 40604 545398 42123 545400
rect 40604 545396 40610 545398
rect 42057 545395 42123 545398
rect 675293 544508 675359 544509
rect 675293 544506 675340 544508
rect 675248 544504 675340 544506
rect 675248 544448 675298 544504
rect 675248 544446 675340 544448
rect 675293 544444 675340 544446
rect 675404 544444 675410 544508
rect 675293 544443 675359 544444
rect 41321 541376 41387 541381
rect 41321 541320 41326 541376
rect 41382 541320 41387 541376
rect 41321 541315 41387 541320
rect 41324 540698 41384 541315
rect 41781 540698 41847 540701
rect 41324 540696 41847 540698
rect 41324 540640 41786 540696
rect 41842 540640 41847 540696
rect 41324 540638 41847 540640
rect 41781 540635 41847 540638
rect 42517 539610 42583 539613
rect 59997 539610 60063 539613
rect 42517 539608 60063 539610
rect 42517 539552 42522 539608
rect 42578 539552 60002 539608
rect 60058 539552 60063 539608
rect 42517 539550 60063 539552
rect 42517 539547 42583 539550
rect 59997 539547 60063 539550
rect 42609 538114 42675 538117
rect 45001 538114 45067 538117
rect 42609 538112 45067 538114
rect 42609 538056 42614 538112
rect 42670 538056 45006 538112
rect 45062 538056 45067 538112
rect 42609 538054 45067 538056
rect 42609 538051 42675 538054
rect 45001 538051 45067 538054
rect 40534 537372 40540 537436
rect 40604 537434 40610 537436
rect 42425 537434 42491 537437
rect 40604 537432 42491 537434
rect 40604 537376 42430 537432
rect 42486 537376 42491 537432
rect 40604 537374 42491 537376
rect 40604 537372 40610 537374
rect 42425 537371 42491 537374
rect 674465 537162 674531 537165
rect 675845 537162 675911 537165
rect 674465 537160 675911 537162
rect 674465 537104 674470 537160
rect 674526 537104 675850 537160
rect 675906 537104 675911 537160
rect 674465 537102 675911 537104
rect 674465 537099 674531 537102
rect 675845 537099 675911 537102
rect 40718 536964 40724 537028
rect 40788 537026 40794 537028
rect 41781 537026 41847 537029
rect 40788 537024 41847 537026
rect 40788 536968 41786 537024
rect 41842 536968 41847 537024
rect 40788 536966 41847 536968
rect 40788 536964 40794 536966
rect 41781 536963 41847 536966
rect 44725 536890 44791 536893
rect 42198 536888 44791 536890
rect 42198 536832 44730 536888
rect 44786 536832 44791 536888
rect 42198 536830 44791 536832
rect 42198 536485 42258 536830
rect 44725 536827 44791 536830
rect 42198 536480 42307 536485
rect 42198 536424 42246 536480
rect 42302 536424 42307 536480
rect 42198 536422 42307 536424
rect 42241 536419 42307 536422
rect 673821 536074 673887 536077
rect 676262 536074 676322 536112
rect 673821 536072 676322 536074
rect 673821 536016 673826 536072
rect 673882 536016 676322 536072
rect 673821 536014 676322 536016
rect 673821 536011 673887 536014
rect 42057 535666 42123 535669
rect 44725 535666 44791 535669
rect 42057 535664 44791 535666
rect 42057 535608 42062 535664
rect 42118 535608 44730 535664
rect 44786 535608 44791 535664
rect 42057 535606 44791 535608
rect 42057 535603 42123 535606
rect 44725 535603 44791 535606
rect 674005 535666 674071 535669
rect 676262 535666 676322 535704
rect 674005 535664 676322 535666
rect 674005 535608 674010 535664
rect 674066 535608 676322 535664
rect 674005 535606 676322 535608
rect 674005 535603 674071 535606
rect 673453 535258 673519 535261
rect 676262 535258 676322 535296
rect 673453 535256 676322 535258
rect 673453 535200 673458 535256
rect 673514 535200 676322 535256
rect 673453 535198 676322 535200
rect 673453 535195 673519 535198
rect 674005 534850 674071 534853
rect 676262 534850 676322 534888
rect 674005 534848 676322 534850
rect 674005 534792 674010 534848
rect 674066 534792 676322 534848
rect 674005 534790 676322 534792
rect 674005 534787 674071 534790
rect 673821 534442 673887 534445
rect 676262 534442 676322 534480
rect 673821 534440 676322 534442
rect 673821 534384 673826 534440
rect 673882 534384 676322 534440
rect 673821 534382 676322 534384
rect 673821 534379 673887 534382
rect 674005 534170 674071 534173
rect 674005 534168 676322 534170
rect 674005 534112 674010 534168
rect 674066 534112 676322 534168
rect 674005 534110 676322 534112
rect 674005 534107 674071 534110
rect 676262 534072 676322 534110
rect 674005 533626 674071 533629
rect 676262 533626 676322 533664
rect 674005 533624 676322 533626
rect 674005 533568 674010 533624
rect 674066 533568 676322 533624
rect 674005 533566 676322 533568
rect 674005 533563 674071 533566
rect 674005 533354 674071 533357
rect 674005 533352 676322 533354
rect 674005 533296 674010 533352
rect 674066 533296 676322 533352
rect 674005 533294 676322 533296
rect 674005 533291 674071 533294
rect 676262 533256 676322 533294
rect 42701 532810 42767 532813
rect 45369 532810 45435 532813
rect 42701 532808 45435 532810
rect 42701 532752 42706 532808
rect 42762 532752 45374 532808
rect 45430 532752 45435 532808
rect 42701 532750 45435 532752
rect 42701 532747 42767 532750
rect 45369 532747 45435 532750
rect 674005 532810 674071 532813
rect 676262 532810 676322 532848
rect 674005 532808 676322 532810
rect 674005 532752 674010 532808
rect 674066 532752 676322 532808
rect 674005 532750 676322 532752
rect 674005 532747 674071 532750
rect 674005 532538 674071 532541
rect 674005 532536 676322 532538
rect 674005 532480 674010 532536
rect 674066 532480 676322 532536
rect 674005 532478 676322 532480
rect 674005 532475 674071 532478
rect 676262 532440 676322 532478
rect 674005 531994 674071 531997
rect 676262 531994 676322 532032
rect 674005 531992 676322 531994
rect 674005 531936 674010 531992
rect 674066 531936 676322 531992
rect 674005 531934 676322 531936
rect 674005 531931 674071 531934
rect 674005 531722 674071 531725
rect 674005 531720 676322 531722
rect 674005 531664 674010 531720
rect 674066 531664 676322 531720
rect 674005 531662 676322 531664
rect 674005 531659 674071 531662
rect 676262 531624 676322 531662
rect 62113 531314 62179 531317
rect 62113 531312 64154 531314
rect 62113 531256 62118 531312
rect 62174 531256 64154 531312
rect 62113 531254 64154 531256
rect 62113 531251 62179 531254
rect 64094 531202 64154 531254
rect 64094 531142 64676 531202
rect 674005 531178 674071 531181
rect 676262 531178 676322 531216
rect 674005 531176 676322 531178
rect 674005 531120 674010 531176
rect 674066 531120 676322 531176
rect 674005 531118 676322 531120
rect 674005 531115 674071 531118
rect 680997 531042 681063 531045
rect 680997 531040 681106 531042
rect 680997 530984 681002 531040
rect 681058 530984 681106 531040
rect 680997 530979 681106 530984
rect 681046 530808 681106 530979
rect 41454 530708 41460 530772
rect 41524 530770 41530 530772
rect 42609 530770 42675 530773
rect 41524 530768 42675 530770
rect 41524 530712 42614 530768
rect 42670 530712 42675 530768
rect 41524 530710 42675 530712
rect 41524 530708 41530 530710
rect 42609 530707 42675 530710
rect 62113 530634 62179 530637
rect 678237 530634 678303 530637
rect 62113 530632 64706 530634
rect 62113 530576 62118 530632
rect 62174 530576 64706 530632
rect 62113 530574 64706 530576
rect 62113 530571 62179 530574
rect 64646 529990 64706 530574
rect 678237 530632 678346 530634
rect 678237 530576 678242 530632
rect 678298 530576 678346 530632
rect 678237 530571 678346 530576
rect 678286 530400 678346 530571
rect 673821 530090 673887 530093
rect 673821 530088 676322 530090
rect 673821 530032 673826 530088
rect 673882 530032 676322 530088
rect 673821 530030 676322 530032
rect 673821 530027 673887 530030
rect 676262 529992 676322 530030
rect 674005 529682 674071 529685
rect 674005 529680 676322 529682
rect 674005 529624 674010 529680
rect 674066 529624 676322 529680
rect 674005 529622 676322 529624
rect 674005 529619 674071 529622
rect 676262 529584 676322 529622
rect 41638 529484 41644 529548
rect 41708 529546 41714 529548
rect 42425 529546 42491 529549
rect 41708 529544 42491 529546
rect 41708 529488 42430 529544
rect 42486 529488 42491 529544
rect 41708 529486 42491 529488
rect 41708 529484 41714 529486
rect 42425 529483 42491 529486
rect 673269 529138 673335 529141
rect 674005 529138 674071 529141
rect 676262 529138 676322 529176
rect 673269 529136 673378 529138
rect 673269 529080 673274 529136
rect 673330 529080 673378 529136
rect 673269 529075 673378 529080
rect 674005 529136 676322 529138
rect 674005 529080 674010 529136
rect 674066 529080 676322 529136
rect 674005 529078 676322 529080
rect 674005 529075 674071 529078
rect 41781 529004 41847 529005
rect 41781 529000 41828 529004
rect 41892 529002 41898 529004
rect 41781 528944 41786 529000
rect 41781 528940 41828 528944
rect 41892 528942 41938 529002
rect 41892 528940 41898 528942
rect 41781 528939 41847 528940
rect 42241 528866 42307 528869
rect 45185 528866 45251 528869
rect 42241 528864 45251 528866
rect 42241 528808 42246 528864
rect 42302 528808 45190 528864
rect 45246 528808 45251 528864
rect 673318 528866 673378 529075
rect 42241 528806 45251 528808
rect 42241 528803 42307 528806
rect 45185 528803 45251 528806
rect 62113 528594 62179 528597
rect 64646 528594 64706 528808
rect 673318 528806 676322 528866
rect 676262 528768 676322 528806
rect 62113 528592 64706 528594
rect 62113 528536 62118 528592
rect 62174 528536 64706 528592
rect 62113 528534 64706 528536
rect 62113 528531 62179 528534
rect 674005 528458 674071 528461
rect 674005 528456 676322 528458
rect 674005 528400 674010 528456
rect 674066 528400 676322 528456
rect 674005 528398 676322 528400
rect 674005 528395 674071 528398
rect 676262 528360 676322 528398
rect 684217 528186 684283 528189
rect 684174 528184 684283 528186
rect 684174 528128 684222 528184
rect 684278 528128 684283 528184
rect 684174 528123 684283 528128
rect 63401 528050 63467 528053
rect 63401 528048 64706 528050
rect 63401 527992 63406 528048
rect 63462 527992 64706 528048
rect 63401 527990 64706 527992
rect 63401 527987 63467 527990
rect 64646 527626 64706 527990
rect 684174 527952 684234 528123
rect 672901 527642 672967 527645
rect 672901 527640 676322 527642
rect 672901 527584 672906 527640
rect 672962 527584 676322 527640
rect 672901 527582 676322 527584
rect 672901 527579 672967 527582
rect 676262 527544 676322 527582
rect 683205 527370 683271 527373
rect 683205 527368 683314 527370
rect 683205 527312 683210 527368
rect 683266 527312 683314 527368
rect 683205 527307 683314 527312
rect 42609 527234 42675 527237
rect 45093 527234 45159 527237
rect 42609 527232 45159 527234
rect 42609 527176 42614 527232
rect 42670 527176 45098 527232
rect 45154 527176 45159 527232
rect 42609 527174 45159 527176
rect 42609 527171 42675 527174
rect 45093 527171 45159 527174
rect 683254 527136 683314 527307
rect 61377 527098 61443 527101
rect 61377 527096 64706 527098
rect 61377 527040 61382 527096
rect 61438 527040 64706 527096
rect 61377 527038 64706 527040
rect 61377 527035 61443 527038
rect 64646 526444 64706 527038
rect 683573 526962 683639 526965
rect 683573 526960 683682 526962
rect 683573 526904 683578 526960
rect 683634 526904 683682 526960
rect 683573 526899 683682 526904
rect 683622 526728 683682 526899
rect 683389 526554 683455 526557
rect 683389 526552 683498 526554
rect 683389 526496 683394 526552
rect 683450 526496 683498 526552
rect 683389 526491 683498 526496
rect 683438 526320 683498 526491
rect 677918 525741 677978 525912
rect 62941 525738 63007 525741
rect 62941 525736 64706 525738
rect 62941 525680 62946 525736
rect 63002 525680 64706 525736
rect 62941 525678 64706 525680
rect 62941 525675 63007 525678
rect 64646 525262 64706 525678
rect 677869 525736 677978 525741
rect 677869 525680 677874 525736
rect 677930 525680 677978 525736
rect 677869 525678 677978 525680
rect 677869 525675 677935 525678
rect 683070 524925 683130 525504
rect 683070 524920 683179 524925
rect 683070 524864 683118 524920
rect 683174 524864 683179 524920
rect 683070 524862 683179 524864
rect 683113 524859 683179 524862
rect 674005 524650 674071 524653
rect 675845 524650 675911 524653
rect 674005 524648 675911 524650
rect 674005 524592 674010 524648
rect 674066 524592 675850 524648
rect 675906 524592 675911 524648
rect 674005 524590 675911 524592
rect 674005 524587 674071 524590
rect 675845 524587 675911 524590
rect 677734 524517 677794 524688
rect 677685 524512 677794 524517
rect 677685 524456 677690 524512
rect 677746 524456 677794 524512
rect 677685 524454 677794 524456
rect 677685 524451 677751 524454
rect 675569 513770 675635 513773
rect 676029 513770 676095 513773
rect 675569 513768 676095 513770
rect 675569 513712 675574 513768
rect 675630 513712 676034 513768
rect 676090 513712 676095 513768
rect 675569 513710 676095 513712
rect 675569 513707 675635 513710
rect 676029 513707 676095 513710
rect 675201 508874 675267 508877
rect 676121 508874 676187 508877
rect 675201 508872 676187 508874
rect 675201 508816 675206 508872
rect 675262 508816 676126 508872
rect 676182 508816 676187 508872
rect 675201 508814 676187 508816
rect 675201 508811 675267 508814
rect 676121 508811 676187 508814
rect 675017 501938 675083 501941
rect 675845 501938 675911 501941
rect 675017 501936 675911 501938
rect 675017 501880 675022 501936
rect 675078 501880 675850 501936
rect 675906 501880 675911 501936
rect 675017 501878 675911 501880
rect 675017 501875 675083 501878
rect 675845 501875 675911 501878
rect 674373 492418 674439 492421
rect 676029 492418 676095 492421
rect 674373 492416 676095 492418
rect 674373 492360 674378 492416
rect 674434 492360 676034 492416
rect 676090 492360 676095 492416
rect 674373 492358 676095 492360
rect 674373 492355 674439 492358
rect 676029 492355 676095 492358
rect 673821 492146 673887 492149
rect 673821 492144 676292 492146
rect 673821 492088 673826 492144
rect 673882 492088 676292 492144
rect 673821 492086 676292 492088
rect 673821 492083 673887 492086
rect 674005 491738 674071 491741
rect 674005 491736 676292 491738
rect 674005 491680 674010 491736
rect 674066 491680 676292 491736
rect 674005 491678 676292 491680
rect 674005 491675 674071 491678
rect 672901 491330 672967 491333
rect 672901 491328 676292 491330
rect 672901 491272 672906 491328
rect 672962 491272 676292 491328
rect 672901 491270 676292 491272
rect 672901 491267 672967 491270
rect 674005 490922 674071 490925
rect 674005 490920 676292 490922
rect 674005 490864 674010 490920
rect 674066 490864 676292 490920
rect 674005 490862 676292 490864
rect 674005 490859 674071 490862
rect 675845 490514 675911 490517
rect 675845 490512 676292 490514
rect 675845 490456 675850 490512
rect 675906 490456 676292 490512
rect 675845 490454 676292 490456
rect 675845 490451 675911 490454
rect 674005 490106 674071 490109
rect 674005 490104 676292 490106
rect 674005 490048 674010 490104
rect 674066 490048 676292 490104
rect 674005 490046 676292 490048
rect 674005 490043 674071 490046
rect 674005 489698 674071 489701
rect 674005 489696 676292 489698
rect 674005 489640 674010 489696
rect 674066 489640 676292 489696
rect 674005 489638 676292 489640
rect 674005 489635 674071 489638
rect 674005 489290 674071 489293
rect 674005 489288 676292 489290
rect 674005 489232 674010 489288
rect 674066 489232 676292 489288
rect 674005 489230 676292 489232
rect 674005 489227 674071 489230
rect 675702 488820 675708 488884
rect 675772 488882 675778 488884
rect 675772 488822 676292 488882
rect 675772 488820 675778 488822
rect 674005 488474 674071 488477
rect 674005 488472 676292 488474
rect 674005 488416 674010 488472
rect 674066 488416 676292 488472
rect 674005 488414 676292 488416
rect 674005 488411 674071 488414
rect 676029 488066 676095 488069
rect 676029 488064 676292 488066
rect 676029 488008 676034 488064
rect 676090 488008 676292 488064
rect 676029 488006 676292 488008
rect 676029 488003 676095 488006
rect 675293 487658 675359 487661
rect 675293 487656 676292 487658
rect 675293 487600 675298 487656
rect 675354 487600 676292 487656
rect 675293 487598 676292 487600
rect 675293 487595 675359 487598
rect 678237 487250 678303 487253
rect 678237 487248 678316 487250
rect 678237 487192 678242 487248
rect 678298 487192 678316 487248
rect 678237 487190 678316 487192
rect 678237 487187 678303 487190
rect 683389 486842 683455 486845
rect 683389 486840 683468 486842
rect 683389 486784 683394 486840
rect 683450 486784 683468 486840
rect 683389 486782 683468 486784
rect 683389 486779 683455 486782
rect 680997 486434 681063 486437
rect 680997 486432 681076 486434
rect 680997 486376 681002 486432
rect 681058 486376 681076 486432
rect 680997 486374 681076 486376
rect 680997 486371 681063 486374
rect 674005 486026 674071 486029
rect 674005 486024 676292 486026
rect 674005 485968 674010 486024
rect 674066 485968 676292 486024
rect 674005 485966 676292 485968
rect 674005 485963 674071 485966
rect 673821 485618 673887 485621
rect 673821 485616 676292 485618
rect 673821 485560 673826 485616
rect 673882 485560 676292 485616
rect 673821 485558 676292 485560
rect 673821 485555 673887 485558
rect 674005 485210 674071 485213
rect 674005 485208 676292 485210
rect 674005 485152 674010 485208
rect 674066 485152 676292 485208
rect 674005 485150 676292 485152
rect 674005 485147 674071 485150
rect 676630 484567 676690 484772
rect 676581 484562 676690 484567
rect 676581 484506 676586 484562
rect 676642 484506 676690 484562
rect 676581 484504 676690 484506
rect 676581 484501 676647 484504
rect 673637 484394 673703 484397
rect 673637 484392 676292 484394
rect 673637 484336 673642 484392
rect 673698 484336 676292 484392
rect 673637 484334 676292 484336
rect 673637 484331 673703 484334
rect 675886 483924 675892 483988
rect 675956 483986 675962 483988
rect 675956 483926 676292 483986
rect 675956 483924 675962 483926
rect 675518 483516 675524 483580
rect 675588 483578 675594 483580
rect 675588 483518 676292 483578
rect 675588 483516 675594 483518
rect 673085 483170 673151 483173
rect 673085 483168 676292 483170
rect 673085 483112 673090 483168
rect 673146 483112 676292 483168
rect 673085 483110 676292 483112
rect 673085 483107 673151 483110
rect 674649 482762 674715 482765
rect 674649 482760 676292 482762
rect 674649 482704 674654 482760
rect 674710 482704 676292 482760
rect 674649 482702 676292 482704
rect 674649 482699 674715 482702
rect 674005 482354 674071 482357
rect 674005 482352 676292 482354
rect 674005 482296 674010 482352
rect 674066 482296 676292 482352
rect 674005 482294 676292 482296
rect 674005 482291 674071 482294
rect 675109 481946 675175 481949
rect 675109 481944 676292 481946
rect 675109 481888 675114 481944
rect 675170 481888 676292 481944
rect 675109 481886 676292 481888
rect 675109 481883 675175 481886
rect 677182 481130 677242 481508
rect 683113 481130 683179 481133
rect 677182 481128 683179 481130
rect 677182 481100 683118 481128
rect 677212 481072 683118 481100
rect 683174 481072 683179 481128
rect 677212 481070 683179 481072
rect 683113 481067 683179 481070
rect 675293 480722 675359 480725
rect 675293 480720 676292 480722
rect 675293 480664 675298 480720
rect 675354 480664 676292 480720
rect 675293 480662 676292 480664
rect 675293 480659 675359 480662
rect 674833 480042 674899 480045
rect 676121 480042 676187 480045
rect 674833 480040 676187 480042
rect 674833 479984 674838 480040
rect 674894 479984 676126 480040
rect 676182 479984 676187 480040
rect 674833 479982 676187 479984
rect 674833 479979 674899 479982
rect 676121 479979 676187 479982
rect 674598 477396 674604 477460
rect 674668 477458 674674 477460
rect 676213 477458 676279 477461
rect 674668 477456 676279 477458
rect 674668 477400 676218 477456
rect 676274 477400 676279 477456
rect 674668 477398 676279 477400
rect 674668 477396 674674 477398
rect 676213 477395 676279 477398
rect 673678 475356 673684 475420
rect 673748 475418 673754 475420
rect 674414 475418 674420 475420
rect 673748 475358 674420 475418
rect 673748 475356 673754 475358
rect 674414 475356 674420 475358
rect 674484 475356 674490 475420
rect 671470 474812 671476 474876
rect 671540 474874 671546 474876
rect 671981 474874 672047 474877
rect 671540 474872 672047 474874
rect 671540 474816 671986 474872
rect 672042 474816 672047 474872
rect 671540 474814 672047 474816
rect 671540 474812 671546 474814
rect 671981 474811 672047 474814
rect 673453 464810 673519 464813
rect 673678 464810 673684 464812
rect 673453 464808 673684 464810
rect 673453 464752 673458 464808
rect 673514 464752 673684 464808
rect 673453 464750 673684 464752
rect 673453 464747 673519 464750
rect 673678 464748 673684 464750
rect 673748 464748 673754 464812
rect 673821 455834 673887 455837
rect 676121 455834 676187 455837
rect 673821 455832 676187 455834
rect 673821 455776 673826 455832
rect 673882 455776 676126 455832
rect 676182 455776 676187 455832
rect 673821 455774 676187 455776
rect 673821 455771 673887 455774
rect 676121 455771 676187 455774
rect 669405 455426 669471 455429
rect 673269 455426 673335 455429
rect 669405 455424 673335 455426
rect 669405 455368 669410 455424
rect 669466 455368 673274 455424
rect 673330 455368 673335 455424
rect 669405 455366 673335 455368
rect 669405 455363 669471 455366
rect 673269 455363 673335 455366
rect 673269 455018 673335 455021
rect 673862 455018 673868 455020
rect 673269 455016 673868 455018
rect 673269 454960 673274 455016
rect 673330 454960 673868 455016
rect 673269 454958 673868 454960
rect 673269 454955 673335 454958
rect 673862 454956 673868 454958
rect 673932 454956 673938 455020
rect 673039 454610 673105 454613
rect 675661 454610 675727 454613
rect 673039 454608 675727 454610
rect 673039 454552 673044 454608
rect 673100 454552 675666 454608
rect 675722 454552 675727 454608
rect 673039 454550 675727 454552
rect 673039 454547 673105 454550
rect 675661 454547 675727 454550
rect 672947 454338 673013 454341
rect 674281 454338 674347 454341
rect 672947 454336 674347 454338
rect 672947 454280 672952 454336
rect 673008 454280 674286 454336
rect 674342 454280 674347 454336
rect 672947 454278 674347 454280
rect 672947 454275 673013 454278
rect 674281 454275 674347 454278
rect 672809 454066 672875 454069
rect 675293 454066 675359 454069
rect 672809 454064 675359 454066
rect 672809 454008 672814 454064
rect 672870 454008 675298 454064
rect 675354 454008 675359 454064
rect 672809 454006 675359 454008
rect 672809 454003 672875 454006
rect 675293 454003 675359 454006
rect 672441 453794 672507 453797
rect 675109 453794 675175 453797
rect 672441 453792 675175 453794
rect 672441 453736 672446 453792
rect 672502 453736 675114 453792
rect 675170 453736 675175 453792
rect 672441 453734 675175 453736
rect 672441 453731 672507 453734
rect 675109 453731 675175 453734
rect 675334 447748 675340 447812
rect 675404 447810 675410 447812
rect 675937 447810 676003 447813
rect 675404 447808 676003 447810
rect 675404 447752 675942 447808
rect 675998 447752 676003 447808
rect 675404 447750 676003 447752
rect 675404 447748 675410 447750
rect 675937 447747 676003 447750
rect 676806 440268 676812 440332
rect 676876 440330 676882 440332
rect 677501 440330 677567 440333
rect 676876 440328 677567 440330
rect 676876 440272 677506 440328
rect 677562 440272 677567 440328
rect 676876 440270 677567 440272
rect 676876 440268 676882 440270
rect 677501 440267 677567 440270
rect 41492 430886 55230 430946
rect 55170 430674 55230 430886
rect 59997 430674 60063 430677
rect 55170 430672 60063 430674
rect 55170 430616 60002 430672
rect 60058 430616 60063 430672
rect 55170 430614 60063 430616
rect 59997 430611 60063 430614
rect 41492 430478 45570 430538
rect 35801 430130 35867 430133
rect 35788 430128 35867 430130
rect 35788 430072 35806 430128
rect 35862 430072 35867 430128
rect 35788 430070 35867 430072
rect 35801 430067 35867 430070
rect 44541 429722 44607 429725
rect 41492 429720 44607 429722
rect 41492 429664 44546 429720
rect 44602 429664 44607 429720
rect 41492 429662 44607 429664
rect 44541 429659 44607 429662
rect 44633 429314 44699 429317
rect 41492 429312 44699 429314
rect 41492 429256 44638 429312
rect 44694 429256 44699 429312
rect 41492 429254 44699 429256
rect 45510 429314 45570 430478
rect 61377 429314 61443 429317
rect 45510 429312 61443 429314
rect 45510 429256 61382 429312
rect 61438 429256 61443 429312
rect 45510 429254 61443 429256
rect 44633 429251 44699 429254
rect 61377 429251 61443 429254
rect 44265 428906 44331 428909
rect 41492 428904 44331 428906
rect 41492 428848 44270 428904
rect 44326 428848 44331 428904
rect 41492 428846 44331 428848
rect 44265 428843 44331 428846
rect 44265 428498 44331 428501
rect 41492 428496 44331 428498
rect 41492 428440 44270 428496
rect 44326 428440 44331 428496
rect 41492 428438 44331 428440
rect 44265 428435 44331 428438
rect 45645 428090 45711 428093
rect 41492 428088 45711 428090
rect 41492 428032 45650 428088
rect 45706 428032 45711 428088
rect 41492 428030 45711 428032
rect 45645 428027 45711 428030
rect 45553 427682 45619 427685
rect 41492 427680 45619 427682
rect 41492 427624 45558 427680
rect 45614 427624 45619 427680
rect 41492 427622 45619 427624
rect 45553 427619 45619 427622
rect 45829 427410 45895 427413
rect 41784 427408 45895 427410
rect 41784 427352 45834 427408
rect 45890 427352 45895 427408
rect 41784 427350 45895 427352
rect 41784 427274 41844 427350
rect 45829 427347 45895 427350
rect 41492 427214 41844 427274
rect 41965 427138 42031 427141
rect 63125 427138 63191 427141
rect 41965 427136 63191 427138
rect 41965 427080 41970 427136
rect 42026 427080 63130 427136
rect 63186 427080 63191 427136
rect 41965 427078 63191 427080
rect 41965 427075 42031 427078
rect 63125 427075 63191 427078
rect 45829 426866 45895 426869
rect 41492 426864 45895 426866
rect 41492 426808 45834 426864
rect 45890 426808 45895 426864
rect 41492 426806 45895 426808
rect 45829 426803 45895 426806
rect 41822 426458 41828 426460
rect 41492 426398 41828 426458
rect 41822 426396 41828 426398
rect 41892 426396 41898 426460
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 41137 425642 41203 425645
rect 41124 425640 41203 425642
rect 41124 425584 41142 425640
rect 41198 425584 41203 425640
rect 41124 425582 41203 425584
rect 41137 425579 41203 425582
rect 40953 425234 41019 425237
rect 40940 425232 41019 425234
rect 40940 425176 40958 425232
rect 41014 425176 41019 425232
rect 40940 425174 41019 425176
rect 40953 425171 41019 425174
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 32029 424418 32095 424421
rect 32029 424416 32108 424418
rect 32029 424360 32034 424416
rect 32090 424360 32108 424416
rect 32029 424358 32108 424360
rect 32029 424355 32095 424358
rect 41873 424282 41939 424285
rect 42190 424282 42196 424284
rect 41873 424280 42196 424282
rect 41873 424224 41878 424280
rect 41934 424224 42196 424280
rect 41873 424222 42196 424224
rect 41873 424219 41939 424222
rect 42190 424220 42196 424222
rect 42260 424220 42266 424284
rect 46013 424010 46079 424013
rect 41492 424008 46079 424010
rect 41492 423952 46018 424008
rect 46074 423952 46079 424008
rect 41492 423950 46079 423952
rect 46013 423947 46079 423950
rect 42793 423602 42859 423605
rect 41492 423600 42859 423602
rect 41492 423544 42798 423600
rect 42854 423544 42859 423600
rect 41492 423542 42859 423544
rect 42793 423539 42859 423542
rect 45001 423194 45067 423197
rect 41492 423192 45067 423194
rect 41492 423136 45006 423192
rect 45062 423136 45067 423192
rect 41492 423134 45067 423136
rect 45001 423131 45067 423134
rect 41822 422786 41828 422788
rect 41492 422726 41828 422786
rect 41822 422724 41828 422726
rect 41892 422724 41898 422788
rect 44449 422378 44515 422381
rect 41492 422376 44515 422378
rect 41492 422320 44454 422376
rect 44510 422320 44515 422376
rect 41492 422318 44515 422320
rect 44449 422315 44515 422318
rect 41822 421970 41828 421972
rect 41492 421910 41828 421970
rect 41822 421908 41828 421910
rect 41892 421908 41898 421972
rect 45369 421562 45435 421565
rect 41492 421560 45435 421562
rect 41492 421504 45374 421560
rect 45430 421504 45435 421560
rect 41492 421502 45435 421504
rect 45369 421499 45435 421502
rect 45185 421154 45251 421157
rect 41492 421152 45251 421154
rect 41492 421096 45190 421152
rect 45246 421096 45251 421152
rect 41492 421094 45251 421096
rect 45185 421091 45251 421094
rect 43253 420746 43319 420749
rect 41492 420744 43319 420746
rect 41492 420688 43258 420744
rect 43314 420688 43319 420744
rect 41492 420686 43319 420688
rect 43253 420683 43319 420686
rect 41462 419930 41522 420308
rect 42517 419930 42583 419933
rect 41462 419928 42583 419930
rect 41462 419900 42522 419928
rect 41492 419872 42522 419900
rect 42578 419872 42583 419928
rect 41492 419870 42583 419872
rect 42517 419867 42583 419870
rect 43069 419522 43135 419525
rect 41492 419520 43135 419522
rect 41492 419464 43074 419520
rect 43130 419464 43135 419520
rect 41492 419462 43135 419464
rect 43069 419459 43135 419462
rect 41137 418842 41203 418845
rect 41454 418842 41460 418844
rect 41137 418840 41460 418842
rect 41137 418784 41142 418840
rect 41198 418784 41460 418840
rect 41137 418782 41460 418784
rect 41137 418779 41203 418782
rect 41454 418780 41460 418782
rect 41524 418780 41530 418844
rect 41638 413340 41644 413404
rect 41708 413402 41714 413404
rect 42190 413402 42196 413404
rect 41708 413342 42196 413402
rect 41708 413340 41714 413342
rect 42190 413340 42196 413342
rect 42260 413340 42266 413404
rect 42057 411906 42123 411909
rect 42517 411906 42583 411909
rect 42057 411904 42583 411906
rect 42057 411848 42062 411904
rect 42118 411848 42522 411904
rect 42578 411848 42583 411904
rect 42057 411846 42583 411848
rect 42057 411843 42123 411846
rect 42517 411843 42583 411846
rect 675334 410484 675340 410548
rect 675404 410546 675410 410548
rect 676029 410546 676095 410549
rect 675404 410544 676095 410546
rect 675404 410488 676034 410544
rect 676090 410488 676095 410544
rect 675404 410486 676095 410488
rect 675404 410484 675410 410486
rect 676029 410483 676095 410486
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 41965 408098 42031 408101
rect 45185 408098 45251 408101
rect 41965 408096 45251 408098
rect 41965 408040 41970 408096
rect 42026 408040 45190 408096
rect 45246 408040 45251 408096
rect 41965 408038 45251 408040
rect 41965 408035 42031 408038
rect 45185 408035 45251 408038
rect 42425 407826 42491 407829
rect 53833 407826 53899 407829
rect 42425 407824 53899 407826
rect 42425 407768 42430 407824
rect 42486 407768 53838 407824
rect 53894 407768 53899 407824
rect 42425 407766 53899 407768
rect 42425 407763 42491 407766
rect 53833 407763 53899 407766
rect 42241 407554 42307 407557
rect 44449 407554 44515 407557
rect 42241 407552 44515 407554
rect 42241 407496 42246 407552
rect 42302 407496 44454 407552
rect 44510 407496 44515 407552
rect 42241 407494 44515 407496
rect 42241 407491 42307 407494
rect 44449 407491 44515 407494
rect 42057 406738 42123 406741
rect 45369 406738 45435 406741
rect 42057 406736 45435 406738
rect 42057 406680 42062 406736
rect 42118 406680 45374 406736
rect 45430 406680 45435 406736
rect 42057 406678 45435 406680
rect 42057 406675 42123 406678
rect 45369 406675 45435 406678
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 40902 405588 40908 405652
rect 40972 405650 40978 405652
rect 42241 405650 42307 405653
rect 40972 405648 42307 405650
rect 40972 405592 42246 405648
rect 42302 405592 42307 405648
rect 40972 405590 42307 405592
rect 40972 405588 40978 405590
rect 42241 405587 42307 405590
rect 42425 405650 42491 405653
rect 44817 405650 44883 405653
rect 42425 405648 44883 405650
rect 42425 405592 42430 405648
rect 42486 405592 44822 405648
rect 44878 405592 44883 405648
rect 42425 405590 44883 405592
rect 42425 405587 42491 405590
rect 44817 405587 44883 405590
rect 62113 404154 62179 404157
rect 62113 404152 64706 404154
rect 62113 404096 62118 404152
rect 62174 404096 64706 404152
rect 62113 404094 64706 404096
rect 62113 404091 62179 404094
rect 64646 403550 64706 404094
rect 676262 403746 676322 403852
rect 663750 403686 676322 403746
rect 657537 403338 657603 403341
rect 663750 403338 663810 403686
rect 674557 403474 674623 403477
rect 674557 403472 676292 403474
rect 674557 403416 674562 403472
rect 674618 403416 676292 403472
rect 674557 403414 676292 403416
rect 674557 403411 674623 403414
rect 657537 403336 663810 403338
rect 657537 403280 657542 403336
rect 657598 403280 663810 403336
rect 657537 403278 663810 403280
rect 657537 403275 657603 403278
rect 676630 402933 676690 403036
rect 42333 402930 42399 402933
rect 45001 402930 45067 402933
rect 42333 402928 45067 402930
rect 42333 402872 42338 402928
rect 42394 402872 45006 402928
rect 45062 402872 45067 402928
rect 42333 402870 45067 402872
rect 42333 402867 42399 402870
rect 45001 402867 45067 402870
rect 676581 402928 676690 402933
rect 676581 402872 676586 402928
rect 676642 402872 676690 402928
rect 676581 402870 676690 402872
rect 676581 402867 676647 402870
rect 62113 402658 62179 402661
rect 676029 402658 676095 402661
rect 62113 402656 64706 402658
rect 62113 402600 62118 402656
rect 62174 402600 64706 402656
rect 62113 402598 64706 402600
rect 62113 402595 62179 402598
rect 64646 402368 64706 402598
rect 676029 402656 676292 402658
rect 676029 402600 676034 402656
rect 676090 402600 676292 402656
rect 676029 402598 676292 402600
rect 676029 402595 676095 402598
rect 674833 402250 674899 402253
rect 674833 402248 676292 402250
rect 674833 402192 674838 402248
rect 674894 402192 676292 402248
rect 674833 402190 676292 402192
rect 674833 402187 674899 402190
rect 672625 401978 672691 401981
rect 672625 401976 676322 401978
rect 672625 401920 672630 401976
rect 672686 401920 676322 401976
rect 672625 401918 676322 401920
rect 672625 401915 672691 401918
rect 41781 401844 41847 401845
rect 41781 401840 41828 401844
rect 41892 401842 41898 401844
rect 41781 401784 41786 401840
rect 41781 401780 41828 401784
rect 41892 401782 41938 401842
rect 676262 401812 676322 401918
rect 41892 401780 41898 401782
rect 41781 401779 41847 401780
rect 672809 401706 672875 401709
rect 674833 401706 674899 401709
rect 672809 401704 674899 401706
rect 672809 401648 672814 401704
rect 672870 401648 674838 401704
rect 674894 401648 674899 401704
rect 672809 401646 674899 401648
rect 672809 401643 672875 401646
rect 674833 401643 674899 401646
rect 673177 401298 673243 401301
rect 676262 401298 676322 401404
rect 673177 401296 676322 401298
rect 673177 401240 673182 401296
rect 673238 401240 676322 401296
rect 673177 401238 676322 401240
rect 673177 401235 673243 401238
rect 677174 401236 677180 401300
rect 677244 401236 677250 401300
rect 62113 400618 62179 400621
rect 64646 400618 64706 401186
rect 677182 400996 677242 401236
rect 652017 400890 652083 400893
rect 676581 400890 676647 400893
rect 652017 400888 676647 400890
rect 652017 400832 652022 400888
rect 652078 400832 676586 400888
rect 676642 400832 676647 400888
rect 652017 400830 676647 400832
rect 652017 400827 652083 400830
rect 676581 400827 676647 400830
rect 62113 400616 64706 400618
rect 62113 400560 62118 400616
rect 62174 400560 64706 400616
rect 62113 400558 64706 400560
rect 673361 400618 673427 400621
rect 673361 400616 676292 400618
rect 673361 400560 673366 400616
rect 673422 400560 676292 400616
rect 673361 400558 676292 400560
rect 62113 400555 62179 400558
rect 673361 400555 673427 400558
rect 676806 400420 676812 400484
rect 676876 400420 676882 400484
rect 42425 400210 42491 400213
rect 46013 400210 46079 400213
rect 42425 400208 46079 400210
rect 42425 400152 42430 400208
rect 42486 400152 46018 400208
rect 46074 400152 46079 400208
rect 42425 400150 46079 400152
rect 42425 400147 42491 400150
rect 46013 400147 46079 400150
rect 63125 400210 63191 400213
rect 63125 400208 64706 400210
rect 63125 400152 63130 400208
rect 63186 400152 64706 400208
rect 676814 400180 676874 400420
rect 63125 400150 64706 400152
rect 63125 400147 63191 400150
rect 40534 400012 40540 400076
rect 40604 400074 40610 400076
rect 41781 400074 41847 400077
rect 40604 400072 41847 400074
rect 40604 400016 41786 400072
rect 41842 400016 41847 400072
rect 40604 400014 41847 400016
rect 40604 400012 40610 400014
rect 41781 400011 41847 400014
rect 64646 400004 64706 400150
rect 673913 399802 673979 399805
rect 673913 399800 676292 399802
rect 673913 399744 673918 399800
rect 673974 399744 676292 399800
rect 673913 399742 676292 399744
rect 673913 399739 673979 399742
rect 62113 399394 62179 399397
rect 674833 399394 674899 399397
rect 62113 399392 64706 399394
rect 62113 399336 62118 399392
rect 62174 399336 64706 399392
rect 62113 399334 64706 399336
rect 62113 399331 62179 399334
rect 41454 398788 41460 398852
rect 41524 398850 41530 398852
rect 41781 398850 41847 398853
rect 41524 398848 41847 398850
rect 41524 398792 41786 398848
rect 41842 398792 41847 398848
rect 64646 398822 64706 399334
rect 674833 399392 676292 399394
rect 674833 399336 674838 399392
rect 674894 399336 676292 399392
rect 674833 399334 676292 399336
rect 674833 399331 674899 399334
rect 41524 398790 41847 398792
rect 41524 398788 41530 398790
rect 41781 398787 41847 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 61377 398306 61443 398309
rect 61377 398304 64706 398306
rect 61377 398248 61382 398304
rect 61438 398248 64706 398304
rect 61377 398246 64706 398248
rect 61377 398243 61443 398246
rect 64646 397640 64706 398246
rect 675017 398170 675083 398173
rect 675017 398168 676292 398170
rect 675017 398112 675022 398168
rect 675078 398112 676292 398168
rect 675017 398110 676292 398112
rect 675017 398107 675083 398110
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 671981 397218 672047 397221
rect 676262 397218 676322 397324
rect 671981 397216 676322 397218
rect 671981 397160 671986 397216
rect 672042 397160 676322 397216
rect 671981 397158 676322 397160
rect 671981 397155 672047 397158
rect 676262 396812 676322 396916
rect 676254 396748 676260 396812
rect 676324 396748 676330 396812
rect 674373 396538 674439 396541
rect 674373 396536 676292 396538
rect 674373 396480 674378 396536
rect 674434 396480 676292 396536
rect 674373 396478 676292 396480
rect 674373 396475 674439 396478
rect 676446 395996 676506 396100
rect 676438 395932 676444 395996
rect 676508 395932 676514 395996
rect 42149 395722 42215 395725
rect 51073 395722 51139 395725
rect 42149 395720 51139 395722
rect 42149 395664 42154 395720
rect 42210 395664 51078 395720
rect 51134 395664 51139 395720
rect 42149 395662 51139 395664
rect 42149 395659 42215 395662
rect 51073 395659 51139 395662
rect 674741 395722 674807 395725
rect 674741 395720 676292 395722
rect 674741 395664 674746 395720
rect 674802 395664 676292 395720
rect 674741 395662 676292 395664
rect 674741 395659 674807 395662
rect 652201 395314 652267 395317
rect 674557 395314 674623 395317
rect 652201 395312 674623 395314
rect 652201 395256 652206 395312
rect 652262 395256 674562 395312
rect 674618 395256 674623 395312
rect 652201 395254 674623 395256
rect 652201 395251 652267 395254
rect 674557 395251 674623 395254
rect 676630 395180 676690 395284
rect 676622 395116 676628 395180
rect 676692 395116 676698 395180
rect 672993 394770 673059 394773
rect 676262 394770 676322 394876
rect 672993 394768 676322 394770
rect 672993 394712 672998 394768
rect 673054 394712 676322 394768
rect 672993 394710 676322 394712
rect 672993 394707 673059 394710
rect 674281 394498 674347 394501
rect 674281 394496 676292 394498
rect 674281 394440 674286 394496
rect 674342 394440 676292 394496
rect 674281 394438 676292 394440
rect 674281 394435 674347 394438
rect 676029 394090 676095 394093
rect 676029 394088 676292 394090
rect 676029 394032 676034 394088
rect 676090 394032 676292 394088
rect 676029 394030 676292 394032
rect 676029 394027 676095 394030
rect 669221 393546 669287 393549
rect 676262 393546 676322 393652
rect 669221 393544 676322 393546
rect 669221 393488 669226 393544
rect 669282 393488 676322 393544
rect 669221 393486 676322 393488
rect 669221 393483 669287 393486
rect 673729 393138 673795 393141
rect 676029 393138 676095 393141
rect 673729 393136 676095 393138
rect 673729 393080 673734 393136
rect 673790 393080 676034 393136
rect 676090 393080 676095 393136
rect 673729 393078 676095 393080
rect 673729 393075 673795 393078
rect 676029 393075 676095 393078
rect 683070 392733 683130 393244
rect 683021 392728 683130 392733
rect 683021 392672 683026 392728
rect 683082 392672 683130 392728
rect 683021 392670 683130 392672
rect 683021 392667 683087 392670
rect 670601 392322 670667 392325
rect 676262 392322 676322 392428
rect 670601 392320 676322 392322
rect 670601 392264 670606 392320
rect 670662 392264 676322 392320
rect 670601 392262 676322 392264
rect 670601 392259 670667 392262
rect 675886 389812 675892 389876
rect 675956 389874 675962 389876
rect 683021 389874 683087 389877
rect 675956 389872 683087 389874
rect 675956 389816 683026 389872
rect 683082 389816 683087 389872
rect 675956 389814 683087 389816
rect 675956 389812 675962 389814
rect 683021 389811 683087 389814
rect 675702 388452 675708 388516
rect 675772 388514 675778 388516
rect 680997 388514 681063 388517
rect 675772 388512 681063 388514
rect 675772 388456 681002 388512
rect 681058 388456 681063 388512
rect 675772 388454 681063 388456
rect 675772 388452 675778 388454
rect 680997 388451 681063 388454
rect 41462 387562 41522 387668
rect 41462 387502 51090 387562
rect 41094 387157 41154 387260
rect 41094 387152 41203 387157
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387094 41203 387096
rect 41137 387091 41203 387094
rect 41278 386749 41338 386852
rect 41278 386744 41387 386749
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386686 41387 386688
rect 41321 386683 41387 386686
rect 44633 386474 44699 386477
rect 41492 386472 44699 386474
rect 41492 386416 44638 386472
rect 44694 386416 44699 386472
rect 41492 386414 44699 386416
rect 51030 386474 51090 387502
rect 61377 386474 61443 386477
rect 51030 386472 61443 386474
rect 51030 386416 61382 386472
rect 61438 386416 61443 386472
rect 51030 386414 61443 386416
rect 44633 386411 44699 386414
rect 61377 386411 61443 386414
rect 668853 386066 668919 386069
rect 675385 386066 675451 386069
rect 668853 386064 675451 386066
rect 40726 385933 40786 386036
rect 668853 386008 668858 386064
rect 668914 386008 675390 386064
rect 675446 386008 675451 386064
rect 668853 386006 675451 386008
rect 668853 386003 668919 386006
rect 675385 386003 675451 386006
rect 40726 385928 40835 385933
rect 40726 385872 40774 385928
rect 40830 385872 40835 385928
rect 40726 385870 40835 385872
rect 40769 385867 40835 385870
rect 41321 385930 41387 385933
rect 63401 385930 63467 385933
rect 41321 385928 63467 385930
rect 41321 385872 41326 385928
rect 41382 385872 63406 385928
rect 63462 385872 63467 385928
rect 41321 385870 63467 385872
rect 41321 385867 41387 385870
rect 63401 385867 63467 385870
rect 44265 385658 44331 385661
rect 41492 385656 44331 385658
rect 41492 385600 44270 385656
rect 44326 385600 44331 385656
rect 41492 385598 44331 385600
rect 44265 385595 44331 385598
rect 675753 385386 675819 385389
rect 676254 385386 676260 385388
rect 675753 385384 676260 385386
rect 675753 385328 675758 385384
rect 675814 385328 676260 385384
rect 675753 385326 676260 385328
rect 675753 385323 675819 385326
rect 676254 385324 676260 385326
rect 676324 385324 676330 385388
rect 45093 385250 45159 385253
rect 41492 385248 45159 385250
rect 41492 385192 45098 385248
rect 45154 385192 45159 385248
rect 41492 385190 45159 385192
rect 45093 385187 45159 385190
rect 45553 384842 45619 384845
rect 41492 384840 45619 384842
rect 41492 384784 45558 384840
rect 45614 384784 45619 384840
rect 41492 384782 45619 384784
rect 45553 384779 45619 384782
rect 46013 384434 46079 384437
rect 41492 384432 46079 384434
rect 41492 384376 46018 384432
rect 46074 384376 46079 384432
rect 41492 384374 46079 384376
rect 46013 384371 46079 384374
rect 45829 384026 45895 384029
rect 41492 384024 45895 384026
rect 41492 383968 45834 384024
rect 45890 383968 45895 384024
rect 41492 383966 45895 383968
rect 45829 383963 45895 383966
rect 45645 383618 45711 383621
rect 41492 383616 45711 383618
rect 41492 383560 45650 383616
rect 45706 383560 45711 383616
rect 41492 383558 45711 383560
rect 45645 383555 45711 383558
rect 47117 383210 47183 383213
rect 41492 383208 47183 383210
rect 41492 383152 47122 383208
rect 47178 383152 47183 383208
rect 41492 383150 47183 383152
rect 47117 383147 47183 383150
rect 654777 382938 654843 382941
rect 668853 382938 668919 382941
rect 654777 382936 668919 382938
rect 654777 382880 654782 382936
rect 654838 382880 668858 382936
rect 668914 382880 668919 382936
rect 654777 382878 668919 382880
rect 654777 382875 654843 382878
rect 668853 382875 668919 382878
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 46933 382394 46999 382397
rect 41492 382392 46999 382394
rect 41492 382336 46938 382392
rect 46994 382336 46999 382392
rect 41492 382334 46999 382336
rect 46933 382331 46999 382334
rect 40910 381853 40970 381956
rect 40910 381848 41019 381853
rect 40910 381792 40958 381848
rect 41014 381792 41019 381848
rect 40910 381790 41019 381792
rect 40953 381787 41019 381790
rect 41137 381850 41203 381853
rect 62941 381850 63007 381853
rect 41137 381848 63007 381850
rect 41137 381792 41142 381848
rect 41198 381792 62946 381848
rect 63002 381792 63007 381848
rect 41137 381790 63007 381792
rect 41137 381787 41203 381790
rect 62941 381787 63007 381790
rect 675753 381714 675819 381717
rect 676438 381714 676444 381716
rect 675753 381712 676444 381714
rect 675753 381656 675758 381712
rect 675814 381656 676444 381712
rect 675753 381654 676444 381656
rect 675753 381651 675819 381654
rect 676438 381652 676444 381654
rect 676508 381652 676514 381716
rect 40174 381445 40234 381548
rect 40174 381440 40283 381445
rect 40174 381384 40222 381440
rect 40278 381384 40283 381440
rect 40174 381382 40283 381384
rect 40217 381379 40283 381382
rect 40769 381442 40835 381445
rect 45277 381442 45343 381445
rect 40769 381440 45343 381442
rect 40769 381384 40774 381440
rect 40830 381384 45282 381440
rect 45338 381384 45343 381440
rect 40769 381382 45343 381384
rect 40769 381379 40835 381382
rect 45277 381379 45343 381382
rect 35206 381037 35266 381140
rect 35157 381032 35266 381037
rect 35157 380976 35162 381032
rect 35218 380976 35266 381032
rect 35157 380974 35266 380976
rect 672993 381034 673059 381037
rect 675385 381034 675451 381037
rect 672993 381032 675451 381034
rect 672993 380976 672998 381032
rect 673054 380976 675390 381032
rect 675446 380976 675451 381032
rect 672993 380974 675451 380976
rect 35157 380971 35223 380974
rect 672993 380971 673059 380974
rect 675385 380971 675451 380974
rect 40542 380628 40602 380732
rect 40534 380564 40540 380628
rect 40604 380564 40610 380628
rect 37966 380221 38026 380324
rect 37917 380216 38026 380221
rect 37917 380160 37922 380216
rect 37978 380160 38026 380216
rect 37917 380158 38026 380160
rect 37917 380155 37983 380158
rect 33734 379813 33794 379916
rect 33734 379808 33843 379813
rect 33734 379752 33782 379808
rect 33838 379752 33843 379808
rect 33734 379750 33843 379752
rect 33777 379747 33843 379750
rect 40953 379810 41019 379813
rect 41454 379810 41460 379812
rect 40953 379808 41460 379810
rect 40953 379752 40958 379808
rect 41014 379752 41460 379808
rect 40953 379750 41460 379752
rect 40953 379747 41019 379750
rect 41454 379748 41460 379750
rect 41524 379748 41530 379812
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 40585 379402 40651 379405
rect 42885 379402 42951 379405
rect 40585 379400 42951 379402
rect 40585 379344 40590 379400
rect 40646 379344 42890 379400
rect 42946 379344 42951 379400
rect 40585 379342 42951 379344
rect 40585 379339 40651 379342
rect 42885 379339 42951 379342
rect 44357 379130 44423 379133
rect 41492 379128 44423 379130
rect 41492 379072 44362 379128
rect 44418 379072 44423 379128
rect 41492 379070 44423 379072
rect 44357 379067 44423 379070
rect 44541 378722 44607 378725
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 41492 378720 44607 378722
rect 41492 378664 44546 378720
rect 44602 378664 44607 378720
rect 41492 378662 44607 378664
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 44541 378659 44607 378662
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 44725 377906 44791 377909
rect 41492 377904 44791 377906
rect 41492 377848 44730 377904
rect 44786 377848 44791 377904
rect 41492 377846 44791 377848
rect 44725 377843 44791 377846
rect 44909 377498 44975 377501
rect 41492 377496 44975 377498
rect 41492 377440 44914 377496
rect 44970 377440 44975 377496
rect 41492 377438 44975 377440
rect 44909 377435 44975 377438
rect 675753 377362 675819 377365
rect 676622 377362 676628 377364
rect 675753 377360 676628 377362
rect 675753 377304 675758 377360
rect 675814 377304 676628 377360
rect 675753 377302 676628 377304
rect 675753 377299 675819 377302
rect 676622 377300 676628 377302
rect 676692 377300 676698 377364
rect 35758 376549 35818 377060
rect 673729 376682 673795 376685
rect 675109 376682 675175 376685
rect 673729 376680 675175 376682
rect 673729 376624 673734 376680
rect 673790 376624 675114 376680
rect 675170 376624 675175 376680
rect 673729 376622 675175 376624
rect 673729 376619 673795 376622
rect 675109 376619 675175 376622
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 35801 376483 35867 376486
rect 44173 376274 44239 376277
rect 41492 376272 44239 376274
rect 41492 376216 44178 376272
rect 44234 376216 44239 376272
rect 41492 376214 44239 376216
rect 44173 376211 44239 376214
rect 35801 374642 35867 374645
rect 41270 374642 41276 374644
rect 35801 374640 41276 374642
rect 35801 374584 35806 374640
rect 35862 374584 41276 374640
rect 35801 374582 41276 374584
rect 35801 374579 35867 374582
rect 41270 374580 41276 374582
rect 41340 374580 41346 374644
rect 652201 373962 652267 373965
rect 649950 373960 652267 373962
rect 649950 373904 652206 373960
rect 652262 373904 652267 373960
rect 649950 373902 652267 373904
rect 649950 373892 650010 373902
rect 652201 373899 652267 373902
rect 675753 373690 675819 373693
rect 676070 373690 676076 373692
rect 675753 373688 676076 373690
rect 675753 373632 675758 373688
rect 675814 373632 676076 373688
rect 675753 373630 676076 373632
rect 675753 373627 675819 373630
rect 676070 373628 676076 373630
rect 676140 373628 676146 373692
rect 651465 373282 651531 373285
rect 649950 373280 651531 373282
rect 649950 373224 651470 373280
rect 651526 373224 651531 373280
rect 649950 373222 651531 373224
rect 37917 372738 37983 372741
rect 41638 372738 41644 372740
rect 37917 372736 41644 372738
rect 37917 372680 37922 372736
rect 37978 372680 41644 372736
rect 37917 372678 41644 372680
rect 37917 372675 37983 372678
rect 41638 372676 41644 372678
rect 41708 372676 41714 372740
rect 649950 372710 650010 373222
rect 651465 373219 651531 373222
rect 675661 373010 675727 373013
rect 675886 373010 675892 373012
rect 675661 373008 675892 373010
rect 675661 372952 675666 373008
rect 675722 372952 675892 373008
rect 675661 372950 675892 372952
rect 675661 372947 675727 372950
rect 675886 372948 675892 372950
rect 675956 372948 675962 373012
rect 671981 372602 672047 372605
rect 675109 372602 675175 372605
rect 671981 372600 675175 372602
rect 671981 372544 671986 372600
rect 672042 372544 675114 372600
rect 675170 372544 675175 372600
rect 671981 372542 675175 372544
rect 671981 372539 672047 372542
rect 675109 372539 675175 372542
rect 652017 372194 652083 372197
rect 649950 372192 652083 372194
rect 649950 372136 652022 372192
rect 652078 372136 652083 372192
rect 649950 372134 652083 372136
rect 33777 371922 33843 371925
rect 41822 371922 41828 371924
rect 33777 371920 41828 371922
rect 33777 371864 33782 371920
rect 33838 371864 41828 371920
rect 33777 371862 41828 371864
rect 33777 371859 33843 371862
rect 41822 371860 41828 371862
rect 41892 371860 41898 371924
rect 649950 371528 650010 372134
rect 652017 372131 652083 372134
rect 651465 370698 651531 370701
rect 649950 370696 651531 370698
rect 649950 370640 651470 370696
rect 651526 370640 651531 370696
rect 649950 370638 651531 370640
rect 649950 370346 650010 370638
rect 651465 370635 651531 370638
rect 41270 368460 41276 368524
rect 41340 368522 41346 368524
rect 41781 368522 41847 368525
rect 41340 368520 41847 368522
rect 41340 368464 41786 368520
rect 41842 368464 41847 368520
rect 41340 368462 41847 368464
rect 41340 368460 41346 368462
rect 41781 368459 41847 368462
rect 42057 366210 42123 366213
rect 42885 366210 42951 366213
rect 42057 366208 42951 366210
rect 42057 366152 42062 366208
rect 42118 366152 42890 366208
rect 42946 366152 42951 366208
rect 42057 366150 42951 366152
rect 42057 366147 42123 366150
rect 42885 366147 42951 366150
rect 42057 364850 42123 364853
rect 44725 364850 44791 364853
rect 42057 364848 44791 364850
rect 42057 364792 42062 364848
rect 42118 364792 44730 364848
rect 44786 364792 44791 364848
rect 42057 364790 44791 364792
rect 42057 364787 42123 364790
rect 44725 364787 44791 364790
rect 42241 364170 42307 364173
rect 44357 364170 44423 364173
rect 42241 364168 44423 364170
rect 42241 364112 42246 364168
rect 42302 364112 44362 364168
rect 44418 364112 44423 364168
rect 42241 364110 44423 364112
rect 42241 364107 42307 364110
rect 44357 364107 44423 364110
rect 40718 363700 40724 363764
rect 40788 363762 40794 363764
rect 41781 363762 41847 363765
rect 40788 363760 41847 363762
rect 40788 363704 41786 363760
rect 41842 363704 41847 363760
rect 40788 363702 41847 363704
rect 40788 363700 40794 363702
rect 41781 363699 41847 363702
rect 42701 363218 42767 363221
rect 46565 363218 46631 363221
rect 42701 363216 46631 363218
rect 42701 363160 42706 363216
rect 42762 363160 46570 363216
rect 46626 363160 46631 363216
rect 42701 363158 46631 363160
rect 42701 363155 42767 363158
rect 46565 363155 46631 363158
rect 42241 362946 42307 362949
rect 45369 362946 45435 362949
rect 42241 362944 45435 362946
rect 42241 362888 42246 362944
rect 42302 362888 45374 362944
rect 45430 362888 45435 362944
rect 42241 362886 45435 362888
rect 42241 362883 42307 362886
rect 45369 362883 45435 362886
rect 42425 361586 42491 361589
rect 44541 361586 44607 361589
rect 42425 361584 44607 361586
rect 42425 361528 42430 361584
rect 42486 361528 44546 361584
rect 44602 361528 44607 361584
rect 42425 361526 44607 361528
rect 42425 361523 42491 361526
rect 44541 361523 44607 361526
rect 62113 360906 62179 360909
rect 62113 360904 64706 360906
rect 62113 360848 62118 360904
rect 62174 360848 64706 360904
rect 62113 360846 64706 360848
rect 62113 360843 62179 360846
rect 64646 360328 64706 360846
rect 41781 360092 41847 360093
rect 41781 360088 41828 360092
rect 41892 360090 41898 360092
rect 41781 360032 41786 360088
rect 41781 360028 41828 360032
rect 41892 360030 41938 360090
rect 41892 360028 41898 360030
rect 41781 360027 41847 360028
rect 62113 359818 62179 359821
rect 62113 359816 64706 359818
rect 62113 359760 62118 359816
rect 62174 359760 64706 359816
rect 62113 359758 64706 359760
rect 62113 359755 62179 359758
rect 41638 359484 41644 359548
rect 41708 359546 41714 359548
rect 41708 359486 41890 359546
rect 41708 359484 41714 359486
rect 41830 359277 41890 359486
rect 41781 359272 41890 359277
rect 41781 359216 41786 359272
rect 41842 359216 41890 359272
rect 41781 359214 41890 359216
rect 41781 359211 41847 359214
rect 64646 359146 64706 359758
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 663750 358670 676292 358730
rect 654777 358594 654843 358597
rect 663750 358594 663810 358670
rect 654777 358592 663810 358594
rect 654777 358536 654782 358592
rect 654838 358536 663810 358592
rect 654777 358534 663810 358536
rect 654777 358531 654843 358534
rect 675569 358322 675635 358325
rect 675569 358320 676292 358322
rect 675569 358264 675574 358320
rect 675630 358264 676292 358320
rect 675569 358262 676292 358264
rect 675569 358259 675635 358262
rect 62113 357778 62179 357781
rect 64646 357778 64706 357964
rect 675937 357914 676003 357917
rect 675937 357912 676292 357914
rect 675937 357856 675942 357912
rect 675998 357856 676292 357912
rect 675937 357854 676292 357856
rect 675937 357851 676003 357854
rect 62113 357776 64706 357778
rect 62113 357720 62118 357776
rect 62174 357720 64706 357776
rect 62113 357718 64706 357720
rect 62113 357715 62179 357718
rect 672809 357506 672875 357509
rect 672809 357504 676292 357506
rect 672809 357448 672814 357504
rect 672870 357448 676292 357504
rect 672809 357446 676292 357448
rect 672809 357443 672875 357446
rect 63401 357370 63467 357373
rect 63401 357368 64706 357370
rect 63401 357312 63406 357368
rect 63462 357312 64706 357368
rect 63401 357310 64706 357312
rect 63401 357307 63467 357310
rect 64646 356782 64706 357310
rect 672349 357098 672415 357101
rect 672349 357096 676292 357098
rect 672349 357040 672354 357096
rect 672410 357040 676292 357096
rect 672349 357038 676292 357040
rect 672349 357035 672415 357038
rect 673177 356826 673243 356829
rect 673177 356824 676230 356826
rect 673177 356768 673182 356824
rect 673238 356768 676230 356824
rect 673177 356766 676230 356768
rect 673177 356763 673243 356766
rect 652017 356690 652083 356693
rect 676170 356690 676230 356766
rect 652017 356688 663810 356690
rect 652017 356632 652022 356688
rect 652078 356632 663810 356688
rect 652017 356630 663810 356632
rect 676170 356630 676292 356690
rect 652017 356627 652083 356630
rect 663750 356554 663810 356630
rect 675937 356554 676003 356557
rect 663750 356552 676003 356554
rect 663750 356496 675942 356552
rect 675998 356496 676003 356552
rect 663750 356494 676003 356496
rect 675937 356491 676003 356494
rect 672533 356282 672599 356285
rect 672533 356280 676292 356282
rect 672533 356224 672538 356280
rect 672594 356224 676292 356280
rect 672533 356222 676292 356224
rect 672533 356219 672599 356222
rect 40534 356084 40540 356148
rect 40604 356146 40610 356148
rect 41781 356146 41847 356149
rect 40604 356144 41847 356146
rect 40604 356088 41786 356144
rect 41842 356088 41847 356144
rect 40604 356086 41847 356088
rect 40604 356084 40610 356086
rect 41781 356083 41847 356086
rect 61377 356010 61443 356013
rect 61377 356008 64706 356010
rect 61377 355952 61382 356008
rect 61438 355952 64706 356008
rect 61377 355950 64706 355952
rect 61377 355947 61443 355950
rect 64646 355600 64706 355950
rect 673361 355874 673427 355877
rect 673361 355872 676292 355874
rect 673361 355816 673366 355872
rect 673422 355816 676292 355872
rect 673361 355814 676292 355816
rect 673361 355811 673427 355814
rect 672165 355466 672231 355469
rect 672165 355464 676292 355466
rect 672165 355408 672170 355464
rect 672226 355408 676292 355464
rect 672165 355406 676292 355408
rect 672165 355403 672231 355406
rect 43805 355194 43871 355197
rect 44817 355194 44883 355197
rect 43805 355192 44883 355194
rect 43805 355136 43810 355192
rect 43866 355136 44822 355192
rect 44878 355136 44883 355192
rect 43805 355134 44883 355136
rect 43805 355131 43871 355134
rect 44817 355131 44883 355134
rect 673913 355058 673979 355061
rect 673913 355056 676292 355058
rect 673913 355000 673918 355056
rect 673974 355000 676292 355056
rect 673913 354998 676292 355000
rect 673913 354995 673979 354998
rect 43621 354922 43687 354925
rect 44633 354922 44699 354925
rect 43621 354920 44699 354922
rect 43621 354864 43626 354920
rect 43682 354864 44638 354920
rect 44694 354864 44699 354920
rect 43621 354862 44699 354864
rect 43621 354859 43687 354862
rect 44633 354859 44699 354862
rect 674097 354650 674163 354653
rect 674097 354648 676292 354650
rect 674097 354592 674102 354648
rect 674158 354592 676292 354648
rect 674097 354590 676292 354592
rect 674097 354587 674163 354590
rect 62941 354514 63007 354517
rect 62941 354512 64706 354514
rect 62941 354456 62946 354512
rect 63002 354456 64706 354512
rect 62941 354454 64706 354456
rect 62941 354451 63007 354454
rect 64646 354418 64706 354454
rect 42425 354378 42491 354381
rect 47117 354378 47183 354381
rect 42425 354376 47183 354378
rect 42425 354320 42430 354376
rect 42486 354320 47122 354376
rect 47178 354320 47183 354376
rect 42425 354318 47183 354320
rect 42425 354315 42491 354318
rect 47117 354315 47183 354318
rect 674741 354242 674807 354245
rect 674741 354240 676292 354242
rect 674741 354184 674746 354240
rect 674802 354184 676292 354240
rect 674741 354182 676292 354184
rect 674741 354179 674807 354182
rect 43069 353970 43135 353973
rect 45829 353970 45895 353973
rect 43069 353968 45895 353970
rect 43069 353912 43074 353968
rect 43130 353912 45834 353968
rect 45890 353912 45895 353968
rect 43069 353910 45895 353912
rect 43069 353907 43135 353910
rect 45829 353907 45895 353910
rect 675845 353834 675911 353837
rect 675845 353832 676292 353834
rect 675845 353776 675850 353832
rect 675906 353776 676292 353832
rect 675845 353774 676292 353776
rect 675845 353771 675911 353774
rect 43253 353698 43319 353701
rect 45829 353698 45895 353701
rect 43253 353696 45895 353698
rect 43253 353640 43258 353696
rect 43314 353640 45834 353696
rect 45890 353640 45895 353696
rect 43253 353638 45895 353640
rect 43253 353635 43319 353638
rect 45829 353635 45895 353638
rect 675518 353364 675524 353428
rect 675588 353426 675594 353428
rect 675588 353366 676292 353426
rect 675588 353364 675594 353366
rect 42149 353290 42215 353293
rect 51717 353290 51783 353293
rect 42149 353288 51783 353290
rect 42149 353232 42154 353288
rect 42210 353232 51722 353288
rect 51778 353232 51783 353288
rect 42149 353230 51783 353232
rect 42149 353227 42215 353230
rect 51717 353227 51783 353230
rect 42333 353018 42399 353021
rect 46933 353018 46999 353021
rect 42333 353016 46999 353018
rect 42333 352960 42338 353016
rect 42394 352960 46938 353016
rect 46994 352960 46999 353016
rect 42333 352958 46999 352960
rect 42333 352955 42399 352958
rect 46933 352955 46999 352958
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 675569 352882 675635 352885
rect 669270 352880 675635 352882
rect 669270 352824 675574 352880
rect 675630 352824 675635 352880
rect 669270 352822 675635 352824
rect 652385 352610 652451 352613
rect 669270 352610 669330 352822
rect 675569 352819 675635 352822
rect 652385 352608 669330 352610
rect 652385 352552 652390 352608
rect 652446 352552 669330 352608
rect 652385 352550 669330 352552
rect 673729 352610 673795 352613
rect 673729 352608 676292 352610
rect 673729 352552 673734 352608
rect 673790 352552 676292 352608
rect 673729 352550 676292 352552
rect 652385 352547 652451 352550
rect 673729 352547 673795 352550
rect 675932 352140 675938 352204
rect 676002 352202 676008 352204
rect 676002 352142 676292 352202
rect 676002 352140 676008 352142
rect 675845 351932 675911 351933
rect 675845 351930 675892 351932
rect 675800 351928 675892 351930
rect 675800 351872 675850 351928
rect 675800 351870 675892 351872
rect 675845 351868 675892 351870
rect 675956 351868 675962 351932
rect 675845 351867 675911 351868
rect 676029 351794 676095 351797
rect 676029 351792 676292 351794
rect 676029 351736 676034 351792
rect 676090 351736 676292 351792
rect 676029 351734 676292 351736
rect 676029 351731 676095 351734
rect 672993 351386 673059 351389
rect 672993 351384 676292 351386
rect 672993 351328 672998 351384
rect 673054 351328 676292 351384
rect 672993 351326 676292 351328
rect 672993 351323 673059 351326
rect 674281 350978 674347 350981
rect 674281 350976 676292 350978
rect 674281 350920 674286 350976
rect 674342 350920 676292 350976
rect 674281 350918 676292 350920
rect 674281 350915 674347 350918
rect 674557 350570 674623 350573
rect 674557 350568 676292 350570
rect 674557 350512 674562 350568
rect 674618 350512 676292 350568
rect 674557 350510 676292 350512
rect 674557 350507 674623 350510
rect 671981 350162 672047 350165
rect 671981 350160 676292 350162
rect 671981 350104 671986 350160
rect 672042 350104 676292 350160
rect 671981 350102 676292 350104
rect 671981 350099 672047 350102
rect 673361 349754 673427 349757
rect 673361 349752 676292 349754
rect 673361 349696 673366 349752
rect 673422 349696 676292 349752
rect 673361 349694 676292 349696
rect 673361 349691 673427 349694
rect 673545 349346 673611 349349
rect 673545 349344 676292 349346
rect 673545 349288 673550 349344
rect 673606 349288 676292 349344
rect 673545 349286 676292 349288
rect 673545 349283 673611 349286
rect 673913 348938 673979 348941
rect 673913 348936 676292 348938
rect 673913 348880 673918 348936
rect 673974 348880 676292 348936
rect 673913 348878 676292 348880
rect 673913 348875 673979 348878
rect 672717 348530 672783 348533
rect 672717 348528 676292 348530
rect 672717 348472 672722 348528
rect 672778 348472 676292 348528
rect 672717 348470 676292 348472
rect 672717 348467 672783 348470
rect 683070 347717 683130 348092
rect 683070 347712 683179 347717
rect 683070 347684 683118 347712
rect 683100 347656 683118 347684
rect 683174 347656 683179 347712
rect 683100 347654 683179 347656
rect 683113 347651 683179 347654
rect 676029 347306 676095 347309
rect 676029 347304 676292 347306
rect 676029 347248 676034 347304
rect 676090 347248 676292 347304
rect 676029 347246 676292 347248
rect 676029 347243 676095 347246
rect 658917 346490 658983 346493
rect 676262 346490 676322 346868
rect 676489 346628 676555 346629
rect 676438 346564 676444 346628
rect 676508 346626 676555 346628
rect 676508 346624 676600 346626
rect 676550 346568 676600 346624
rect 676508 346566 676600 346568
rect 676508 346564 676555 346566
rect 676489 346563 676555 346564
rect 683113 346490 683179 346493
rect 658917 346488 676322 346490
rect 658917 346432 658922 346488
rect 658978 346432 676322 346488
rect 658917 346430 676322 346432
rect 676814 346488 683179 346490
rect 676814 346432 683118 346488
rect 683174 346432 683179 346488
rect 676814 346430 683179 346432
rect 658917 346427 658983 346430
rect 676814 346220 676874 346430
rect 683113 346427 683179 346430
rect 676806 346156 676812 346220
rect 676876 346156 676882 346220
rect 669957 345674 670023 345677
rect 676029 345674 676095 345677
rect 669957 345672 676095 345674
rect 669957 345616 669962 345672
rect 670018 345616 676034 345672
rect 676090 345616 676095 345672
rect 669957 345614 676095 345616
rect 669957 345611 670023 345614
rect 676029 345611 676095 345614
rect 35758 344317 35818 344556
rect 35758 344312 35867 344317
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35758 344254 35867 344256
rect 35801 344251 35867 344254
rect 35574 343909 35634 344148
rect 35574 343904 35683 343909
rect 35574 343848 35622 343904
rect 35678 343848 35683 343904
rect 35574 343846 35683 343848
rect 35617 343843 35683 343846
rect 40401 343906 40467 343909
rect 46013 343906 46079 343909
rect 40401 343904 46079 343906
rect 40401 343848 40406 343904
rect 40462 343848 46018 343904
rect 46074 343848 46079 343904
rect 40401 343846 46079 343848
rect 40401 343843 40467 343846
rect 46013 343843 46079 343846
rect 35758 343501 35818 343740
rect 35758 343496 35867 343501
rect 35758 343440 35806 343496
rect 35862 343440 35867 343496
rect 35758 343438 35867 343440
rect 35801 343435 35867 343438
rect 45185 343362 45251 343365
rect 41492 343360 45251 343362
rect 41492 343304 45190 343360
rect 45246 343304 45251 343360
rect 41492 343302 45251 343304
rect 45185 343299 45251 343302
rect 44398 342954 44404 342956
rect 41492 342894 44404 342954
rect 44398 342892 44404 342894
rect 44468 342892 44474 342956
rect 45001 342546 45067 342549
rect 41492 342544 45067 342546
rect 41492 342488 45006 342544
rect 45062 342488 45067 342544
rect 41492 342486 45067 342488
rect 45001 342483 45067 342486
rect 40217 342274 40283 342277
rect 45461 342274 45527 342277
rect 40217 342272 45527 342274
rect 40217 342216 40222 342272
rect 40278 342216 45466 342272
rect 45522 342216 45527 342272
rect 40217 342214 45527 342216
rect 40217 342211 40283 342214
rect 45461 342211 45527 342214
rect 39622 341869 39682 342108
rect 35801 341866 35867 341869
rect 35758 341864 35867 341866
rect 35758 341808 35806 341864
rect 35862 341808 35867 341864
rect 35758 341803 35867 341808
rect 39622 341864 39731 341869
rect 39622 341808 39670 341864
rect 39726 341808 39731 341864
rect 39622 341806 39731 341808
rect 39665 341803 39731 341806
rect 39849 341866 39915 341869
rect 39849 341864 45570 341866
rect 39849 341808 39854 341864
rect 39910 341808 45570 341864
rect 39849 341806 45570 341808
rect 39849 341803 39915 341806
rect 35758 341700 35818 341803
rect 45510 341730 45570 341806
rect 62941 341730 63007 341733
rect 45510 341728 63007 341730
rect 45510 341672 62946 341728
rect 63002 341672 63007 341728
rect 45510 341670 63007 341672
rect 62941 341667 63007 341670
rect 44214 341594 44220 341596
rect 42014 341534 44220 341594
rect 42014 341322 42074 341534
rect 44214 341532 44220 341534
rect 44284 341532 44290 341596
rect 62757 341458 62823 341461
rect 45510 341456 62823 341458
rect 45510 341400 62762 341456
rect 62818 341400 62823 341456
rect 45510 341398 62823 341400
rect 41492 341262 42074 341322
rect 42241 341322 42307 341325
rect 45510 341322 45570 341398
rect 62757 341395 62823 341398
rect 42241 341320 45570 341322
rect 42241 341264 42246 341320
rect 42302 341264 45570 341320
rect 42241 341262 45570 341264
rect 42241 341259 42307 341262
rect 35801 341050 35867 341053
rect 35758 341048 35867 341050
rect 35758 340992 35806 341048
rect 35862 340992 35867 341048
rect 35758 340987 35867 340992
rect 40125 341050 40191 341053
rect 40125 341048 40418 341050
rect 40125 340992 40130 341048
rect 40186 340992 40418 341048
rect 40125 340990 40418 340992
rect 40125 340987 40191 340990
rect 35758 340884 35818 340987
rect 40358 340778 40418 340990
rect 45645 340778 45711 340781
rect 675569 340780 675635 340781
rect 675518 340778 675524 340780
rect 40358 340776 45711 340778
rect 40358 340720 45650 340776
rect 45706 340720 45711 340776
rect 40358 340718 45711 340720
rect 675478 340718 675524 340778
rect 675588 340776 675635 340780
rect 675630 340720 675635 340776
rect 45645 340715 45711 340718
rect 675518 340716 675524 340718
rect 675588 340716 675635 340720
rect 675569 340715 675635 340716
rect 42742 340506 42748 340508
rect 41492 340446 42748 340506
rect 42742 340444 42748 340446
rect 42812 340444 42818 340508
rect 39665 340234 39731 340237
rect 44582 340234 44588 340236
rect 39665 340232 44588 340234
rect 39665 340176 39670 340232
rect 39726 340176 44588 340232
rect 39665 340174 44588 340176
rect 39665 340171 39731 340174
rect 44582 340172 44588 340174
rect 44652 340172 44658 340236
rect 675753 340234 675819 340237
rect 676438 340234 676444 340236
rect 675753 340232 676444 340234
rect 675753 340176 675758 340232
rect 675814 340176 676444 340232
rect 675753 340174 676444 340176
rect 675753 340171 675819 340174
rect 676438 340172 676444 340174
rect 676508 340172 676514 340236
rect 35574 339829 35634 340068
rect 35525 339824 35634 339829
rect 35801 339826 35867 339829
rect 35525 339768 35530 339824
rect 35586 339768 35634 339824
rect 35525 339766 35634 339768
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35525 339763 35591 339766
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 46933 339282 46999 339285
rect 41492 339280 46999 339282
rect 41492 339224 46938 339280
rect 46994 339224 46999 339280
rect 41492 339222 46999 339224
rect 46933 339219 46999 339222
rect 45553 338874 45619 338877
rect 41492 338872 45619 338874
rect 41492 338816 45558 338872
rect 45614 338816 45619 338872
rect 41492 338814 45619 338816
rect 45553 338811 45619 338814
rect 653397 338738 653463 338741
rect 675109 338738 675175 338741
rect 653397 338736 675175 338738
rect 653397 338680 653402 338736
rect 653458 338680 675114 338736
rect 675170 338680 675175 338736
rect 653397 338678 675175 338680
rect 653397 338675 653463 338678
rect 675109 338675 675175 338678
rect 41462 338194 41522 338436
rect 41638 338194 41644 338196
rect 41462 338134 41644 338194
rect 41638 338132 41644 338134
rect 41708 338132 41714 338196
rect 41278 337922 41338 338028
rect 45369 337922 45435 337925
rect 41278 337920 45435 337922
rect 41278 337864 45374 337920
rect 45430 337864 45435 337920
rect 41278 337862 45435 337864
rect 45369 337859 45435 337862
rect 675661 337786 675727 337789
rect 675886 337786 675892 337788
rect 675661 337784 675892 337786
rect 675661 337728 675666 337784
rect 675722 337728 675892 337784
rect 675661 337726 675892 337728
rect 675661 337723 675727 337726
rect 675886 337724 675892 337726
rect 675956 337724 675962 337788
rect 42926 337650 42932 337652
rect 41492 337590 42932 337650
rect 42926 337588 42932 337590
rect 42996 337588 43002 337652
rect 43110 337242 43116 337244
rect 41492 337182 43116 337242
rect 43110 337180 43116 337182
rect 43180 337180 43186 337244
rect 672993 337242 673059 337245
rect 675109 337242 675175 337245
rect 672993 337240 675175 337242
rect 672993 337184 672998 337240
rect 673054 337184 675114 337240
rect 675170 337184 675175 337240
rect 672993 337182 675175 337184
rect 672993 337179 673059 337182
rect 675109 337179 675175 337182
rect 40718 336908 40724 336972
rect 40788 336908 40794 336972
rect 40726 336804 40786 336908
rect 37089 336562 37155 336565
rect 42006 336562 42012 336564
rect 37089 336560 42012 336562
rect 37089 336504 37094 336560
rect 37150 336504 42012 336560
rect 37089 336502 42012 336504
rect 37089 336499 37155 336502
rect 42006 336500 42012 336502
rect 42076 336500 42082 336564
rect 41462 336154 41522 336396
rect 41462 336094 44466 336154
rect 35758 335749 35818 335988
rect 35758 335744 35867 335749
rect 35758 335688 35806 335744
rect 35862 335688 35867 335744
rect 35758 335686 35867 335688
rect 35801 335683 35867 335686
rect 38837 335746 38903 335749
rect 41822 335746 41828 335748
rect 38837 335744 41828 335746
rect 38837 335688 38842 335744
rect 38898 335688 41828 335744
rect 38837 335686 41828 335688
rect 38837 335683 38903 335686
rect 41822 335684 41828 335686
rect 41892 335684 41898 335748
rect 40542 335340 40602 335580
rect 40534 335276 40540 335340
rect 40604 335276 40610 335340
rect 41462 334930 41522 335172
rect 41462 334870 41890 334930
rect 35758 334525 35818 334764
rect 41830 334658 41890 334870
rect 44406 334661 44466 336094
rect 673361 335610 673427 335613
rect 675109 335610 675175 335613
rect 673361 335608 675175 335610
rect 673361 335552 673366 335608
rect 673422 335552 675114 335608
rect 675170 335552 675175 335608
rect 673361 335550 675175 335552
rect 673361 335547 673427 335550
rect 675109 335547 675175 335550
rect 44173 334658 44239 334661
rect 41830 334656 44239 334658
rect 41830 334600 44178 334656
rect 44234 334600 44239 334656
rect 41830 334598 44239 334600
rect 44173 334595 44239 334598
rect 44357 334656 44466 334661
rect 44357 334600 44362 334656
rect 44418 334600 44466 334656
rect 44357 334598 44466 334600
rect 44357 334595 44423 334598
rect 35758 334520 35867 334525
rect 35758 334464 35806 334520
rect 35862 334464 35867 334520
rect 35758 334462 35867 334464
rect 35801 334459 35867 334462
rect 41462 334114 41522 334356
rect 51717 334114 51783 334117
rect 41462 334112 51783 334114
rect 41462 334056 51722 334112
rect 51778 334056 51783 334112
rect 41462 334054 51783 334056
rect 51717 334051 51783 334054
rect 673729 333978 673795 333981
rect 675109 333978 675175 333981
rect 673729 333976 675175 333978
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 673729 333920 673734 333976
rect 673790 333920 675114 333976
rect 675170 333920 675175 333976
rect 673729 333918 675175 333920
rect 673729 333915 673795 333918
rect 675109 333915 675175 333918
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 50337 333162 50403 333165
rect 41492 333160 50403 333162
rect 41492 333104 50342 333160
rect 50398 333104 50403 333160
rect 41492 333102 50403 333104
rect 50337 333099 50403 333102
rect 40309 332890 40375 332893
rect 42885 332890 42951 332893
rect 40309 332888 42951 332890
rect 40309 332832 40314 332888
rect 40370 332832 42890 332888
rect 42946 332832 42951 332888
rect 40309 332830 42951 332832
rect 40309 332827 40375 332830
rect 42885 332827 42951 332830
rect 673545 332754 673611 332757
rect 675109 332754 675175 332757
rect 673545 332752 675175 332754
rect 673545 332696 673550 332752
rect 673606 332696 675114 332752
rect 675170 332696 675175 332752
rect 673545 332694 675175 332696
rect 673545 332691 673611 332694
rect 675109 332691 675175 332694
rect 39849 332482 39915 332485
rect 43069 332482 43135 332485
rect 39849 332480 43135 332482
rect 39849 332424 39854 332480
rect 39910 332424 43074 332480
rect 43130 332424 43135 332480
rect 39849 332422 43135 332424
rect 39849 332419 39915 332422
rect 43069 332419 43135 332422
rect 671981 332346 672047 332349
rect 675109 332346 675175 332349
rect 671981 332344 675175 332346
rect 671981 332288 671986 332344
rect 672042 332288 675114 332344
rect 675170 332288 675175 332344
rect 671981 332286 675175 332288
rect 671981 332283 672047 332286
rect 675109 332283 675175 332286
rect 673913 331258 673979 331261
rect 675109 331258 675175 331261
rect 673913 331256 675175 331258
rect 673913 331200 673918 331256
rect 673974 331200 675114 331256
rect 675170 331200 675175 331256
rect 673913 331198 675175 331200
rect 673913 331195 673979 331198
rect 675109 331195 675175 331198
rect 652385 329762 652451 329765
rect 649950 329760 652451 329762
rect 649950 329704 652390 329760
rect 652446 329704 652451 329760
rect 649950 329702 652451 329704
rect 649950 329234 650010 329702
rect 652385 329699 652451 329702
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 651373 328130 651439 328133
rect 649950 328128 651439 328130
rect 649950 328072 651378 328128
rect 651434 328072 651439 328128
rect 649950 328070 651439 328072
rect 649950 328052 650010 328070
rect 651373 328067 651439 328070
rect 42425 327042 42491 327045
rect 45277 327042 45343 327045
rect 42425 327040 45343 327042
rect 42425 326984 42430 327040
rect 42486 326984 45282 327040
rect 45338 326984 45343 327040
rect 42425 326982 45343 326984
rect 42425 326979 42491 326982
rect 45277 326979 45343 326982
rect 652017 326906 652083 326909
rect 650502 326904 652083 326906
rect 650502 326900 652022 326904
rect 649980 326848 652022 326900
rect 652078 326848 652083 326904
rect 649980 326846 652083 326848
rect 649980 326840 650562 326846
rect 652017 326843 652083 326846
rect 649950 325682 650010 325710
rect 651373 325682 651439 325685
rect 649950 325680 651439 325682
rect 649950 325624 651378 325680
rect 651434 325624 651439 325680
rect 649950 325622 651439 325624
rect 651373 325619 651439 325622
rect 675293 325546 675359 325549
rect 676254 325546 676260 325548
rect 675293 325544 676260 325546
rect 675293 325488 675298 325544
rect 675354 325488 676260 325544
rect 675293 325486 676260 325488
rect 675293 325483 675359 325486
rect 676254 325484 676260 325486
rect 676324 325484 676330 325548
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 675109 325274 675175 325277
rect 676806 325274 676812 325276
rect 675109 325272 676812 325274
rect 675109 325216 675114 325272
rect 675170 325216 676812 325272
rect 675109 325214 676812 325216
rect 675109 325211 675175 325214
rect 676806 325212 676812 325214
rect 676876 325212 676882 325276
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 42057 322826 42123 322829
rect 44357 322826 44423 322829
rect 42057 322824 44423 322826
rect 42057 322768 42062 322824
rect 42118 322768 44362 322824
rect 44418 322768 44423 322824
rect 42057 322766 44423 322768
rect 42057 322763 42123 322766
rect 44357 322763 44423 322766
rect 42057 321194 42123 321197
rect 42885 321194 42951 321197
rect 42057 321192 42951 321194
rect 42057 321136 42062 321192
rect 42118 321136 42890 321192
rect 42946 321136 42951 321192
rect 42057 321134 42951 321136
rect 42057 321131 42123 321134
rect 42885 321131 42951 321134
rect 42609 320786 42675 320789
rect 53833 320786 53899 320789
rect 42609 320784 53899 320786
rect 42609 320728 42614 320784
rect 42670 320728 53838 320784
rect 53894 320728 53899 320784
rect 42609 320726 53899 320728
rect 42609 320723 42675 320726
rect 53833 320723 53899 320726
rect 42149 320514 42215 320517
rect 43069 320514 43135 320517
rect 42149 320512 43135 320514
rect 42149 320456 42154 320512
rect 42210 320456 43074 320512
rect 43130 320456 43135 320512
rect 42149 320454 43135 320456
rect 42149 320451 42215 320454
rect 43069 320451 43135 320454
rect 41873 319972 41939 319973
rect 41822 319970 41828 319972
rect 41782 319910 41828 319970
rect 41892 319968 41939 319972
rect 41934 319912 41939 319968
rect 41822 319908 41828 319910
rect 41892 319908 41939 319912
rect 41873 319907 41939 319908
rect 42057 319970 42123 319973
rect 44173 319970 44239 319973
rect 42057 319968 44239 319970
rect 42057 319912 42062 319968
rect 42118 319912 44178 319968
rect 44234 319912 44239 319968
rect 42057 319910 44239 319912
rect 42057 319907 42123 319910
rect 44173 319907 44239 319910
rect 42425 319698 42491 319701
rect 53097 319698 53163 319701
rect 42425 319696 53163 319698
rect 42425 319640 42430 319696
rect 42486 319640 53102 319696
rect 53158 319640 53163 319696
rect 42425 319638 53163 319640
rect 42425 319635 42491 319638
rect 53097 319635 53163 319638
rect 40718 318956 40724 319020
rect 40788 319018 40794 319020
rect 42241 319018 42307 319021
rect 40788 319016 42307 319018
rect 40788 318960 42246 319016
rect 42302 318960 42307 319016
rect 40788 318958 42307 318960
rect 40788 318956 40794 318958
rect 42241 318955 42307 318958
rect 40534 317324 40540 317388
rect 40604 317386 40610 317388
rect 41781 317386 41847 317389
rect 40604 317384 41847 317386
rect 40604 317328 41786 317384
rect 41842 317328 41847 317384
rect 40604 317326 41847 317328
rect 40604 317324 40610 317326
rect 41781 317323 41847 317326
rect 62113 317386 62179 317389
rect 62113 317384 64706 317386
rect 62113 317328 62118 317384
rect 62174 317328 64706 317384
rect 62113 317326 64706 317328
rect 62113 317323 62179 317326
rect 64646 317106 64706 317326
rect 42149 316026 42215 316029
rect 43110 316026 43116 316028
rect 42149 316024 43116 316026
rect 42149 315968 42154 316024
rect 42210 315968 43116 316024
rect 42149 315966 43116 315968
rect 42149 315963 42215 315966
rect 43110 315964 43116 315966
rect 43180 315964 43186 316028
rect 62113 316026 62179 316029
rect 62113 316024 64706 316026
rect 62113 315968 62118 316024
rect 62174 315968 64706 316024
rect 62113 315966 64706 315968
rect 62113 315963 62179 315966
rect 64646 315924 64706 315966
rect 42149 315482 42215 315485
rect 45553 315482 45619 315485
rect 42149 315480 45619 315482
rect 42149 315424 42154 315480
rect 42210 315424 45558 315480
rect 45614 315424 45619 315480
rect 42149 315422 45619 315424
rect 42149 315419 42215 315422
rect 45553 315419 45619 315422
rect 62113 314802 62179 314805
rect 62113 314800 64706 314802
rect 62113 314744 62118 314800
rect 62174 314744 64706 314800
rect 62113 314742 64706 314744
rect 62113 314739 62179 314742
rect 63125 314122 63191 314125
rect 63125 314120 64706 314122
rect 63125 314064 63130 314120
rect 63186 314064 64706 314120
rect 63125 314062 64706 314064
rect 63125 314059 63191 314062
rect 42057 313716 42123 313717
rect 42006 313714 42012 313716
rect 41966 313654 42012 313714
rect 42076 313712 42123 313716
rect 42118 313656 42123 313712
rect 42006 313652 42012 313654
rect 42076 313652 42123 313656
rect 42057 313651 42123 313652
rect 64646 313560 64706 314062
rect 676213 313986 676279 313989
rect 676213 313984 676322 313986
rect 676213 313928 676218 313984
rect 676274 313928 676322 313984
rect 676213 313923 676322 313928
rect 676262 313684 676322 313923
rect 653397 313306 653463 313309
rect 653397 313304 676292 313306
rect 653397 313248 653402 313304
rect 653458 313248 676292 313304
rect 653397 313246 676292 313248
rect 653397 313243 653463 313246
rect 62941 313034 63007 313037
rect 674649 313034 674715 313037
rect 62941 313032 64706 313034
rect 62941 312976 62946 313032
rect 63002 312976 64706 313032
rect 62941 312974 64706 312976
rect 62941 312971 63007 312974
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 64646 312378 64706 312974
rect 674649 313032 675034 313034
rect 674649 312976 674654 313032
rect 674710 312976 675034 313032
rect 674649 312974 675034 312976
rect 674649 312971 674715 312974
rect 674974 312898 675034 312974
rect 674974 312838 676292 312898
rect 673361 312762 673427 312765
rect 674833 312762 674899 312765
rect 673361 312760 674899 312762
rect 673361 312704 673366 312760
rect 673422 312704 674838 312760
rect 674894 312704 674899 312760
rect 673361 312702 674899 312704
rect 673361 312699 673427 312702
rect 674833 312699 674899 312702
rect 672349 312490 672415 312493
rect 672349 312488 676292 312490
rect 672349 312432 672354 312488
rect 672410 312432 676292 312488
rect 672349 312430 676292 312432
rect 672349 312427 672415 312430
rect 674833 312082 674899 312085
rect 674833 312080 676292 312082
rect 674833 312024 674838 312080
rect 674894 312024 676292 312080
rect 674833 312022 676292 312024
rect 674833 312019 674899 312022
rect 664437 311946 664503 311949
rect 674649 311946 674715 311949
rect 664437 311944 674715 311946
rect 664437 311888 664442 311944
rect 664498 311888 674654 311944
rect 674710 311888 674715 311944
rect 664437 311886 674715 311888
rect 664437 311883 664503 311886
rect 674649 311883 674715 311886
rect 62757 311810 62823 311813
rect 62757 311808 64706 311810
rect 62757 311752 62762 311808
rect 62818 311752 64706 311808
rect 62757 311750 64706 311752
rect 62757 311747 62823 311750
rect 64646 311196 64706 311750
rect 672533 311674 672599 311677
rect 672533 311672 676292 311674
rect 672533 311616 672538 311672
rect 672594 311616 676292 311672
rect 672533 311614 676292 311616
rect 672533 311611 672599 311614
rect 673177 311266 673243 311269
rect 673177 311264 676292 311266
rect 673177 311208 673182 311264
rect 673238 311208 676292 311264
rect 673177 311206 676292 311208
rect 673177 311203 673243 311206
rect 672165 310858 672231 310861
rect 672165 310856 676292 310858
rect 672165 310800 672170 310856
rect 672226 310800 676292 310856
rect 672165 310798 676292 310800
rect 672165 310795 672231 310798
rect 42425 310450 42491 310453
rect 46933 310450 46999 310453
rect 42425 310448 46999 310450
rect 42425 310392 42430 310448
rect 42486 310392 46938 310448
rect 46994 310392 46999 310448
rect 42425 310390 46999 310392
rect 42425 310387 42491 310390
rect 46933 310387 46999 310390
rect 674189 310450 674255 310453
rect 674189 310448 676292 310450
rect 674189 310392 674194 310448
rect 674250 310392 676292 310448
rect 674189 310390 676292 310392
rect 674189 310387 674255 310390
rect 674373 310042 674439 310045
rect 674373 310040 676292 310042
rect 674373 309984 674378 310040
rect 674434 309984 676292 310040
rect 674373 309982 676292 309984
rect 674373 309979 674439 309982
rect 652293 309906 652359 309909
rect 652293 309904 663810 309906
rect 652293 309848 652298 309904
rect 652354 309848 663810 309904
rect 652293 309846 663810 309848
rect 652293 309843 652359 309846
rect 663750 309362 663810 309846
rect 674557 309634 674623 309637
rect 674557 309632 676292 309634
rect 674557 309576 674562 309632
rect 674618 309576 676292 309632
rect 674557 309574 676292 309576
rect 674557 309571 674623 309574
rect 675845 309362 675911 309365
rect 663750 309360 675911 309362
rect 663750 309304 675850 309360
rect 675906 309304 675911 309360
rect 663750 309302 675911 309304
rect 675845 309299 675911 309302
rect 676032 309166 676292 309226
rect 42057 309090 42123 309093
rect 59905 309090 59971 309093
rect 42057 309088 59971 309090
rect 42057 309032 42062 309088
rect 42118 309032 59910 309088
rect 59966 309032 59971 309088
rect 42057 309030 59971 309032
rect 42057 309027 42123 309030
rect 59905 309027 59971 309030
rect 675702 309028 675708 309092
rect 675772 309090 675778 309092
rect 676032 309090 676092 309166
rect 675772 309030 676092 309090
rect 675772 309028 675778 309030
rect 675702 308756 675708 308820
rect 675772 308818 675778 308820
rect 675772 308758 676292 308818
rect 675772 308756 675778 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675109 308002 675175 308005
rect 675109 308000 676292 308002
rect 675109 307944 675114 308000
rect 675170 307944 676292 308000
rect 675109 307942 676292 307944
rect 675109 307939 675175 307942
rect 676029 307594 676095 307597
rect 676029 307592 676292 307594
rect 676029 307536 676034 307592
rect 676090 307536 676292 307592
rect 676029 307534 676292 307536
rect 676029 307531 676095 307534
rect 675886 307124 675892 307188
rect 675956 307186 675962 307188
rect 675956 307126 676292 307186
rect 675956 307124 675962 307126
rect 679617 306778 679683 306781
rect 679604 306776 679683 306778
rect 679604 306720 679622 306776
rect 679678 306720 679683 306776
rect 679604 306718 679683 306720
rect 679617 306715 679683 306718
rect 677593 306370 677659 306373
rect 677580 306368 677659 306370
rect 677580 306312 677598 306368
rect 677654 306312 677659 306368
rect 677580 306310 677659 306312
rect 677593 306307 677659 306310
rect 676489 305962 676555 305965
rect 676476 305960 676555 305962
rect 676476 305904 676494 305960
rect 676550 305904 676555 305960
rect 676476 305902 676555 305904
rect 676489 305899 676555 305902
rect 672993 305554 673059 305557
rect 672993 305552 676292 305554
rect 672993 305496 672998 305552
rect 673054 305496 676292 305552
rect 672993 305494 676292 305496
rect 672993 305491 673059 305494
rect 674373 305146 674439 305149
rect 674373 305144 676292 305146
rect 674373 305088 674378 305144
rect 674434 305088 676292 305144
rect 674373 305086 676292 305088
rect 674373 305083 674439 305086
rect 676029 304738 676095 304741
rect 676029 304736 676292 304738
rect 676029 304680 676034 304736
rect 676090 304680 676292 304736
rect 676029 304678 676292 304680
rect 676029 304675 676095 304678
rect 672533 304330 672599 304333
rect 672533 304328 676292 304330
rect 672533 304272 672538 304328
rect 672594 304272 676292 304328
rect 672533 304270 676292 304272
rect 672533 304267 672599 304270
rect 674005 303922 674071 303925
rect 674005 303920 676292 303922
rect 674005 303864 674010 303920
rect 674066 303864 676292 303920
rect 674005 303862 676292 303864
rect 674005 303859 674071 303862
rect 673637 303514 673703 303517
rect 673637 303512 676292 303514
rect 673637 303456 673642 303512
rect 673698 303456 676292 303512
rect 673637 303454 676292 303456
rect 673637 303451 673703 303454
rect 651373 303378 651439 303381
rect 649950 303376 651439 303378
rect 649950 303320 651378 303376
rect 651434 303320 651439 303376
rect 649950 303318 651439 303320
rect 649950 302776 650010 303318
rect 651373 303315 651439 303318
rect 683070 302701 683130 303076
rect 683021 302696 683130 302701
rect 683021 302640 683026 302696
rect 683082 302668 683130 302696
rect 683082 302640 683100 302668
rect 683021 302638 683100 302640
rect 683021 302635 683087 302638
rect 671521 302290 671587 302293
rect 671521 302288 676292 302290
rect 671521 302232 671526 302288
rect 671582 302232 676292 302288
rect 671521 302230 676292 302232
rect 671521 302227 671587 302230
rect 652293 302154 652359 302157
rect 649950 302152 652359 302154
rect 649950 302096 652298 302152
rect 652354 302096 652359 302152
rect 649950 302094 652359 302096
rect 649950 301594 650010 302094
rect 652293 302091 652359 302094
rect 674925 301882 674991 301885
rect 675845 301882 675911 301885
rect 674925 301880 675911 301882
rect 674925 301824 674930 301880
rect 674986 301824 675850 301880
rect 675906 301824 675911 301880
rect 674925 301822 675911 301824
rect 674925 301819 674991 301822
rect 675845 301819 675911 301822
rect 53097 301338 53163 301341
rect 41492 301336 53163 301338
rect 41492 301280 53102 301336
rect 53158 301280 53163 301336
rect 41492 301278 53163 301280
rect 53097 301275 53163 301278
rect 35617 300930 35683 300933
rect 35604 300928 35683 300930
rect 35604 300872 35622 300928
rect 35678 300872 35683 300928
rect 35604 300870 35683 300872
rect 35617 300867 35683 300870
rect 654777 300930 654843 300933
rect 676262 300930 676322 301852
rect 676489 301612 676555 301613
rect 676438 301548 676444 301612
rect 676508 301610 676555 301612
rect 676508 301608 676600 301610
rect 676550 301552 676600 301608
rect 676508 301550 676600 301552
rect 676508 301548 676555 301550
rect 676489 301547 676555 301548
rect 654777 300928 676322 300930
rect 654777 300872 654782 300928
rect 654838 300872 676322 300928
rect 654777 300870 676322 300872
rect 654777 300867 654843 300870
rect 651465 300658 651531 300661
rect 649950 300656 651531 300658
rect 649950 300600 651470 300656
rect 651526 300600 651531 300656
rect 649950 300598 651531 300600
rect 46197 300522 46263 300525
rect 41492 300520 46263 300522
rect 41492 300464 46202 300520
rect 46258 300464 46263 300520
rect 41492 300462 46263 300464
rect 46197 300459 46263 300462
rect 649950 300412 650010 300598
rect 651465 300595 651531 300598
rect 676029 300658 676095 300661
rect 676254 300658 676260 300660
rect 676029 300656 676260 300658
rect 676029 300600 676034 300656
rect 676090 300600 676260 300656
rect 676029 300598 676260 300600
rect 676029 300595 676095 300598
rect 676254 300596 676260 300598
rect 676324 300596 676330 300660
rect 44398 300114 44404 300116
rect 41492 300054 44404 300114
rect 44398 300052 44404 300054
rect 44468 300052 44474 300116
rect 44173 299706 44239 299709
rect 41492 299704 44239 299706
rect 41492 299648 44178 299704
rect 44234 299648 44239 299704
rect 41492 299646 44239 299648
rect 44173 299643 44239 299646
rect 675702 299372 675708 299436
rect 675772 299434 675778 299436
rect 683021 299434 683087 299437
rect 675772 299432 683087 299434
rect 675772 299376 683026 299432
rect 683082 299376 683087 299432
rect 675772 299374 683087 299376
rect 675772 299372 675778 299374
rect 683021 299371 683087 299374
rect 44582 299298 44588 299300
rect 41492 299238 44588 299298
rect 44582 299236 44588 299238
rect 44652 299236 44658 299300
rect 35801 298890 35867 298893
rect 35788 298888 35867 298890
rect 35788 298832 35806 298888
rect 35862 298832 35867 298888
rect 35788 298830 35867 298832
rect 35801 298827 35867 298830
rect 41781 298754 41847 298757
rect 62757 298754 62823 298757
rect 41781 298752 62823 298754
rect 41781 298696 41786 298752
rect 41842 298696 62762 298752
rect 62818 298696 62823 298752
rect 41781 298694 62823 298696
rect 649950 298754 650010 299230
rect 651465 298754 651531 298757
rect 649950 298752 651531 298754
rect 649950 298696 651470 298752
rect 651526 298696 651531 298752
rect 649950 298694 651531 298696
rect 41781 298691 41847 298694
rect 62757 298691 62823 298694
rect 651465 298691 651531 298694
rect 44214 298482 44220 298484
rect 41492 298422 44220 298482
rect 44214 298420 44220 298422
rect 44284 298420 44290 298484
rect 45001 298074 45067 298077
rect 41492 298072 45067 298074
rect 41492 298016 45006 298072
rect 45062 298016 45067 298072
rect 41492 298014 45067 298016
rect 45001 298011 45067 298014
rect 42742 297666 42748 297668
rect 41492 297606 42748 297666
rect 42742 297604 42748 297606
rect 42812 297604 42818 297668
rect 649950 297530 650010 298048
rect 651465 297530 651531 297533
rect 649950 297528 651531 297530
rect 649950 297472 651470 297528
rect 651526 297472 651531 297528
rect 649950 297470 651531 297472
rect 651465 297467 651531 297470
rect 44357 297258 44423 297261
rect 41492 297256 44423 297258
rect 41492 297200 44362 297256
rect 44418 297200 44423 297256
rect 41492 297198 44423 297200
rect 44357 297195 44423 297198
rect 42006 296850 42012 296852
rect 41492 296790 42012 296850
rect 42006 296788 42012 296790
rect 42076 296788 42082 296852
rect 649950 296850 650010 296866
rect 652661 296850 652727 296853
rect 649950 296848 652727 296850
rect 649950 296792 652666 296848
rect 652722 296792 652727 296848
rect 649950 296790 652727 296792
rect 652661 296787 652727 296790
rect 675334 296788 675340 296852
rect 675404 296850 675410 296852
rect 676121 296850 676187 296853
rect 675404 296848 676187 296850
rect 675404 296792 676126 296848
rect 676182 296792 676187 296848
rect 675404 296790 676187 296792
rect 675404 296788 675410 296790
rect 676121 296787 676187 296790
rect 41781 296578 41847 296581
rect 42793 296578 42859 296581
rect 41781 296576 42859 296578
rect 41781 296520 41786 296576
rect 41842 296520 42798 296576
rect 42854 296520 42859 296576
rect 41781 296518 42859 296520
rect 41781 296515 41847 296518
rect 42793 296515 42859 296518
rect 675518 296516 675524 296580
rect 675588 296578 675594 296580
rect 675937 296578 676003 296581
rect 675588 296576 676003 296578
rect 675588 296520 675942 296576
rect 675998 296520 676003 296576
rect 675588 296518 676003 296520
rect 675588 296516 675594 296518
rect 675937 296515 676003 296518
rect 35433 296442 35499 296445
rect 35420 296440 35499 296442
rect 35420 296384 35438 296440
rect 35494 296384 35499 296440
rect 35420 296382 35499 296384
rect 35433 296379 35499 296382
rect 35617 296034 35683 296037
rect 35604 296032 35683 296034
rect 35604 295976 35622 296032
rect 35678 295976 35683 296032
rect 35604 295974 35683 295976
rect 35617 295971 35683 295974
rect 35801 295626 35867 295629
rect 35788 295624 35867 295626
rect 35788 295568 35806 295624
rect 35862 295568 35867 295624
rect 35788 295566 35867 295568
rect 35801 295563 35867 295566
rect 62113 295490 62179 295493
rect 64646 295490 64706 295684
rect 62113 295488 64706 295490
rect 62113 295432 62118 295488
rect 62174 295432 64706 295488
rect 62113 295430 64706 295432
rect 62113 295427 62179 295430
rect 41781 295354 41847 295357
rect 43161 295354 43227 295357
rect 41781 295352 43227 295354
rect 41781 295296 41786 295352
rect 41842 295296 43166 295352
rect 43222 295296 43227 295352
rect 41781 295294 43227 295296
rect 649950 295354 650010 295684
rect 652109 295354 652175 295357
rect 649950 295352 652175 295354
rect 649950 295296 652114 295352
rect 652170 295296 652175 295352
rect 649950 295294 652175 295296
rect 41781 295291 41847 295294
rect 43161 295291 43227 295294
rect 652109 295291 652175 295294
rect 675334 295292 675340 295356
rect 675404 295354 675410 295356
rect 675569 295354 675635 295357
rect 675404 295352 675635 295354
rect 675404 295296 675574 295352
rect 675630 295296 675635 295352
rect 675404 295294 675635 295296
rect 675404 295292 675410 295294
rect 675569 295291 675635 295294
rect 35801 295218 35867 295221
rect 35788 295216 35867 295218
rect 35788 295160 35806 295216
rect 35862 295160 35867 295216
rect 35788 295158 35867 295160
rect 35801 295155 35867 295158
rect 33777 294810 33843 294813
rect 33764 294808 33843 294810
rect 33764 294752 33782 294808
rect 33838 294752 33843 294808
rect 33764 294750 33843 294752
rect 33777 294747 33843 294750
rect 675753 294538 675819 294541
rect 676622 294538 676628 294540
rect 675753 294536 676628 294538
rect 32397 294402 32463 294405
rect 32397 294400 32476 294402
rect 32397 294344 32402 294400
rect 32458 294344 32476 294400
rect 32397 294342 32476 294344
rect 32397 294339 32463 294342
rect 62113 294130 62179 294133
rect 64646 294130 64706 294502
rect 649950 294266 650010 294502
rect 675753 294480 675758 294536
rect 675814 294480 676628 294536
rect 675753 294478 676628 294480
rect 675753 294475 675819 294478
rect 676622 294476 676628 294478
rect 676692 294476 676698 294540
rect 651465 294266 651531 294269
rect 649950 294264 651531 294266
rect 649950 294208 651470 294264
rect 651526 294208 651531 294264
rect 649950 294206 651531 294208
rect 651465 294203 651531 294206
rect 62113 294128 64706 294130
rect 62113 294072 62118 294128
rect 62174 294072 64706 294128
rect 62113 294070 64706 294072
rect 62113 294067 62179 294070
rect 44725 293994 44791 293997
rect 41492 293992 44791 293994
rect 41492 293936 44730 293992
rect 44786 293936 44791 293992
rect 41492 293934 44791 293936
rect 44725 293931 44791 293934
rect 662413 293858 662479 293861
rect 675201 293858 675267 293861
rect 662413 293856 675267 293858
rect 662413 293800 662418 293856
rect 662474 293800 675206 293856
rect 675262 293800 675267 293856
rect 662413 293798 675267 293800
rect 662413 293795 662479 293798
rect 675201 293795 675267 293798
rect 44541 293586 44607 293589
rect 41492 293584 44607 293586
rect 41492 293528 44546 293584
rect 44602 293528 44607 293584
rect 41492 293526 44607 293528
rect 44541 293523 44607 293526
rect 35801 293178 35867 293181
rect 35788 293176 35867 293178
rect 35788 293120 35806 293176
rect 35862 293120 35867 293176
rect 35788 293118 35867 293120
rect 35801 293115 35867 293118
rect 35801 292770 35867 292773
rect 35788 292768 35867 292770
rect 35788 292712 35806 292768
rect 35862 292712 35867 292768
rect 35788 292710 35867 292712
rect 35801 292707 35867 292710
rect 62297 292770 62363 292773
rect 64646 292770 64706 293320
rect 649950 293042 650010 293320
rect 651465 293042 651531 293045
rect 649950 293040 651531 293042
rect 649950 292984 651470 293040
rect 651526 292984 651531 293040
rect 649950 292982 651531 292984
rect 651465 292979 651531 292982
rect 62297 292768 64706 292770
rect 62297 292712 62302 292768
rect 62358 292712 64706 292768
rect 62297 292710 64706 292712
rect 62297 292707 62363 292710
rect 41362 292528 41368 292592
rect 41432 292528 41438 292592
rect 41370 292362 41430 292528
rect 62113 292498 62179 292501
rect 62113 292496 64706 292498
rect 62113 292440 62118 292496
rect 62174 292440 64706 292496
rect 62113 292438 64706 292440
rect 62113 292435 62179 292438
rect 41370 292302 41492 292362
rect 41781 292226 41847 292229
rect 43621 292226 43687 292229
rect 41781 292224 43687 292226
rect 41781 292168 41786 292224
rect 41842 292168 43626 292224
rect 43682 292168 43687 292224
rect 41781 292166 43687 292168
rect 41781 292163 41847 292166
rect 43621 292163 43687 292166
rect 64646 292138 64706 292438
rect 675569 292228 675635 292229
rect 675518 292164 675524 292228
rect 675588 292226 675635 292228
rect 675588 292224 675680 292226
rect 675630 292168 675680 292224
rect 675588 292166 675680 292168
rect 675588 292164 675635 292166
rect 675569 292163 675635 292164
rect 41781 291954 41847 291957
rect 41492 291952 41847 291954
rect 41492 291896 41786 291952
rect 41842 291896 41847 291952
rect 41492 291894 41847 291896
rect 41781 291891 41847 291894
rect 41822 291546 41828 291548
rect 41492 291486 41828 291546
rect 41822 291484 41828 291486
rect 41892 291484 41898 291548
rect 649950 291546 650010 292138
rect 652385 291546 652451 291549
rect 649950 291544 652451 291546
rect 649950 291488 652390 291544
rect 652446 291488 652451 291544
rect 649950 291486 652451 291488
rect 652385 291483 652451 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 35801 291138 35867 291141
rect 35788 291136 35867 291138
rect 35788 291080 35806 291136
rect 35862 291080 35867 291136
rect 35788 291078 35867 291080
rect 35801 291075 35867 291078
rect 62113 291002 62179 291005
rect 62113 291000 64154 291002
rect 62113 290944 62118 291000
rect 62174 290986 64154 291000
rect 62174 290944 64676 290986
rect 62113 290942 64676 290944
rect 62113 290939 62179 290942
rect 64094 290926 64676 290942
rect 50521 290730 50587 290733
rect 41492 290728 50587 290730
rect 41492 290672 50526 290728
rect 50582 290672 50587 290728
rect 41492 290670 50587 290672
rect 50521 290667 50587 290670
rect 649950 290458 650010 290956
rect 675753 290866 675819 290869
rect 676254 290866 676260 290868
rect 675753 290864 676260 290866
rect 675753 290808 675758 290864
rect 675814 290808 676260 290864
rect 675753 290806 676260 290808
rect 675753 290803 675819 290806
rect 676254 290804 676260 290806
rect 676324 290804 676330 290868
rect 651465 290458 651531 290461
rect 649950 290456 651531 290458
rect 649950 290400 651470 290456
rect 651526 290400 651531 290456
rect 649950 290398 651531 290400
rect 651465 290395 651531 290398
rect 35617 290322 35683 290325
rect 35604 290320 35683 290322
rect 35604 290264 35622 290320
rect 35678 290264 35683 290320
rect 35604 290262 35683 290264
rect 35617 290259 35683 290262
rect 41781 290322 41847 290325
rect 43345 290322 43411 290325
rect 41781 290320 43411 290322
rect 41781 290264 41786 290320
rect 41842 290264 43350 290320
rect 43406 290264 43411 290320
rect 41781 290262 43411 290264
rect 41781 290259 41847 290262
rect 43345 290259 43411 290262
rect 48957 289914 49023 289917
rect 41492 289912 49023 289914
rect 41492 289856 48962 289912
rect 49018 289856 49023 289912
rect 41492 289854 49023 289856
rect 48957 289851 49023 289854
rect 62757 289778 62823 289781
rect 62757 289776 64706 289778
rect 62757 289720 62762 289776
rect 62818 289720 64706 289776
rect 62757 289718 64706 289720
rect 62757 289715 62823 289718
rect 40718 289172 40724 289236
rect 40788 289234 40794 289236
rect 41781 289234 41847 289237
rect 40788 289232 41847 289234
rect 40788 289176 41786 289232
rect 41842 289176 41847 289232
rect 40788 289174 41847 289176
rect 649950 289234 650010 289774
rect 651465 289234 651531 289237
rect 649950 289232 651531 289234
rect 649950 289176 651470 289232
rect 651526 289176 651531 289232
rect 649950 289174 651531 289176
rect 40788 289172 40794 289174
rect 41781 289171 41847 289174
rect 651465 289171 651531 289174
rect 62113 288554 62179 288557
rect 64646 288554 64706 288592
rect 62113 288552 64706 288554
rect 62113 288496 62118 288552
rect 62174 288496 64706 288552
rect 62113 288494 64706 288496
rect 649950 288554 650010 288592
rect 651741 288554 651807 288557
rect 649950 288552 651807 288554
rect 649950 288496 651746 288552
rect 651802 288496 651807 288552
rect 649950 288494 651807 288496
rect 62113 288491 62179 288494
rect 651741 288491 651807 288494
rect 672533 287874 672599 287877
rect 675109 287874 675175 287877
rect 672533 287872 675175 287874
rect 672533 287816 672538 287872
rect 672594 287816 675114 287872
rect 675170 287816 675175 287872
rect 672533 287814 675175 287816
rect 672533 287811 672599 287814
rect 675109 287811 675175 287814
rect 651465 287466 651531 287469
rect 649766 287464 651531 287466
rect 63125 287194 63191 287197
rect 64646 287194 64706 287410
rect 649766 287408 651470 287464
rect 651526 287408 651531 287464
rect 649766 287406 651531 287408
rect 651465 287403 651531 287406
rect 63125 287192 64706 287194
rect 63125 287136 63130 287192
rect 63186 287136 64706 287192
rect 63125 287134 64706 287136
rect 63125 287131 63191 287134
rect 674005 286514 674071 286517
rect 675385 286514 675451 286517
rect 674005 286512 675451 286514
rect 674005 286456 674010 286512
rect 674066 286456 675390 286512
rect 675446 286456 675451 286512
rect 674005 286454 675451 286456
rect 674005 286451 674071 286454
rect 675385 286451 675451 286454
rect 62113 285970 62179 285973
rect 64646 285970 64706 286228
rect 62113 285968 64706 285970
rect 62113 285912 62118 285968
rect 62174 285912 64706 285968
rect 62113 285910 64706 285912
rect 649950 285970 650010 286228
rect 651465 285970 651531 285973
rect 649950 285968 651531 285970
rect 649950 285912 651470 285968
rect 651526 285912 651531 285968
rect 649950 285910 651531 285912
rect 62113 285907 62179 285910
rect 651465 285907 651531 285910
rect 672993 285562 673059 285565
rect 675109 285562 675175 285565
rect 672993 285560 675175 285562
rect 672993 285504 672998 285560
rect 673054 285504 675114 285560
rect 675170 285504 675175 285560
rect 672993 285502 675175 285504
rect 672993 285499 673059 285502
rect 675109 285499 675175 285502
rect 32397 284882 32463 284885
rect 41638 284882 41644 284884
rect 32397 284880 41644 284882
rect 32397 284824 32402 284880
rect 32458 284824 41644 284880
rect 32397 284822 41644 284824
rect 32397 284819 32463 284822
rect 41638 284820 41644 284822
rect 41708 284820 41714 284884
rect 62113 284474 62179 284477
rect 64646 284474 64706 285046
rect 649950 284746 650010 285046
rect 651465 284746 651531 284749
rect 649950 284744 651531 284746
rect 649950 284688 651470 284744
rect 651526 284688 651531 284744
rect 649950 284686 651531 284688
rect 651465 284683 651531 284686
rect 62113 284472 64706 284474
rect 62113 284416 62118 284472
rect 62174 284416 64706 284472
rect 62113 284414 64706 284416
rect 62113 284411 62179 284414
rect 40677 284338 40743 284341
rect 42006 284338 42012 284340
rect 40677 284336 42012 284338
rect 40677 284280 40682 284336
rect 40738 284280 42012 284336
rect 40677 284278 42012 284280
rect 40677 284275 40743 284278
rect 42006 284276 42012 284278
rect 42076 284276 42082 284340
rect 668117 283930 668183 283933
rect 672809 283930 672875 283933
rect 668117 283928 672875 283930
rect 668117 283872 668122 283928
rect 668178 283872 672814 283928
rect 672870 283872 672875 283928
rect 668117 283870 672875 283872
rect 668117 283867 668183 283870
rect 672809 283867 672875 283870
rect 62757 283250 62823 283253
rect 64646 283250 64706 283864
rect 62757 283248 64706 283250
rect 62757 283192 62762 283248
rect 62818 283192 64706 283248
rect 62757 283190 64706 283192
rect 649950 283250 650010 283864
rect 675661 283658 675727 283661
rect 675886 283658 675892 283660
rect 675661 283656 675892 283658
rect 675661 283600 675666 283656
rect 675722 283600 675892 283656
rect 675661 283598 675892 283600
rect 675661 283595 675727 283598
rect 675886 283596 675892 283598
rect 675956 283596 675962 283660
rect 652109 283522 652175 283525
rect 674373 283522 674439 283525
rect 652109 283520 674439 283522
rect 652109 283464 652114 283520
rect 652170 283464 674378 283520
rect 674434 283464 674439 283520
rect 652109 283462 674439 283464
rect 652109 283459 652175 283462
rect 674373 283459 674439 283462
rect 652569 283250 652635 283253
rect 649950 283248 652635 283250
rect 649950 283192 652574 283248
rect 652630 283192 652635 283248
rect 649950 283190 652635 283192
rect 62757 283187 62823 283190
rect 652569 283187 652635 283190
rect 675661 282844 675727 282845
rect 675661 282840 675708 282844
rect 675772 282842 675778 282844
rect 675661 282784 675666 282840
rect 675661 282780 675708 282784
rect 675772 282782 675818 282842
rect 675772 282780 675778 282782
rect 675661 282779 675727 282780
rect 62941 282162 63007 282165
rect 64646 282162 64706 282682
rect 62941 282160 64706 282162
rect 62941 282104 62946 282160
rect 63002 282104 64706 282160
rect 62941 282102 64706 282104
rect 649950 282162 650010 282682
rect 651925 282162 651991 282165
rect 649950 282160 651991 282162
rect 649950 282104 651930 282160
rect 651986 282104 651991 282160
rect 649950 282102 651991 282104
rect 62941 282099 63007 282102
rect 651925 282099 651991 282102
rect 62113 280938 62179 280941
rect 64646 280938 64706 281500
rect 62113 280936 64706 280938
rect 62113 280880 62118 280936
rect 62174 280880 64706 280936
rect 62113 280878 64706 280880
rect 649950 280938 650010 281500
rect 675753 281210 675819 281213
rect 676070 281210 676076 281212
rect 675753 281208 676076 281210
rect 675753 281152 675758 281208
rect 675814 281152 676076 281208
rect 675753 281150 676076 281152
rect 675753 281147 675819 281150
rect 676070 281148 676076 281150
rect 676140 281148 676146 281212
rect 651649 280938 651715 280941
rect 649950 280936 651715 280938
rect 649950 280880 651654 280936
rect 651710 280880 651715 280936
rect 649950 280878 651715 280880
rect 62113 280875 62179 280878
rect 651649 280875 651715 280878
rect 61377 280394 61443 280397
rect 651465 280394 651531 280397
rect 61377 280392 64706 280394
rect 61377 280336 61382 280392
rect 61438 280336 64706 280392
rect 61377 280334 64706 280336
rect 61377 280331 61443 280334
rect 64646 280318 64706 280334
rect 649950 280392 651531 280394
rect 649950 280336 651470 280392
rect 651526 280336 651531 280392
rect 649950 280334 651531 280336
rect 649950 280318 650010 280334
rect 651465 280331 651531 280334
rect 42425 278762 42491 278765
rect 58617 278762 58683 278765
rect 42425 278760 58683 278762
rect 42425 278704 42430 278760
rect 42486 278704 58622 278760
rect 58678 278704 58683 278760
rect 42425 278702 58683 278704
rect 42425 278699 42491 278702
rect 58617 278699 58683 278702
rect 40902 278428 40908 278492
rect 40972 278490 40978 278492
rect 41781 278490 41847 278493
rect 40972 278488 41847 278490
rect 40972 278432 41786 278488
rect 41842 278432 41847 278488
rect 40972 278430 41847 278432
rect 40972 278428 40978 278430
rect 41781 278427 41847 278430
rect 42057 277810 42123 277813
rect 43621 277810 43687 277813
rect 42057 277808 43687 277810
rect 42057 277752 42062 277808
rect 42118 277752 43626 277808
rect 43682 277752 43687 277808
rect 42057 277750 43687 277752
rect 42057 277747 42123 277750
rect 43621 277747 43687 277750
rect 40718 277068 40724 277132
rect 40788 277130 40794 277132
rect 41781 277130 41847 277133
rect 40788 277128 41847 277130
rect 40788 277072 41786 277128
rect 41842 277072 41847 277128
rect 40788 277070 41847 277072
rect 40788 277068 40794 277070
rect 41781 277067 41847 277070
rect 42057 276722 42123 276725
rect 42609 276722 42675 276725
rect 42057 276720 42675 276722
rect 42057 276664 42062 276720
rect 42118 276664 42614 276720
rect 42670 276664 42675 276720
rect 42057 276662 42675 276664
rect 42057 276659 42123 276662
rect 42609 276659 42675 276662
rect 42241 275906 42307 275909
rect 57237 275906 57303 275909
rect 42241 275904 57303 275906
rect 42241 275848 42246 275904
rect 42302 275848 57242 275904
rect 57298 275848 57303 275904
rect 42241 275846 57303 275848
rect 42241 275843 42307 275846
rect 57237 275843 57303 275846
rect 537293 275090 537359 275093
rect 538121 275090 538187 275093
rect 537293 275088 538187 275090
rect 537293 275032 537298 275088
rect 537354 275032 538126 275088
rect 538182 275032 538187 275088
rect 537293 275030 538187 275032
rect 537293 275027 537359 275030
rect 538121 275027 538187 275030
rect 542261 274818 542327 274821
rect 543181 274818 543247 274821
rect 542261 274816 543247 274818
rect 542261 274760 542266 274816
rect 542322 274760 543186 274816
rect 543242 274760 543247 274816
rect 542261 274758 543247 274760
rect 542261 274755 542327 274758
rect 543181 274755 543247 274758
rect 539317 274546 539383 274549
rect 543825 274546 543891 274549
rect 539317 274544 543891 274546
rect 539317 274488 539322 274544
rect 539378 274488 543830 274544
rect 543886 274488 543891 274544
rect 539317 274486 543891 274488
rect 539317 274483 539383 274486
rect 543825 274483 543891 274486
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 544009 273322 544075 273325
rect 552565 273322 552631 273325
rect 544009 273320 552631 273322
rect 544009 273264 544014 273320
rect 544070 273264 552570 273320
rect 552626 273264 552631 273320
rect 544009 273262 552631 273264
rect 544009 273259 544075 273262
rect 552565 273259 552631 273262
rect 42333 273186 42399 273189
rect 44541 273186 44607 273189
rect 42333 273184 44607 273186
rect 42333 273128 42338 273184
rect 42394 273128 44546 273184
rect 44602 273128 44607 273184
rect 42333 273126 44607 273128
rect 42333 273123 42399 273126
rect 44541 273123 44607 273126
rect 42425 272914 42491 272917
rect 44725 272914 44791 272917
rect 42425 272912 44791 272914
rect 42425 272856 42430 272912
rect 42486 272856 44730 272912
rect 44786 272856 44791 272912
rect 42425 272854 44791 272856
rect 42425 272851 42491 272854
rect 44725 272851 44791 272854
rect 489913 272778 489979 272781
rect 495709 272778 495775 272781
rect 489913 272776 495775 272778
rect 489913 272720 489918 272776
rect 489974 272720 495714 272776
rect 495770 272720 495775 272776
rect 489913 272718 495775 272720
rect 489913 272715 489979 272718
rect 495709 272715 495775 272718
rect 470409 272642 470475 272645
rect 470593 272642 470659 272645
rect 470409 272640 470659 272642
rect 470409 272584 470414 272640
rect 470470 272584 470598 272640
rect 470654 272584 470659 272640
rect 470409 272582 470659 272584
rect 470409 272579 470475 272582
rect 470593 272579 470659 272582
rect 41965 272372 42031 272373
rect 41965 272368 42012 272372
rect 42076 272370 42082 272372
rect 462221 272370 462287 272373
rect 470409 272370 470475 272373
rect 41965 272312 41970 272368
rect 41965 272308 42012 272312
rect 42076 272310 42122 272370
rect 462221 272368 470475 272370
rect 462221 272312 462226 272368
rect 462282 272312 470414 272368
rect 470470 272312 470475 272368
rect 462221 272310 470475 272312
rect 42076 272308 42082 272310
rect 41965 272307 42031 272308
rect 462221 272307 462287 272310
rect 470409 272307 470475 272310
rect 470593 271962 470659 271965
rect 478045 271962 478111 271965
rect 470593 271960 478111 271962
rect 470593 271904 470598 271960
rect 470654 271904 478050 271960
rect 478106 271904 478111 271960
rect 470593 271902 478111 271904
rect 470593 271899 470659 271902
rect 478045 271899 478111 271902
rect 523861 271146 523927 271149
rect 525333 271146 525399 271149
rect 523861 271144 525399 271146
rect 523861 271088 523866 271144
rect 523922 271088 525338 271144
rect 525394 271088 525399 271144
rect 523861 271086 525399 271088
rect 523861 271083 523927 271086
rect 525333 271083 525399 271086
rect 656157 271146 656223 271149
rect 683113 271146 683179 271149
rect 656157 271144 683179 271146
rect 656157 271088 656162 271144
rect 656218 271088 683118 271144
rect 683174 271088 683179 271144
rect 656157 271086 683179 271088
rect 656157 271083 656223 271086
rect 683113 271083 683179 271086
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 530393 270194 530459 270197
rect 534073 270194 534139 270197
rect 530393 270192 534139 270194
rect 530393 270136 530398 270192
rect 530454 270136 534078 270192
rect 534134 270136 534139 270192
rect 530393 270134 534139 270136
rect 530393 270131 530459 270134
rect 534073 270131 534139 270134
rect 41873 270060 41939 270061
rect 41822 270058 41828 270060
rect 41782 269998 41828 270058
rect 41892 270056 41939 270060
rect 41934 270000 41939 270056
rect 41822 269996 41828 269998
rect 41892 269996 41939 270000
rect 41873 269995 41939 269996
rect 537753 269922 537819 269925
rect 538305 269922 538371 269925
rect 537753 269920 538371 269922
rect 537753 269864 537758 269920
rect 537814 269864 538310 269920
rect 538366 269864 538371 269920
rect 537753 269862 538371 269864
rect 537753 269859 537819 269862
rect 538305 269859 538371 269862
rect 665817 268562 665883 268565
rect 676262 268562 676322 268668
rect 683113 268562 683179 268565
rect 665817 268560 676322 268562
rect 665817 268504 665822 268560
rect 665878 268504 676322 268560
rect 665817 268502 676322 268504
rect 683070 268560 683179 268562
rect 683070 268504 683118 268560
rect 683174 268504 683179 268560
rect 665817 268499 665883 268502
rect 683070 268499 683179 268504
rect 683070 268260 683130 268499
rect 674373 267882 674439 267885
rect 674373 267880 676292 267882
rect 674373 267824 674378 267880
rect 674434 267824 676292 267880
rect 674373 267822 676292 267824
rect 674373 267819 674439 267822
rect 673361 267474 673427 267477
rect 673361 267472 676292 267474
rect 673361 267416 673366 267472
rect 673422 267416 676292 267472
rect 673361 267414 676292 267416
rect 673361 267411 673427 267414
rect 40677 267066 40743 267069
rect 63125 267066 63191 267069
rect 40677 267064 63191 267066
rect 40677 267008 40682 267064
rect 40738 267008 63130 267064
rect 63186 267008 63191 267064
rect 40677 267006 63191 267008
rect 40677 267003 40743 267006
rect 63125 267003 63191 267006
rect 673913 267066 673979 267069
rect 673913 267064 676292 267066
rect 673913 267008 673918 267064
rect 673974 267008 676292 267064
rect 673913 267006 676292 267008
rect 673913 267003 673979 267006
rect 673177 266658 673243 266661
rect 673177 266656 676292 266658
rect 673177 266600 673182 266656
rect 673238 266600 676292 266656
rect 673177 266598 676292 266600
rect 673177 266595 673243 266598
rect 42149 266250 42215 266253
rect 54477 266250 54543 266253
rect 42149 266248 54543 266250
rect 42149 266192 42154 266248
rect 42210 266192 54482 266248
rect 54538 266192 54543 266248
rect 42149 266190 54543 266192
rect 42149 266187 42215 266190
rect 54477 266187 54543 266190
rect 674373 266250 674439 266253
rect 674373 266248 676292 266250
rect 674373 266192 674378 266248
rect 674434 266192 676292 266248
rect 674373 266190 676292 266192
rect 674373 266187 674439 266190
rect 674189 265842 674255 265845
rect 674189 265840 676292 265842
rect 674189 265784 674194 265840
rect 674250 265784 676292 265840
rect 674189 265782 676292 265784
rect 674189 265779 674255 265782
rect 674097 265434 674163 265437
rect 674097 265432 676292 265434
rect 674097 265376 674102 265432
rect 674158 265376 676292 265432
rect 674097 265374 676292 265376
rect 674097 265371 674163 265374
rect 674557 265026 674623 265029
rect 674557 265024 676292 265026
rect 674557 264968 674562 265024
rect 674618 264968 676292 265024
rect 674557 264966 676292 264968
rect 674557 264963 674623 264966
rect 674649 264618 674715 264621
rect 674649 264616 676292 264618
rect 674649 264560 674654 264616
rect 674710 264560 676292 264616
rect 674649 264558 676292 264560
rect 674649 264555 674715 264558
rect 674966 264148 674972 264212
rect 675036 264210 675042 264212
rect 675036 264150 676292 264210
rect 675036 264148 675042 264150
rect 676070 263604 676076 263668
rect 676140 263666 676146 263668
rect 676262 263666 676322 263772
rect 676140 263606 676322 263666
rect 676140 263604 676146 263606
rect 681046 263261 681106 263364
rect 680997 263256 681106 263261
rect 680997 263200 681002 263256
rect 681058 263200 681106 263256
rect 680997 263198 681106 263200
rect 680997 263195 681063 263198
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 674281 262578 674347 262581
rect 674281 262576 676292 262578
rect 674281 262520 674286 262576
rect 674342 262520 676292 262576
rect 674281 262518 676292 262520
rect 674281 262515 674347 262518
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671889 262170 671955 262173
rect 671889 262168 676292 262170
rect 671889 262112 671894 262168
rect 671950 262112 676292 262168
rect 671889 262110 676292 262112
rect 671889 262107 671955 262110
rect 676814 261628 676874 261732
rect 676806 261564 676812 261628
rect 676876 261564 676882 261628
rect 670417 261354 670483 261357
rect 670417 261352 676292 261354
rect 670417 261296 670422 261352
rect 670478 261296 676292 261352
rect 670417 261294 676292 261296
rect 670417 261291 670483 261294
rect 671705 260946 671771 260949
rect 671705 260944 676292 260946
rect 671705 260888 671710 260944
rect 671766 260888 676292 260944
rect 671705 260886 676292 260888
rect 671705 260883 671771 260886
rect 673361 260538 673427 260541
rect 673361 260536 676292 260538
rect 673361 260480 673366 260536
rect 673422 260480 676292 260536
rect 673361 260478 676292 260480
rect 673361 260475 673427 260478
rect 554313 259994 554379 259997
rect 676998 259996 677058 260100
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 676990 259932 676996 259996
rect 677060 259932 677066 259996
rect 670233 259722 670299 259725
rect 670233 259720 676292 259722
rect 670233 259664 670238 259720
rect 670294 259664 676292 259720
rect 670233 259662 676292 259664
rect 670233 259659 670299 259662
rect 674741 259314 674807 259317
rect 674741 259312 676292 259314
rect 674741 259256 674746 259312
rect 674802 259256 676292 259312
rect 674741 259254 676292 259256
rect 674741 259251 674807 259254
rect 673177 258906 673243 258909
rect 673177 258904 676292 258906
rect 673177 258848 673182 258904
rect 673238 258848 676292 258904
rect 673177 258846 676292 258848
rect 673177 258843 673243 258846
rect 671337 258498 671403 258501
rect 671337 258496 676292 258498
rect 671337 258440 671342 258496
rect 671398 258440 676292 258496
rect 671337 258438 676292 258440
rect 671337 258435 671403 258438
rect 46197 258090 46263 258093
rect 41492 258088 46263 258090
rect 41492 258032 46202 258088
rect 46258 258032 46263 258088
rect 41492 258030 46263 258032
rect 46197 258027 46263 258030
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 41462 257546 41522 257652
rect 683070 257549 683130 258060
rect 41462 257486 51090 257546
rect 35758 257141 35818 257244
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 44173 256866 44239 256869
rect 41492 256864 44239 256866
rect 41492 256808 44178 256864
rect 44234 256808 44239 256864
rect 41492 256806 44239 256808
rect 44173 256803 44239 256806
rect 51030 256730 51090 257486
rect 683021 257544 683130 257549
rect 683021 257488 683026 257544
rect 683082 257488 683130 257544
rect 683021 257486 683130 257488
rect 683021 257483 683087 257486
rect 676262 257141 676322 257244
rect 676213 257136 676322 257141
rect 676213 257080 676218 257136
rect 676274 257080 676322 257136
rect 676213 257078 676322 257080
rect 676213 257075 676279 257078
rect 59997 256730 60063 256733
rect 51030 256728 60063 256730
rect 51030 256672 60002 256728
rect 60058 256672 60063 256728
rect 51030 256670 60063 256672
rect 59997 256667 60063 256670
rect 650637 256730 650703 256733
rect 676262 256730 676322 256836
rect 650637 256728 676322 256730
rect 650637 256672 650642 256728
rect 650698 256672 676322 256728
rect 650637 256670 676322 256672
rect 650637 256667 650703 256670
rect 44817 256458 44883 256461
rect 41492 256456 44883 256458
rect 41492 256400 44822 256456
rect 44878 256400 44883 256456
rect 41492 256398 44883 256400
rect 44817 256395 44883 256398
rect 670785 256458 670851 256461
rect 676213 256458 676279 256461
rect 670785 256456 676279 256458
rect 670785 256400 670790 256456
rect 670846 256400 676218 256456
rect 676274 256400 676279 256456
rect 670785 256398 676279 256400
rect 670785 256395 670851 256398
rect 676213 256395 676279 256398
rect 35758 255917 35818 256020
rect 35758 255912 35867 255917
rect 35758 255856 35806 255912
rect 35862 255856 35867 255912
rect 35758 255854 35867 255856
rect 35801 255851 35867 255854
rect 39757 255914 39823 255917
rect 42793 255914 42859 255917
rect 39757 255912 42859 255914
rect 39757 255856 39762 255912
rect 39818 255856 42798 255912
rect 42854 255856 42859 255912
rect 39757 255854 42859 255856
rect 39757 255851 39823 255854
rect 42793 255851 42859 255854
rect 45553 255642 45619 255645
rect 553485 255642 553551 255645
rect 41492 255640 45619 255642
rect 41492 255584 45558 255640
rect 45614 255584 45619 255640
rect 41492 255582 45619 255584
rect 552460 255640 553551 255642
rect 552460 255584 553490 255640
rect 553546 255584 553551 255640
rect 552460 255582 553551 255584
rect 45553 255579 45619 255582
rect 553485 255579 553551 255582
rect 45001 255234 45067 255237
rect 41492 255232 45067 255234
rect 41492 255176 45006 255232
rect 45062 255176 45067 255232
rect 41492 255174 45067 255176
rect 45001 255171 45067 255174
rect 675293 254962 675359 254965
rect 680997 254962 681063 254965
rect 675293 254960 681063 254962
rect 675293 254904 675298 254960
rect 675354 254904 681002 254960
rect 681058 254904 681063 254960
rect 675293 254902 681063 254904
rect 675293 254899 675359 254902
rect 680997 254899 681063 254902
rect 44633 254826 44699 254829
rect 41492 254824 44699 254826
rect 41492 254768 44638 254824
rect 44694 254768 44699 254824
rect 41492 254766 44699 254768
rect 44633 254763 44699 254766
rect 675017 254690 675083 254693
rect 676029 254690 676095 254693
rect 675017 254688 676095 254690
rect 675017 254632 675022 254688
rect 675078 254632 676034 254688
rect 676090 254632 676095 254688
rect 675017 254630 676095 254632
rect 675017 254627 675083 254630
rect 676029 254627 676095 254630
rect 44357 254418 44423 254421
rect 41492 254416 44423 254418
rect 41492 254360 44362 254416
rect 44418 254360 44423 254416
rect 41492 254358 44423 254360
rect 44357 254355 44423 254358
rect 35758 253877 35818 253980
rect 35758 253872 35867 253877
rect 35758 253816 35806 253872
rect 35862 253816 35867 253872
rect 35758 253814 35867 253816
rect 35801 253811 35867 253814
rect 39573 253874 39639 253877
rect 42793 253874 42859 253877
rect 39573 253872 42859 253874
rect 39573 253816 39578 253872
rect 39634 253816 42798 253872
rect 42854 253816 42859 253872
rect 39573 253814 42859 253816
rect 39573 253811 39639 253814
rect 42793 253811 42859 253814
rect 35574 253469 35634 253572
rect 35574 253464 35683 253469
rect 554405 253466 554471 253469
rect 35574 253408 35622 253464
rect 35678 253408 35683 253464
rect 35574 253406 35683 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 35617 253403 35683 253406
rect 554405 253403 554471 253406
rect 35758 253061 35818 253164
rect 35758 253056 35867 253061
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252998 35867 253000
rect 35801 252995 35867 252998
rect 40953 253058 41019 253061
rect 43253 253058 43319 253061
rect 40953 253056 43319 253058
rect 40953 253000 40958 253056
rect 41014 253000 43258 253056
rect 43314 253000 43319 253056
rect 40953 252998 43319 253000
rect 40953 252995 41019 252998
rect 43253 252995 43319 252998
rect 44357 252786 44423 252789
rect 41492 252784 44423 252786
rect 41492 252728 44362 252784
rect 44418 252728 44423 252784
rect 41492 252726 44423 252728
rect 44357 252723 44423 252726
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 40493 252242 40559 252245
rect 42425 252242 42491 252245
rect 40493 252240 42491 252242
rect 40493 252184 40498 252240
rect 40554 252184 42430 252240
rect 42486 252184 42491 252240
rect 40493 252182 42491 252184
rect 40493 252179 40559 252182
rect 42425 252179 42491 252182
rect 45001 251970 45067 251973
rect 41492 251968 45067 251970
rect 41492 251912 45006 251968
rect 45062 251912 45067 251968
rect 41492 251910 45067 251912
rect 45001 251907 45067 251910
rect 44173 251562 44239 251565
rect 41492 251560 44239 251562
rect 41492 251504 44178 251560
rect 44234 251504 44239 251560
rect 41492 251502 44239 251504
rect 44173 251499 44239 251502
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 45921 251154 45987 251157
rect 41492 251152 45987 251154
rect 41492 251096 45926 251152
rect 45982 251096 45987 251152
rect 41492 251094 45987 251096
rect 45921 251091 45987 251094
rect 670969 250882 671035 250885
rect 675477 250882 675543 250885
rect 670969 250880 675543 250882
rect 670969 250824 670974 250880
rect 671030 250824 675482 250880
rect 675538 250824 675543 250880
rect 670969 250822 675543 250824
rect 670969 250819 671035 250822
rect 675477 250819 675543 250822
rect 35758 250613 35818 250716
rect 35758 250608 35867 250613
rect 35758 250552 35806 250608
rect 35862 250552 35867 250608
rect 35758 250550 35867 250552
rect 35801 250547 35867 250550
rect 40542 250204 40602 250308
rect 40534 250140 40540 250204
rect 40604 250140 40610 250204
rect 675753 250202 675819 250205
rect 676806 250202 676812 250204
rect 675753 250200 676812 250202
rect 675753 250144 675758 250200
rect 675814 250144 676812 250200
rect 675753 250142 676812 250144
rect 675753 250139 675819 250142
rect 676806 250140 676812 250142
rect 676876 250140 676882 250204
rect 40726 249796 40786 249900
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 674966 249732 674972 249796
rect 675036 249732 675042 249796
rect 674974 249522 675034 249732
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 675385 249522 675451 249525
rect 674974 249520 675451 249522
rect 35758 249389 35818 249492
rect 674974 249464 675390 249520
rect 675446 249464 675451 249520
rect 674974 249462 675451 249464
rect 675385 249459 675451 249462
rect 35758 249384 35867 249389
rect 35758 249328 35806 249384
rect 35862 249328 35867 249384
rect 35758 249326 35867 249328
rect 35801 249323 35867 249326
rect 39389 249386 39455 249389
rect 43161 249386 43227 249389
rect 39389 249384 43227 249386
rect 39389 249328 39394 249384
rect 39450 249328 43166 249384
rect 43222 249328 43227 249384
rect 39389 249326 43227 249328
rect 39389 249323 39455 249326
rect 43161 249323 43227 249326
rect 675017 249250 675083 249253
rect 676078 249250 676138 249596
rect 675017 249248 676138 249250
rect 675017 249192 675022 249248
rect 675078 249192 676138 249248
rect 675017 249190 676138 249192
rect 675017 249187 675083 249190
rect 45185 249114 45251 249117
rect 554037 249114 554103 249117
rect 41492 249112 45251 249114
rect 41492 249056 45190 249112
rect 45246 249056 45251 249112
rect 41492 249054 45251 249056
rect 552460 249112 554103 249114
rect 552460 249056 554042 249112
rect 554098 249056 554103 249112
rect 552460 249054 554103 249056
rect 45185 249051 45251 249054
rect 554037 249051 554103 249054
rect 45737 248706 45803 248709
rect 41492 248704 45803 248706
rect 41492 248648 45742 248704
rect 45798 248648 45803 248704
rect 41492 248646 45803 248648
rect 45737 248643 45803 248646
rect 46105 248298 46171 248301
rect 41492 248296 46171 248298
rect 41492 248240 46110 248296
rect 46166 248240 46171 248296
rect 41492 248238 46171 248240
rect 46105 248235 46171 248238
rect 664437 248026 664503 248029
rect 670969 248026 671035 248029
rect 664437 248024 671035 248026
rect 664437 247968 664442 248024
rect 664498 247968 670974 248024
rect 671030 247968 671035 248024
rect 664437 247966 671035 247968
rect 664437 247963 664503 247966
rect 670969 247963 671035 247966
rect 35574 247757 35634 247860
rect 35574 247752 35683 247757
rect 35574 247696 35622 247752
rect 35678 247696 35683 247752
rect 35574 247694 35683 247696
rect 35617 247691 35683 247694
rect 49141 247482 49207 247485
rect 41492 247480 49207 247482
rect 41492 247424 49146 247480
rect 49202 247424 49207 247480
rect 41492 247422 49207 247424
rect 49141 247419 49207 247422
rect 670417 247210 670483 247213
rect 675293 247210 675359 247213
rect 670417 247208 675359 247210
rect 670417 247152 670422 247208
rect 670478 247152 675298 247208
rect 675354 247152 675359 247208
rect 670417 247150 675359 247152
rect 670417 247147 670483 247150
rect 675293 247147 675359 247150
rect 35758 246941 35818 247044
rect 35758 246936 35867 246941
rect 35758 246880 35806 246936
rect 35862 246880 35867 246936
rect 35758 246878 35867 246880
rect 35801 246875 35867 246878
rect 41505 246938 41571 246941
rect 43621 246938 43687 246941
rect 553853 246938 553919 246941
rect 41505 246936 43687 246938
rect 41505 246880 41510 246936
rect 41566 246880 43626 246936
rect 43682 246880 43687 246936
rect 41505 246878 43687 246880
rect 552460 246936 553919 246938
rect 552460 246880 553858 246936
rect 553914 246880 553919 246936
rect 552460 246878 553919 246880
rect 41505 246875 41571 246878
rect 43621 246875 43687 246878
rect 553853 246875 553919 246878
rect 671705 246938 671771 246941
rect 675201 246938 675267 246941
rect 671705 246936 675267 246938
rect 671705 246880 671710 246936
rect 671766 246880 675206 246936
rect 675262 246880 675267 246936
rect 671705 246878 675267 246880
rect 671705 246875 671771 246878
rect 675201 246875 675267 246878
rect 47577 246666 47643 246669
rect 41492 246664 47643 246666
rect 41492 246608 47582 246664
rect 47638 246608 47643 246664
rect 41492 246606 47643 246608
rect 47577 246603 47643 246606
rect 672073 246258 672139 246261
rect 673310 246258 673316 246260
rect 672073 246256 673316 246258
rect 672073 246200 672078 246256
rect 672134 246200 673316 246256
rect 672073 246198 673316 246200
rect 672073 246195 672139 246198
rect 673310 246196 673316 246198
rect 673380 246196 673386 246260
rect 670233 245578 670299 245581
rect 675201 245578 675267 245581
rect 670233 245576 675267 245578
rect 670233 245520 670238 245576
rect 670294 245520 675206 245576
rect 675262 245520 675267 245576
rect 670233 245518 675267 245520
rect 670233 245515 670299 245518
rect 675201 245515 675267 245518
rect 39205 245034 39271 245037
rect 42977 245034 43043 245037
rect 39205 245032 43043 245034
rect 39205 244976 39210 245032
rect 39266 244976 42982 245032
rect 43038 244976 43043 245032
rect 39205 244974 43043 244976
rect 39205 244971 39271 244974
rect 42977 244971 43043 244974
rect 554497 244762 554563 244765
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 554497 244699 554563 244702
rect 674281 243674 674347 243677
rect 675201 243674 675267 243677
rect 674281 243672 675267 243674
rect 674281 243616 674286 243672
rect 674342 243616 675206 243672
rect 675262 243616 675267 243672
rect 674281 243614 675267 243616
rect 674281 243611 674347 243614
rect 675201 243611 675267 243614
rect 553669 242586 553735 242589
rect 552460 242584 553735 242586
rect 552460 242528 553674 242584
rect 553730 242528 553735 242584
rect 552460 242526 553735 242528
rect 553669 242523 553735 242526
rect 675753 242314 675819 242317
rect 676990 242314 676996 242316
rect 675753 242312 676996 242314
rect 675753 242256 675758 242312
rect 675814 242256 676996 242312
rect 675753 242254 676996 242256
rect 675753 242251 675819 242254
rect 676990 242252 676996 242254
rect 677060 242252 677066 242316
rect 674097 241906 674163 241909
rect 676806 241906 676812 241908
rect 674097 241904 676812 241906
rect 674097 241848 674102 241904
rect 674158 241848 676812 241904
rect 674097 241846 676812 241848
rect 674097 241843 674163 241846
rect 676806 241844 676812 241846
rect 676876 241844 676882 241908
rect 674373 241634 674439 241637
rect 674966 241634 674972 241636
rect 674373 241632 674972 241634
rect 674373 241576 674378 241632
rect 674434 241576 674972 241632
rect 674373 241574 674972 241576
rect 674373 241571 674439 241574
rect 674966 241572 674972 241574
rect 675036 241572 675042 241636
rect 673177 241090 673243 241093
rect 675385 241090 675451 241093
rect 673177 241088 675451 241090
rect 673177 241032 673182 241088
rect 673238 241032 675390 241088
rect 675446 241032 675451 241088
rect 673177 241030 675451 241032
rect 673177 241027 673243 241030
rect 675385 241027 675451 241030
rect 554497 240410 554563 240413
rect 552460 240408 554563 240410
rect 552460 240352 554502 240408
rect 554558 240352 554563 240408
rect 552460 240350 554563 240352
rect 554497 240347 554563 240350
rect 673361 240274 673427 240277
rect 675385 240274 675451 240277
rect 673361 240272 675451 240274
rect 673361 240216 673366 240272
rect 673422 240216 675390 240272
rect 675446 240216 675451 240272
rect 673361 240214 675451 240216
rect 673361 240211 673427 240214
rect 675385 240211 675451 240214
rect 42057 240138 42123 240141
rect 44173 240138 44239 240141
rect 42057 240136 44239 240138
rect 42057 240080 42062 240136
rect 42118 240080 44178 240136
rect 44234 240080 44239 240136
rect 42057 240078 44239 240080
rect 42057 240075 42123 240078
rect 44173 240075 44239 240078
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 42006 237356 42012 237420
rect 42076 237418 42082 237420
rect 42425 237418 42491 237421
rect 42076 237416 42491 237418
rect 42076 237360 42430 237416
rect 42486 237360 42491 237416
rect 42076 237358 42491 237360
rect 42076 237356 42082 237358
rect 42425 237355 42491 237358
rect 673085 236738 673151 236741
rect 673913 236738 673979 236741
rect 673085 236736 673979 236738
rect 673085 236680 673090 236736
rect 673146 236680 673918 236736
rect 673974 236680 673979 236736
rect 673085 236678 673979 236680
rect 673085 236675 673151 236678
rect 673913 236675 673979 236678
rect 40718 236540 40724 236604
rect 40788 236602 40794 236604
rect 41781 236602 41847 236605
rect 40788 236600 41847 236602
rect 40788 236544 41786 236600
rect 41842 236544 41847 236600
rect 40788 236542 41847 236544
rect 40788 236540 40794 236542
rect 41781 236539 41847 236542
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 42425 235922 42491 235925
rect 46105 235922 46171 235925
rect 42425 235920 46171 235922
rect 42425 235864 42430 235920
rect 42486 235864 46110 235920
rect 46166 235864 46171 235920
rect 42425 235862 46171 235864
rect 42425 235859 42491 235862
rect 46105 235859 46171 235862
rect 674557 235242 674623 235245
rect 675845 235242 675911 235245
rect 674557 235240 675911 235242
rect 674557 235184 674562 235240
rect 674618 235184 675850 235240
rect 675906 235184 675911 235240
rect 674557 235182 675911 235184
rect 674557 235179 674623 235182
rect 675845 235179 675911 235182
rect 673269 234970 673335 234973
rect 672950 234968 673335 234970
rect 672950 234912 673274 234968
rect 673330 234912 673335 234968
rect 672950 234910 673335 234912
rect 672950 234698 673010 234910
rect 673269 234907 673335 234910
rect 674833 234698 674899 234701
rect 672950 234638 673194 234698
rect 669773 234290 669839 234293
rect 673134 234290 673194 234638
rect 669773 234288 673194 234290
rect 669773 234232 669778 234288
rect 669834 234232 673194 234288
rect 669773 234230 673194 234232
rect 673410 234696 674899 234698
rect 673410 234640 674838 234696
rect 674894 234640 674899 234696
rect 673410 234638 674899 234640
rect 669773 234227 669839 234230
rect 670417 234018 670483 234021
rect 673410 234018 673470 234638
rect 674833 234635 674899 234638
rect 670417 234016 673470 234018
rect 670417 233960 670422 234016
rect 670478 233960 673470 234016
rect 670417 233958 673470 233960
rect 670417 233955 670483 233958
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 674097 233882 674163 233885
rect 676029 233882 676095 233885
rect 674097 233880 676095 233882
rect 674097 233824 674102 233880
rect 674158 233824 676034 233880
rect 676090 233824 676095 233880
rect 674097 233822 676095 233824
rect 674097 233819 674163 233822
rect 676029 233819 676095 233822
rect 42425 233474 42491 233477
rect 45737 233474 45803 233477
rect 42425 233472 45803 233474
rect 42425 233416 42430 233472
rect 42486 233416 45742 233472
rect 45798 233416 45803 233472
rect 42425 233414 45803 233416
rect 42425 233411 42491 233414
rect 45737 233411 45803 233414
rect 42425 233202 42491 233205
rect 45001 233202 45067 233205
rect 42425 233200 45067 233202
rect 42425 233144 42430 233200
rect 42486 233144 45006 233200
rect 45062 233144 45067 233200
rect 42425 233142 45067 233144
rect 42425 233139 42491 233142
rect 45001 233139 45067 233142
rect 40534 233004 40540 233068
rect 40604 233066 40610 233068
rect 42241 233066 42307 233069
rect 40604 233064 42307 233066
rect 40604 233008 42246 233064
rect 42302 233008 42307 233064
rect 40604 233006 42307 233008
rect 40604 233004 40610 233006
rect 42241 233003 42307 233006
rect 671889 232522 671955 232525
rect 675845 232522 675911 232525
rect 671889 232520 675911 232522
rect 671889 232464 671894 232520
rect 671950 232464 675850 232520
rect 675906 232464 675911 232520
rect 671889 232462 675911 232464
rect 671889 232459 671955 232462
rect 675845 232459 675911 232462
rect 671889 231570 671955 231573
rect 675845 231570 675911 231573
rect 671889 231568 675911 231570
rect 671889 231512 671894 231568
rect 671950 231512 675850 231568
rect 675906 231512 675911 231568
rect 671889 231510 675911 231512
rect 671889 231507 671955 231510
rect 675845 231507 675911 231510
rect 42057 231026 42123 231029
rect 45185 231026 45251 231029
rect 42057 231024 45251 231026
rect 42057 230968 42062 231024
rect 42118 230968 45190 231024
rect 45246 230968 45251 231024
rect 42057 230966 45251 230968
rect 42057 230963 42123 230966
rect 45185 230963 45251 230966
rect 142429 230482 142495 230485
rect 144085 230482 144151 230485
rect 142429 230480 144151 230482
rect 142429 230424 142434 230480
rect 142490 230424 144090 230480
rect 144146 230424 144151 230480
rect 142429 230422 144151 230424
rect 142429 230419 142495 230422
rect 144085 230419 144151 230422
rect 665817 230482 665883 230485
rect 674669 230482 674735 230485
rect 665817 230480 674735 230482
rect 665817 230424 665822 230480
rect 665878 230424 674674 230480
rect 674730 230424 674735 230480
rect 665817 230422 674735 230424
rect 665817 230419 665883 230422
rect 674669 230419 674735 230422
rect 674833 230482 674899 230485
rect 676673 230482 676739 230485
rect 674833 230480 676739 230482
rect 674833 230424 674838 230480
rect 674894 230424 676678 230480
rect 676734 230424 676739 230480
rect 674833 230422 676739 230424
rect 674833 230419 674899 230422
rect 676673 230419 676739 230422
rect 674966 230148 674972 230212
rect 675036 230210 675042 230212
rect 676029 230210 676095 230213
rect 675036 230208 676095 230210
rect 675036 230152 676034 230208
rect 676090 230152 676095 230208
rect 675036 230150 676095 230152
rect 675036 230148 675042 230150
rect 676029 230147 676095 230150
rect 156689 229938 156755 229941
rect 157425 229938 157491 229941
rect 156689 229936 157491 229938
rect 156689 229880 156694 229936
rect 156750 229880 157430 229936
rect 157486 229880 157491 229936
rect 156689 229878 157491 229880
rect 156689 229875 156755 229878
rect 157425 229875 157491 229878
rect 147581 229802 147647 229805
rect 147949 229802 148015 229805
rect 147581 229800 148015 229802
rect 147581 229744 147586 229800
rect 147642 229744 147954 229800
rect 148010 229744 148015 229800
rect 147581 229742 148015 229744
rect 147581 229739 147647 229742
rect 147949 229739 148015 229742
rect 652569 229802 652635 229805
rect 674046 229802 674052 229804
rect 652569 229800 674052 229802
rect 652569 229744 652574 229800
rect 652630 229744 674052 229800
rect 652569 229742 674052 229744
rect 652569 229739 652635 229742
rect 674046 229740 674052 229742
rect 674116 229740 674122 229804
rect 143993 229530 144059 229533
rect 145373 229530 145439 229533
rect 143993 229528 145439 229530
rect 143993 229472 143998 229528
rect 144054 229472 145378 229528
rect 145434 229472 145439 229528
rect 143993 229470 145439 229472
rect 143993 229467 144059 229470
rect 145373 229467 145439 229470
rect 146201 229394 146267 229397
rect 147765 229394 147831 229397
rect 146201 229392 147831 229394
rect 146201 229336 146206 229392
rect 146262 229336 147770 229392
rect 147826 229336 147831 229392
rect 146201 229334 147831 229336
rect 146201 229331 146267 229334
rect 147765 229331 147831 229334
rect 150341 229394 150407 229397
rect 157057 229394 157123 229397
rect 150341 229392 157123 229394
rect 150341 229336 150346 229392
rect 150402 229336 157062 229392
rect 157118 229336 157123 229392
rect 150341 229334 157123 229336
rect 150341 229331 150407 229334
rect 157057 229331 157123 229334
rect 663701 229394 663767 229397
rect 674465 229394 674531 229397
rect 663701 229392 674531 229394
rect 663701 229336 663706 229392
rect 663762 229336 674470 229392
rect 674526 229336 674531 229392
rect 663701 229334 674531 229336
rect 663701 229331 663767 229334
rect 674465 229331 674531 229334
rect 140037 229122 140103 229125
rect 147121 229122 147187 229125
rect 140037 229120 147187 229122
rect 140037 229064 140042 229120
rect 140098 229064 147126 229120
rect 147182 229064 147187 229120
rect 140037 229062 147187 229064
rect 140037 229059 140103 229062
rect 147121 229059 147187 229062
rect 665173 229122 665239 229125
rect 673453 229122 673519 229125
rect 665173 229120 673519 229122
rect 665173 229064 665178 229120
rect 665234 229064 673458 229120
rect 673514 229064 673519 229120
rect 665173 229062 673519 229064
rect 665173 229059 665239 229062
rect 673453 229059 673519 229062
rect 41965 228988 42031 228989
rect 41965 228984 42012 228988
rect 42076 228986 42082 228988
rect 169293 228986 169359 228989
rect 172145 228986 172211 228989
rect 41965 228928 41970 228984
rect 41965 228924 42012 228928
rect 42076 228926 42122 228986
rect 169293 228984 172211 228986
rect 169293 228928 169298 228984
rect 169354 228928 172150 228984
rect 172206 228928 172211 228984
rect 169293 228926 172211 228928
rect 42076 228924 42082 228926
rect 41965 228923 42031 228924
rect 169293 228923 169359 228926
rect 172145 228923 172211 228926
rect 166809 228850 166875 228853
rect 169109 228850 169175 228853
rect 166809 228848 169175 228850
rect 166809 228792 166814 228848
rect 166870 228792 169114 228848
rect 169170 228792 169175 228848
rect 166809 228790 169175 228792
rect 166809 228787 166875 228790
rect 169109 228787 169175 228790
rect 173157 228850 173223 228853
rect 174813 228850 174879 228853
rect 173157 228848 174879 228850
rect 173157 228792 173162 228848
rect 173218 228792 174818 228848
rect 174874 228792 174879 228848
rect 173157 228790 174879 228792
rect 173157 228787 173223 228790
rect 174813 228787 174879 228790
rect 219617 228714 219683 228717
rect 220537 228714 220603 228717
rect 219617 228712 220603 228714
rect 219617 228656 219622 228712
rect 219678 228656 220542 228712
rect 220598 228656 220603 228712
rect 219617 228654 220603 228656
rect 219617 228651 219683 228654
rect 220537 228651 220603 228654
rect 674097 228578 674163 228581
rect 676397 228578 676463 228581
rect 674097 228576 676463 228578
rect 674097 228520 674102 228576
rect 674158 228520 676402 228576
rect 676458 228520 676463 228576
rect 674097 228518 676463 228520
rect 674097 228515 674163 228518
rect 676397 228515 676463 228518
rect 166809 228442 166875 228445
rect 172329 228442 172395 228445
rect 166809 228440 172395 228442
rect 166809 228384 166814 228440
rect 166870 228384 172334 228440
rect 172390 228384 172395 228440
rect 166809 228382 172395 228384
rect 166809 228379 166875 228382
rect 172329 228379 172395 228382
rect 139301 228306 139367 228309
rect 142981 228306 143047 228309
rect 139301 228304 143047 228306
rect 139301 228248 139306 228304
rect 139362 228248 142986 228304
rect 143042 228248 143047 228304
rect 139301 228246 143047 228248
rect 139301 228243 139367 228246
rect 142981 228243 143047 228246
rect 160001 228170 160067 228173
rect 166809 228170 166875 228173
rect 160001 228168 166875 228170
rect 160001 228112 160006 228168
rect 160062 228112 166814 228168
rect 166870 228112 166875 228168
rect 160001 228110 166875 228112
rect 160001 228107 160067 228110
rect 166809 228107 166875 228110
rect 171225 227626 171291 227629
rect 172145 227626 172211 227629
rect 171225 227624 172211 227626
rect 171225 227568 171230 227624
rect 171286 227568 172150 227624
rect 172206 227568 172211 227624
rect 171225 227566 172211 227568
rect 171225 227563 171291 227566
rect 172145 227563 172211 227566
rect 156689 227490 156755 227493
rect 166533 227490 166599 227493
rect 156689 227488 166599 227490
rect 156689 227432 156694 227488
rect 156750 227432 166538 227488
rect 166594 227432 166599 227488
rect 156689 227430 166599 227432
rect 156689 227427 156755 227430
rect 166533 227427 166599 227430
rect 169477 227354 169543 227357
rect 171685 227354 171751 227357
rect 169477 227352 171751 227354
rect 169477 227296 169482 227352
rect 169538 227296 171690 227352
rect 171746 227296 171751 227352
rect 169477 227294 171751 227296
rect 169477 227291 169543 227294
rect 171685 227291 171751 227294
rect 673453 227082 673519 227085
rect 677041 227082 677107 227085
rect 673453 227080 677107 227082
rect 673453 227024 673458 227080
rect 673514 227024 677046 227080
rect 677102 227024 677107 227080
rect 673453 227022 677107 227024
rect 673453 227019 673519 227022
rect 677041 227019 677107 227022
rect 673453 226810 673519 226813
rect 674097 226810 674163 226813
rect 673453 226808 674163 226810
rect 673453 226752 673458 226808
rect 673514 226752 674102 226808
rect 674158 226752 674163 226808
rect 673453 226750 674163 226752
rect 673453 226747 673519 226750
rect 674097 226747 674163 226750
rect 654777 226402 654843 226405
rect 672717 226402 672783 226405
rect 654777 226400 672783 226402
rect 654777 226344 654782 226400
rect 654838 226344 672722 226400
rect 672778 226344 672783 226400
rect 654777 226342 672783 226344
rect 654777 226339 654843 226342
rect 672717 226339 672783 226342
rect 202597 226266 202663 226269
rect 205081 226266 205147 226269
rect 202597 226264 205147 226266
rect 202597 226208 202602 226264
rect 202658 226208 205086 226264
rect 205142 226208 205147 226264
rect 202597 226206 205147 226208
rect 202597 226203 202663 226206
rect 205081 226203 205147 226206
rect 42241 226130 42307 226133
rect 44357 226130 44423 226133
rect 42241 226128 44423 226130
rect 42241 226072 42246 226128
rect 42302 226072 44362 226128
rect 44418 226072 44423 226128
rect 42241 226070 44423 226072
rect 42241 226067 42307 226070
rect 44357 226067 44423 226070
rect 141141 226130 141207 226133
rect 145189 226130 145255 226133
rect 141141 226128 145255 226130
rect 141141 226072 141146 226128
rect 141202 226072 145194 226128
rect 145250 226072 145255 226128
rect 141141 226070 145255 226072
rect 141141 226067 141207 226070
rect 145189 226067 145255 226070
rect 672257 226130 672323 226133
rect 674833 226130 674899 226133
rect 672257 226128 674899 226130
rect 672257 226072 672262 226128
rect 672318 226072 674838 226128
rect 674894 226072 674899 226128
rect 672257 226070 674899 226072
rect 672257 226067 672323 226070
rect 674833 226067 674899 226070
rect 672625 225858 672691 225861
rect 675017 225858 675083 225861
rect 672625 225856 675083 225858
rect 672625 225800 672630 225856
rect 672686 225800 675022 225856
rect 675078 225800 675083 225856
rect 672625 225798 675083 225800
rect 672625 225795 672691 225798
rect 675017 225795 675083 225798
rect 672257 225722 672323 225725
rect 663750 225720 672323 225722
rect 663750 225664 672262 225720
rect 672318 225664 672323 225720
rect 663750 225662 672323 225664
rect 42609 225586 42675 225589
rect 62941 225586 63007 225589
rect 42609 225584 63007 225586
rect 42609 225528 42614 225584
rect 42670 225528 62946 225584
rect 63002 225528 63007 225584
rect 42609 225526 63007 225528
rect 42609 225523 42675 225526
rect 62941 225523 63007 225526
rect 656157 225586 656223 225589
rect 663750 225586 663810 225662
rect 672257 225659 672323 225662
rect 656157 225584 663810 225586
rect 656157 225528 656162 225584
rect 656218 225528 663810 225584
rect 656157 225526 663810 225528
rect 656157 225523 656223 225526
rect 672073 225450 672139 225453
rect 663934 225448 672139 225450
rect 663934 225392 672078 225448
rect 672134 225392 672139 225448
rect 663934 225390 672139 225392
rect 653397 225314 653463 225317
rect 663934 225314 663994 225390
rect 672073 225387 672139 225390
rect 653397 225312 663994 225314
rect 653397 225256 653402 225312
rect 653458 225256 663994 225312
rect 653397 225254 663994 225256
rect 672257 225314 672323 225317
rect 675201 225314 675267 225317
rect 672257 225312 675267 225314
rect 672257 225256 672262 225312
rect 672318 225256 675206 225312
rect 675262 225256 675267 225312
rect 672257 225254 675267 225256
rect 653397 225251 653463 225254
rect 672257 225251 672323 225254
rect 675201 225251 675267 225254
rect 672027 225178 672093 225181
rect 664118 225176 672093 225178
rect 664118 225120 672032 225176
rect 672088 225120 672093 225176
rect 664118 225118 672093 225120
rect 657721 225042 657787 225045
rect 664118 225042 664178 225118
rect 672027 225115 672093 225118
rect 657721 225040 664178 225042
rect 657721 224984 657726 225040
rect 657782 224984 664178 225040
rect 657721 224982 664178 224984
rect 657721 224979 657787 224982
rect 42425 224906 42491 224909
rect 45921 224906 45987 224909
rect 42425 224904 45987 224906
rect 42425 224848 42430 224904
rect 42486 224848 45926 224904
rect 45982 224848 45987 224904
rect 42425 224846 45987 224848
rect 42425 224843 42491 224846
rect 45921 224843 45987 224846
rect 557073 224770 557139 224773
rect 561673 224770 561739 224773
rect 671153 224772 671219 224773
rect 671102 224770 671108 224772
rect 557073 224768 561739 224770
rect 557073 224712 557078 224768
rect 557134 224712 561678 224768
rect 561734 224712 561739 224768
rect 557073 224710 561739 224712
rect 671062 224710 671108 224770
rect 671172 224768 671219 224772
rect 671214 224712 671219 224768
rect 557073 224707 557139 224710
rect 561673 224707 561739 224710
rect 671102 224708 671108 224710
rect 671172 224708 671219 224712
rect 671153 224707 671219 224708
rect 672717 224770 672783 224773
rect 673361 224770 673427 224773
rect 672717 224768 673427 224770
rect 672717 224712 672722 224768
rect 672778 224712 673366 224768
rect 673422 224712 673427 224768
rect 672717 224710 673427 224712
rect 672717 224707 672783 224710
rect 673361 224707 673427 224710
rect 671813 224498 671879 224501
rect 663750 224496 671879 224498
rect 663750 224440 671818 224496
rect 671874 224440 671879 224496
rect 663750 224438 671879 224440
rect 657537 223954 657603 223957
rect 663750 223954 663810 224438
rect 671813 224435 671879 224438
rect 671245 224226 671311 224229
rect 673453 224226 673519 224229
rect 671245 224224 673519 224226
rect 671245 224168 671250 224224
rect 671306 224168 673458 224224
rect 673514 224168 673519 224224
rect 671245 224166 673519 224168
rect 671245 224163 671311 224166
rect 673453 224163 673519 224166
rect 657537 223952 663810 223954
rect 657537 223896 657542 223952
rect 657598 223896 663810 223952
rect 657537 223894 663810 223896
rect 657537 223891 657603 223894
rect 664437 223818 664503 223821
rect 669037 223818 669103 223821
rect 664437 223816 669103 223818
rect 664437 223760 664442 223816
rect 664498 223760 669042 223816
rect 669098 223760 669103 223816
rect 664437 223758 669103 223760
rect 664437 223755 664503 223758
rect 669037 223755 669103 223758
rect 671245 223818 671311 223821
rect 672073 223818 672139 223821
rect 671245 223816 672139 223818
rect 671245 223760 671250 223816
rect 671306 223760 672078 223816
rect 672134 223760 672139 223816
rect 671245 223758 672139 223760
rect 671245 223755 671311 223758
rect 672073 223755 672139 223758
rect 678237 223818 678303 223821
rect 678237 223816 678346 223818
rect 678237 223760 678242 223816
rect 678298 223760 678346 223816
rect 678237 223755 678346 223760
rect 678286 223516 678346 223755
rect 671015 223410 671081 223413
rect 672441 223410 672507 223413
rect 671015 223408 672507 223410
rect 671015 223352 671020 223408
rect 671076 223352 672446 223408
rect 672502 223352 672507 223408
rect 671015 223350 672507 223352
rect 671015 223347 671081 223350
rect 672441 223347 672507 223350
rect 42149 223274 42215 223277
rect 55857 223274 55923 223277
rect 42149 223272 55923 223274
rect 42149 223216 42154 223272
rect 42210 223216 55862 223272
rect 55918 223216 55923 223272
rect 42149 223214 55923 223216
rect 42149 223211 42215 223214
rect 55857 223211 55923 223214
rect 151905 223138 151971 223141
rect 156781 223138 156847 223141
rect 671153 223140 671219 223141
rect 151905 223136 156847 223138
rect 151905 223080 151910 223136
rect 151966 223080 156786 223136
rect 156842 223080 156847 223136
rect 151905 223078 156847 223080
rect 151905 223075 151971 223078
rect 156781 223075 156847 223078
rect 671102 223076 671108 223140
rect 671172 223138 671219 223140
rect 683573 223138 683639 223141
rect 671172 223136 671264 223138
rect 671214 223080 671264 223136
rect 671172 223078 671264 223080
rect 683573 223136 683652 223138
rect 683573 223080 683578 223136
rect 683634 223080 683652 223136
rect 683573 223078 683652 223080
rect 671172 223076 671219 223078
rect 671153 223075 671219 223076
rect 683573 223075 683639 223078
rect 147305 223002 147371 223005
rect 151445 223002 151511 223005
rect 147305 223000 151511 223002
rect 147305 222944 147310 223000
rect 147366 222944 151450 223000
rect 151506 222944 151511 223000
rect 147305 222942 151511 222944
rect 147305 222939 147371 222942
rect 151445 222939 151511 222942
rect 650637 222866 650703 222869
rect 672717 222866 672783 222869
rect 650637 222864 672783 222866
rect 650637 222808 650642 222864
rect 650698 222808 672722 222864
rect 672778 222808 672783 222864
rect 650637 222806 672783 222808
rect 650637 222803 650703 222806
rect 672717 222803 672783 222806
rect 151629 222730 151695 222733
rect 152089 222730 152155 222733
rect 151629 222728 152155 222730
rect 151629 222672 151634 222728
rect 151690 222672 152094 222728
rect 152150 222672 152155 222728
rect 151629 222670 152155 222672
rect 151629 222667 151695 222670
rect 152089 222667 152155 222670
rect 683205 222730 683271 222733
rect 683205 222728 683284 222730
rect 683205 222672 683210 222728
rect 683266 222672 683284 222728
rect 683205 222670 683284 222672
rect 683205 222667 683271 222670
rect 659101 222594 659167 222597
rect 669037 222594 669103 222597
rect 659101 222592 669103 222594
rect 659101 222536 659106 222592
rect 659162 222536 669042 222592
rect 669098 222536 669103 222592
rect 659101 222534 669103 222536
rect 659101 222531 659167 222534
rect 669037 222531 669103 222534
rect 145925 222322 145991 222325
rect 147121 222322 147187 222325
rect 145925 222320 147187 222322
rect 145925 222264 145930 222320
rect 145986 222264 147126 222320
rect 147182 222264 147187 222320
rect 145925 222262 147187 222264
rect 145925 222259 145991 222262
rect 147121 222259 147187 222262
rect 557901 222322 557967 222325
rect 563145 222322 563211 222325
rect 557901 222320 563211 222322
rect 557901 222264 557906 222320
rect 557962 222264 563150 222320
rect 563206 222264 563211 222320
rect 557901 222262 563211 222264
rect 557901 222259 557967 222262
rect 563145 222259 563211 222262
rect 674373 222322 674439 222325
rect 674373 222320 676292 222322
rect 674373 222264 674378 222320
rect 674434 222264 676292 222320
rect 674373 222262 676292 222264
rect 674373 222259 674439 222262
rect 552933 222186 552999 222189
rect 553577 222186 553643 222189
rect 552933 222184 553643 222186
rect 552933 222128 552938 222184
rect 552994 222128 553582 222184
rect 553638 222128 553643 222184
rect 552933 222126 553643 222128
rect 552933 222123 552999 222126
rect 553577 222123 553643 222126
rect 540881 222050 540947 222053
rect 543825 222050 543891 222053
rect 540881 222048 543891 222050
rect 540881 221992 540886 222048
rect 540942 221992 543830 222048
rect 543886 221992 543891 222048
rect 540881 221990 543891 221992
rect 540881 221987 540947 221990
rect 543825 221987 543891 221990
rect 544193 222050 544259 222053
rect 546585 222050 546651 222053
rect 544193 222048 546651 222050
rect 544193 221992 544198 222048
rect 544254 221992 546590 222048
rect 546646 221992 546651 222048
rect 544193 221990 546651 221992
rect 544193 221987 544259 221990
rect 546585 221987 546651 221990
rect 559557 222050 559623 222053
rect 562869 222050 562935 222053
rect 559557 222048 562935 222050
rect 559557 221992 559562 222048
rect 559618 221992 562874 222048
rect 562930 221992 562935 222048
rect 559557 221990 562935 221992
rect 559557 221987 559623 221990
rect 562869 221987 562935 221990
rect 547137 221914 547203 221917
rect 558545 221914 558611 221917
rect 547137 221912 558611 221914
rect 547137 221856 547142 221912
rect 547198 221856 558550 221912
rect 558606 221856 558611 221912
rect 547137 221854 558611 221856
rect 547137 221851 547203 221854
rect 558545 221851 558611 221854
rect 674230 221852 674236 221916
rect 674300 221914 674306 221916
rect 674300 221854 676292 221914
rect 674300 221852 674306 221854
rect 184657 221778 184723 221781
rect 185761 221778 185827 221781
rect 184657 221776 185827 221778
rect 184657 221720 184662 221776
rect 184718 221720 185766 221776
rect 185822 221720 185827 221776
rect 184657 221718 185827 221720
rect 184657 221715 184723 221718
rect 185761 221715 185827 221718
rect 543089 221778 543155 221781
rect 544009 221778 544075 221781
rect 543089 221776 544075 221778
rect 543089 221720 543094 221776
rect 543150 221720 544014 221776
rect 544070 221720 544075 221776
rect 543089 221718 544075 221720
rect 543089 221715 543155 221718
rect 544009 221715 544075 221718
rect 562685 221778 562751 221781
rect 568941 221778 569007 221781
rect 562685 221776 569007 221778
rect 562685 221720 562690 221776
rect 562746 221720 568946 221776
rect 569002 221720 569007 221776
rect 562685 221718 569007 221720
rect 562685 221715 562751 221718
rect 568941 221715 569007 221718
rect 651465 221778 651531 221781
rect 668025 221778 668091 221781
rect 651465 221776 668091 221778
rect 651465 221720 651470 221776
rect 651526 221720 668030 221776
rect 668086 221720 668091 221776
rect 651465 221718 668091 221720
rect 651465 221715 651531 221718
rect 668025 221715 668091 221718
rect 161933 221642 161999 221645
rect 164325 221642 164391 221645
rect 161933 221640 164391 221642
rect 161933 221584 161938 221640
rect 161994 221584 164330 221640
rect 164386 221584 164391 221640
rect 161933 221582 164391 221584
rect 161933 221579 161999 221582
rect 164325 221579 164391 221582
rect 513373 221642 513439 221645
rect 513373 221640 514770 221642
rect 513373 221584 513378 221640
rect 513434 221584 514770 221640
rect 513373 221582 514770 221584
rect 513373 221579 513439 221582
rect 514710 221506 514770 221582
rect 598933 221506 598999 221509
rect 514710 221504 598999 221506
rect 514710 221448 598938 221504
rect 598994 221448 598999 221504
rect 514710 221446 598999 221448
rect 598933 221443 598999 221446
rect 649901 221506 649967 221509
rect 674833 221506 674899 221509
rect 649901 221504 674899 221506
rect 649901 221448 649906 221504
rect 649962 221448 674838 221504
rect 674894 221448 674899 221504
rect 649901 221446 674899 221448
rect 649901 221443 649967 221446
rect 674833 221443 674899 221446
rect 676029 221506 676095 221509
rect 676029 221504 676292 221506
rect 676029 221448 676034 221504
rect 676090 221448 676292 221504
rect 676029 221446 676292 221448
rect 676029 221443 676095 221446
rect 176469 221370 176535 221373
rect 177297 221370 177363 221373
rect 176469 221368 177363 221370
rect 176469 221312 176474 221368
rect 176530 221312 177302 221368
rect 177358 221312 177363 221368
rect 176469 221310 177363 221312
rect 176469 221307 176535 221310
rect 177297 221307 177363 221310
rect 520181 221234 520247 221237
rect 618253 221234 618319 221237
rect 520181 221232 618319 221234
rect 520181 221176 520186 221232
rect 520242 221176 618258 221232
rect 618314 221176 618319 221232
rect 520181 221174 618319 221176
rect 520181 221171 520247 221174
rect 618253 221171 618319 221174
rect 667013 221098 667079 221101
rect 667013 221096 676292 221098
rect 667013 221040 667018 221096
rect 667074 221040 676292 221096
rect 667013 221038 676292 221040
rect 667013 221035 667079 221038
rect 158345 220962 158411 220965
rect 166717 220962 166783 220965
rect 158345 220960 166783 220962
rect 158345 220904 158350 220960
rect 158406 220904 166722 220960
rect 166778 220904 166783 220960
rect 158345 220902 166783 220904
rect 158345 220899 158411 220902
rect 166717 220899 166783 220902
rect 166901 220962 166967 220965
rect 175457 220962 175523 220965
rect 166901 220960 175523 220962
rect 166901 220904 166906 220960
rect 166962 220904 175462 220960
rect 175518 220904 175523 220960
rect 166901 220902 175523 220904
rect 166901 220899 166967 220902
rect 175457 220899 175523 220902
rect 497825 220962 497891 220965
rect 631317 220962 631383 220965
rect 497825 220960 631383 220962
rect 497825 220904 497830 220960
rect 497886 220904 631322 220960
rect 631378 220904 631383 220960
rect 497825 220902 631383 220904
rect 497825 220899 497891 220902
rect 631317 220899 631383 220902
rect 176469 220826 176535 220829
rect 179873 220826 179939 220829
rect 176469 220824 179939 220826
rect 176469 220768 176474 220824
rect 176530 220768 179878 220824
rect 179934 220768 179939 220824
rect 176469 220766 179939 220768
rect 176469 220763 176535 220766
rect 179873 220763 179939 220766
rect 563145 220690 563211 220693
rect 564801 220690 564867 220693
rect 653029 220690 653095 220693
rect 667841 220690 667907 220693
rect 563145 220688 564867 220690
rect 563145 220632 563150 220688
rect 563206 220632 564806 220688
rect 564862 220632 564867 220688
rect 563145 220630 564867 220632
rect 563145 220627 563211 220630
rect 564801 220627 564867 220630
rect 565310 220630 570338 220690
rect 151721 220554 151787 220557
rect 156965 220554 157031 220557
rect 151721 220552 157031 220554
rect 151721 220496 151726 220552
rect 151782 220496 156970 220552
rect 157026 220496 157031 220552
rect 151721 220494 157031 220496
rect 151721 220491 151787 220494
rect 156965 220491 157031 220494
rect 140773 220418 140839 220421
rect 142337 220418 142403 220421
rect 140773 220416 142403 220418
rect 140773 220360 140778 220416
rect 140834 220360 142342 220416
rect 142398 220360 142403 220416
rect 140773 220358 142403 220360
rect 140773 220355 140839 220358
rect 142337 220355 142403 220358
rect 144821 220418 144887 220421
rect 151445 220418 151511 220421
rect 553945 220418 554011 220421
rect 144821 220416 151511 220418
rect 144821 220360 144826 220416
rect 144882 220360 151450 220416
rect 151506 220360 151511 220416
rect 144821 220358 151511 220360
rect 144821 220355 144887 220358
rect 151445 220355 151511 220358
rect 553534 220416 554011 220418
rect 553534 220360 553950 220416
rect 554006 220360 554011 220416
rect 553534 220358 554011 220360
rect 166901 220282 166967 220285
rect 167085 220282 167151 220285
rect 166901 220280 167151 220282
rect 166901 220224 166906 220280
rect 166962 220224 167090 220280
rect 167146 220224 167151 220280
rect 166901 220222 167151 220224
rect 166901 220219 166967 220222
rect 167085 220219 167151 220222
rect 552841 220282 552907 220285
rect 553534 220282 553594 220358
rect 553945 220355 554011 220358
rect 563329 220418 563395 220421
rect 565310 220418 565370 220630
rect 563329 220416 565370 220418
rect 563329 220360 563334 220416
rect 563390 220360 565370 220416
rect 563329 220358 565370 220360
rect 565629 220418 565695 220421
rect 569953 220418 570019 220421
rect 565629 220416 570019 220418
rect 565629 220360 565634 220416
rect 565690 220360 569958 220416
rect 570014 220360 570019 220416
rect 565629 220358 570019 220360
rect 563329 220355 563395 220358
rect 565629 220355 565695 220358
rect 569953 220355 570019 220358
rect 552841 220280 553594 220282
rect 552841 220224 552846 220280
rect 552902 220224 553594 220280
rect 552841 220222 553594 220224
rect 570278 220282 570338 220630
rect 653029 220688 667907 220690
rect 653029 220632 653034 220688
rect 653090 220632 667846 220688
rect 667902 220632 667907 220688
rect 653029 220630 667907 220632
rect 653029 220627 653095 220630
rect 667841 220627 667907 220630
rect 675886 220628 675892 220692
rect 675956 220690 675962 220692
rect 675956 220630 676292 220690
rect 675956 220628 675962 220630
rect 572989 220554 573055 220557
rect 589641 220554 589707 220557
rect 675017 220554 675083 220557
rect 572989 220552 589707 220554
rect 572989 220496 572994 220552
rect 573050 220496 589646 220552
rect 589702 220496 589707 220552
rect 572989 220494 589707 220496
rect 572989 220491 573055 220494
rect 589641 220491 589707 220494
rect 669270 220552 675083 220554
rect 669270 220496 675022 220552
rect 675078 220496 675083 220552
rect 669270 220494 675083 220496
rect 572621 220418 572687 220421
rect 572805 220418 572871 220421
rect 572621 220416 572871 220418
rect 572621 220360 572626 220416
rect 572682 220360 572810 220416
rect 572866 220360 572871 220416
rect 572621 220358 572871 220360
rect 572621 220355 572687 220358
rect 572805 220355 572871 220358
rect 644749 220418 644815 220421
rect 669270 220418 669330 220494
rect 675017 220491 675083 220494
rect 644749 220416 669330 220418
rect 644749 220360 644754 220416
rect 644810 220360 669330 220416
rect 644749 220358 669330 220360
rect 644749 220355 644815 220358
rect 573357 220282 573423 220285
rect 586329 220282 586395 220285
rect 570278 220248 572546 220282
rect 573357 220280 586395 220282
rect 570278 220222 572730 220248
rect 552841 220219 552907 220222
rect 572486 220188 572730 220222
rect 573357 220224 573362 220280
rect 573418 220224 586334 220280
rect 586390 220224 586395 220280
rect 573357 220222 586395 220224
rect 573357 220219 573423 220222
rect 586329 220219 586395 220222
rect 672625 220282 672691 220285
rect 672625 220280 676292 220282
rect 672625 220224 672630 220280
rect 672686 220224 676292 220280
rect 672625 220222 676292 220224
rect 672625 220219 672691 220222
rect 142153 220146 142219 220149
rect 150893 220146 150959 220149
rect 142153 220144 150959 220146
rect 142153 220088 142158 220144
rect 142214 220088 150898 220144
rect 150954 220088 150959 220144
rect 142153 220086 150959 220088
rect 142153 220083 142219 220086
rect 150893 220083 150959 220086
rect 151077 220146 151143 220149
rect 151905 220146 151971 220149
rect 151077 220144 151971 220146
rect 151077 220088 151082 220144
rect 151138 220088 151910 220144
rect 151966 220088 151971 220144
rect 151077 220086 151971 220088
rect 151077 220083 151143 220086
rect 151905 220083 151971 220086
rect 180517 220146 180583 220149
rect 185761 220146 185827 220149
rect 180517 220144 185827 220146
rect 180517 220088 180522 220144
rect 180578 220088 185766 220144
rect 185822 220088 185827 220144
rect 180517 220086 185827 220088
rect 572670 220146 572730 220188
rect 572989 220146 573055 220149
rect 572670 220144 573055 220146
rect 572670 220088 572994 220144
rect 573050 220088 573055 220144
rect 572670 220086 573055 220088
rect 180517 220083 180583 220086
rect 185761 220083 185827 220086
rect 572989 220083 573055 220086
rect 562869 220010 562935 220013
rect 563513 220010 563579 220013
rect 562869 220008 563579 220010
rect 562869 219952 562874 220008
rect 562930 219952 563518 220008
rect 563574 219952 563579 220008
rect 562869 219950 563579 219952
rect 562869 219947 562935 219950
rect 563513 219947 563579 219950
rect 564801 220010 564867 220013
rect 572529 220010 572595 220013
rect 564801 220008 572595 220010
rect 564801 219952 564806 220008
rect 564862 219952 572534 220008
rect 572590 219952 572595 220008
rect 564801 219950 572595 219952
rect 564801 219947 564867 219950
rect 572529 219947 572595 219950
rect 586329 220010 586395 220013
rect 589457 220010 589523 220013
rect 586329 220008 589523 220010
rect 586329 219952 586334 220008
rect 586390 219952 589462 220008
rect 589518 219952 589523 220008
rect 586329 219950 589523 219952
rect 586329 219947 586395 219950
rect 589457 219947 589523 219950
rect 202413 219874 202479 219877
rect 203149 219874 203215 219877
rect 202413 219872 203215 219874
rect 202413 219816 202418 219872
rect 202474 219816 203154 219872
rect 203210 219816 203215 219872
rect 202413 219814 203215 219816
rect 202413 219811 202479 219814
rect 203149 219811 203215 219814
rect 683389 219874 683455 219877
rect 683389 219872 683468 219874
rect 683389 219816 683394 219872
rect 683450 219816 683468 219872
rect 683389 219814 683468 219816
rect 683389 219811 683455 219814
rect 141969 219738 142035 219741
rect 144177 219738 144243 219741
rect 141969 219736 144243 219738
rect 141969 219680 141974 219736
rect 142030 219680 144182 219736
rect 144238 219680 144243 219736
rect 141969 219678 144243 219680
rect 141969 219675 142035 219678
rect 144177 219675 144243 219678
rect 515213 219738 515279 219741
rect 617241 219738 617307 219741
rect 515213 219736 617307 219738
rect 515213 219680 515218 219736
rect 515274 219680 617246 219736
rect 617302 219680 617307 219736
rect 515213 219678 617307 219680
rect 515213 219675 515279 219678
rect 617241 219675 617307 219678
rect 668025 219738 668091 219741
rect 671337 219738 671403 219741
rect 668025 219736 671403 219738
rect 668025 219680 668030 219736
rect 668086 219680 671342 219736
rect 671398 219680 671403 219736
rect 668025 219678 671403 219680
rect 668025 219675 668091 219678
rect 671337 219675 671403 219678
rect 486969 219466 487035 219469
rect 611629 219466 611695 219469
rect 486969 219464 611695 219466
rect 486969 219408 486974 219464
rect 487030 219408 611634 219464
rect 611690 219408 611695 219464
rect 486969 219406 611695 219408
rect 486969 219403 487035 219406
rect 611629 219403 611695 219406
rect 667749 219466 667815 219469
rect 667749 219464 676292 219466
rect 667749 219408 667754 219464
rect 667810 219408 676292 219464
rect 667749 219406 676292 219408
rect 667749 219403 667815 219406
rect 553209 219194 553275 219197
rect 560201 219194 560267 219197
rect 553209 219192 560267 219194
rect 553209 219136 553214 219192
rect 553270 219136 560206 219192
rect 560262 219136 560267 219192
rect 553209 219134 560267 219136
rect 553209 219131 553275 219134
rect 560201 219131 560267 219134
rect 567101 219194 567167 219197
rect 568297 219194 568363 219197
rect 567101 219192 568363 219194
rect 567101 219136 567106 219192
rect 567162 219136 568302 219192
rect 568358 219136 568363 219192
rect 567101 219134 568363 219136
rect 567101 219131 567167 219134
rect 568297 219131 568363 219134
rect 672073 219058 672139 219061
rect 669270 219056 672139 219058
rect 669270 219000 672078 219056
rect 672134 219000 672139 219056
rect 669270 218998 672139 219000
rect 492673 218922 492739 218925
rect 493777 218922 493843 218925
rect 492673 218920 493843 218922
rect 492673 218864 492678 218920
rect 492734 218864 493782 218920
rect 493838 218864 493843 218920
rect 492673 218862 493843 218864
rect 492673 218859 492739 218862
rect 493777 218859 493843 218862
rect 494697 218922 494763 218925
rect 655421 218922 655487 218925
rect 669270 218922 669330 218998
rect 672073 218995 672139 218998
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 494697 218920 605850 218922
rect 494697 218864 494702 218920
rect 494758 218864 605850 218920
rect 494697 218862 605850 218864
rect 494697 218859 494763 218862
rect 171041 218650 171107 218653
rect 172881 218650 172947 218653
rect 171041 218648 172947 218650
rect 171041 218592 171046 218648
rect 171102 218592 172886 218648
rect 172942 218592 172947 218648
rect 171041 218590 172947 218592
rect 171041 218587 171107 218590
rect 172881 218587 172947 218590
rect 490373 218650 490439 218653
rect 497457 218650 497523 218653
rect 603349 218650 603415 218653
rect 490373 218648 493978 218650
rect 490373 218592 490378 218648
rect 490434 218592 493978 218648
rect 490373 218590 493978 218592
rect 490373 218587 490439 218590
rect 493918 218378 493978 218590
rect 497457 218648 603415 218650
rect 497457 218592 497462 218648
rect 497518 218592 603354 218648
rect 603410 218592 603415 218648
rect 497457 218590 603415 218592
rect 605790 218650 605850 218862
rect 655421 218920 669330 218922
rect 655421 218864 655426 218920
rect 655482 218864 669330 218920
rect 655421 218862 669330 218864
rect 655421 218859 655487 218862
rect 631133 218650 631199 218653
rect 605790 218648 631199 218650
rect 605790 218592 631138 218648
rect 631194 218592 631199 218648
rect 605790 218590 631199 218592
rect 497457 218587 497523 218590
rect 603349 218587 603415 218590
rect 631133 218587 631199 218590
rect 648521 218650 648587 218653
rect 675109 218650 675175 218653
rect 683297 218650 683363 218653
rect 648521 218648 675175 218650
rect 648521 218592 648526 218648
rect 648582 218592 675114 218648
rect 675170 218592 675175 218648
rect 648521 218590 675175 218592
rect 683284 218648 683363 218650
rect 683284 218592 683302 218648
rect 683358 218592 683363 218648
rect 683284 218590 683363 218592
rect 648521 218587 648587 218590
rect 675109 218587 675175 218590
rect 683297 218587 683363 218590
rect 594793 218378 594859 218381
rect 493918 218376 594859 218378
rect 493918 218320 594798 218376
rect 594854 218320 594859 218376
rect 493918 218318 594859 218320
rect 594793 218315 594859 218318
rect 675886 218180 675892 218244
rect 675956 218242 675962 218244
rect 675956 218182 676292 218242
rect 675956 218180 675962 218182
rect 487797 218106 487863 218109
rect 627453 218106 627519 218109
rect 487797 218104 627519 218106
rect 487797 218048 487802 218104
rect 487858 218048 627458 218104
rect 627514 218048 627519 218104
rect 487797 218046 627519 218048
rect 487797 218043 487863 218046
rect 627453 218043 627519 218046
rect 35801 217970 35867 217973
rect 61285 217970 61351 217973
rect 35801 217968 61351 217970
rect 35801 217912 35806 217968
rect 35862 217912 61290 217968
rect 61346 217912 61351 217968
rect 35801 217910 61351 217912
rect 35801 217907 35867 217910
rect 61285 217907 61351 217910
rect 508497 217834 508563 217837
rect 510153 217836 510219 217837
rect 509182 217834 509188 217836
rect 508497 217832 509188 217834
rect 508497 217776 508502 217832
rect 508558 217776 509188 217832
rect 508497 217774 509188 217776
rect 508497 217771 508563 217774
rect 509182 217772 509188 217774
rect 509252 217772 509258 217836
rect 510102 217834 510108 217836
rect 510062 217774 510108 217834
rect 510172 217832 510219 217836
rect 522573 217836 522639 217837
rect 522573 217834 522620 217836
rect 510214 217776 510219 217832
rect 510102 217772 510108 217774
rect 510172 217772 510219 217776
rect 522528 217832 522620 217834
rect 522528 217776 522578 217832
rect 522528 217774 522620 217776
rect 510153 217771 510219 217772
rect 522573 217772 522620 217774
rect 522684 217772 522690 217836
rect 555693 217834 555759 217837
rect 562685 217834 562751 217837
rect 555693 217832 562751 217834
rect 555693 217776 555698 217832
rect 555754 217776 562690 217832
rect 562746 217776 562751 217832
rect 555693 217774 562751 217776
rect 522573 217771 522639 217772
rect 555693 217771 555759 217774
rect 562685 217771 562751 217774
rect 562869 217834 562935 217837
rect 563513 217834 563579 217837
rect 566917 217836 566983 217837
rect 566917 217834 566964 217836
rect 562869 217832 563579 217834
rect 562869 217776 562874 217832
rect 562930 217776 563518 217832
rect 563574 217776 563579 217832
rect 562869 217774 563579 217776
rect 566872 217832 566964 217834
rect 566872 217776 566922 217832
rect 566872 217774 566964 217776
rect 562869 217771 562935 217774
rect 563513 217771 563579 217774
rect 566917 217772 566964 217774
rect 567028 217772 567034 217836
rect 572069 217834 572135 217837
rect 574093 217834 574159 217837
rect 572069 217832 574159 217834
rect 572069 217776 572074 217832
rect 572130 217776 574098 217832
rect 574154 217776 574159 217832
rect 572069 217774 574159 217776
rect 566917 217771 566983 217772
rect 572069 217771 572135 217774
rect 574093 217771 574159 217774
rect 574318 217772 574324 217836
rect 574388 217834 574394 217836
rect 574829 217834 574895 217837
rect 574388 217832 574895 217834
rect 574388 217776 574834 217832
rect 574890 217776 574895 217832
rect 574388 217774 574895 217776
rect 574388 217772 574394 217774
rect 574829 217771 574895 217774
rect 675017 217834 675083 217837
rect 675017 217832 676292 217834
rect 675017 217776 675022 217832
rect 675078 217776 676292 217832
rect 675017 217774 676292 217776
rect 675017 217771 675083 217774
rect 505645 217562 505711 217565
rect 595161 217562 595227 217565
rect 505645 217560 595227 217562
rect 505645 217504 505650 217560
rect 505706 217504 595166 217560
rect 595222 217504 595227 217560
rect 505645 217502 595227 217504
rect 505645 217499 505711 217502
rect 595161 217499 595227 217502
rect 662045 217562 662111 217565
rect 675569 217562 675635 217565
rect 662045 217560 675635 217562
rect 662045 217504 662050 217560
rect 662106 217504 675574 217560
rect 675630 217504 675635 217560
rect 662045 217502 675635 217504
rect 662045 217499 662111 217502
rect 675569 217499 675635 217502
rect 675702 217364 675708 217428
rect 675772 217426 675778 217428
rect 675772 217366 676292 217426
rect 675772 217364 675778 217366
rect 493777 217292 493843 217293
rect 493726 217228 493732 217292
rect 493796 217290 493843 217292
rect 495341 217290 495407 217293
rect 498561 217290 498627 217293
rect 596357 217290 596423 217293
rect 493796 217288 493888 217290
rect 493838 217232 493888 217288
rect 493796 217230 493888 217232
rect 495341 217288 495450 217290
rect 495341 217232 495346 217288
rect 495402 217232 495450 217288
rect 493796 217228 493843 217230
rect 493777 217227 493843 217228
rect 495341 217227 495450 217232
rect 498561 217288 596423 217290
rect 498561 217232 498566 217288
rect 498622 217232 596362 217288
rect 596418 217232 596423 217288
rect 498561 217230 596423 217232
rect 498561 217227 498627 217230
rect 596357 217227 596423 217230
rect 656801 217290 656867 217293
rect 672441 217290 672507 217293
rect 656801 217288 672507 217290
rect 656801 217232 656806 217288
rect 656862 217232 672446 217288
rect 672502 217232 672507 217288
rect 656801 217230 672507 217232
rect 656801 217227 656867 217230
rect 672441 217227 672507 217230
rect 488671 217154 488737 217157
rect 488671 217152 489930 217154
rect 488671 217096 488676 217152
rect 488732 217096 489930 217152
rect 488671 217094 489930 217096
rect 488671 217091 488737 217094
rect 489870 216746 489930 217094
rect 495390 217018 495450 217227
rect 600773 217154 600839 217157
rect 601509 217154 601575 217157
rect 600773 217152 601575 217154
rect 600773 217096 600778 217152
rect 600834 217096 601514 217152
rect 601570 217096 601575 217152
rect 600773 217094 601575 217096
rect 600773 217091 600839 217094
rect 601509 217091 601575 217094
rect 595713 217018 595779 217021
rect 495390 217016 595779 217018
rect 495390 216960 595718 217016
rect 595774 216960 595779 217016
rect 495390 216958 595779 216960
rect 595713 216955 595779 216958
rect 674649 217018 674715 217021
rect 674649 217016 676292 217018
rect 674649 216960 674654 217016
rect 674710 216960 676292 217016
rect 674649 216958 676292 216960
rect 674649 216955 674715 216958
rect 574093 216746 574159 216749
rect 489870 216744 574159 216746
rect 489870 216688 574098 216744
rect 574154 216688 574159 216744
rect 489870 216686 574159 216688
rect 574093 216683 574159 216686
rect 574318 216684 574324 216748
rect 574388 216746 574394 216748
rect 574645 216746 574711 216749
rect 574388 216744 574711 216746
rect 574388 216688 574650 216744
rect 574706 216688 574711 216744
rect 574388 216686 574711 216688
rect 574388 216684 574394 216686
rect 574645 216683 574711 216686
rect 671889 216610 671955 216613
rect 671889 216608 676292 216610
rect 671889 216552 671894 216608
rect 671950 216552 676292 216608
rect 671889 216550 676292 216552
rect 671889 216547 671955 216550
rect 674373 216338 674439 216341
rect 669270 216336 674439 216338
rect 669270 216280 674378 216336
rect 674434 216280 674439 216336
rect 669270 216278 674439 216280
rect 566958 216140 566964 216204
rect 567028 216202 567034 216204
rect 627913 216202 627979 216205
rect 567028 216200 627979 216202
rect 567028 216144 627918 216200
rect 627974 216144 627979 216200
rect 567028 216142 627979 216144
rect 567028 216140 567034 216142
rect 627913 216139 627979 216142
rect 665541 216202 665607 216205
rect 669270 216202 669330 216278
rect 674373 216275 674439 216278
rect 665541 216200 669330 216202
rect 665541 216144 665546 216200
rect 665602 216144 669330 216200
rect 665541 216142 669330 216144
rect 674833 216202 674899 216205
rect 674833 216200 676292 216202
rect 674833 216144 674838 216200
rect 674894 216144 676292 216200
rect 674833 216142 676292 216144
rect 665541 216139 665607 216142
rect 674833 216139 674899 216142
rect 673453 216066 673519 216069
rect 669454 216064 673519 216066
rect 669454 216008 673458 216064
rect 673514 216008 673519 216064
rect 669454 216006 673519 216008
rect 509182 215868 509188 215932
rect 509252 215930 509258 215932
rect 598473 215930 598539 215933
rect 509252 215928 598539 215930
rect 509252 215872 598478 215928
rect 598534 215872 598539 215928
rect 509252 215870 598539 215872
rect 509252 215868 509258 215870
rect 598473 215867 598539 215870
rect 652845 215930 652911 215933
rect 669454 215930 669514 216006
rect 673453 216003 673519 216006
rect 652845 215928 669514 215930
rect 652845 215872 652850 215928
rect 652906 215872 669514 215928
rect 652845 215870 669514 215872
rect 652845 215867 652911 215870
rect 673177 215794 673243 215797
rect 673177 215792 676292 215794
rect 673177 215736 673182 215792
rect 673238 215736 676292 215792
rect 673177 215734 676292 215736
rect 673177 215731 673243 215734
rect 674373 215522 674439 215525
rect 675937 215522 676003 215525
rect 674373 215520 676003 215522
rect 674373 215464 674378 215520
rect 674434 215464 675942 215520
rect 675998 215464 676003 215520
rect 674373 215462 676003 215464
rect 674373 215459 674439 215462
rect 675937 215459 676003 215462
rect 522614 215324 522620 215388
rect 522684 215386 522690 215388
rect 618897 215386 618963 215389
rect 522684 215384 618963 215386
rect 522684 215328 618902 215384
rect 618958 215328 618963 215384
rect 522684 215326 618963 215328
rect 522684 215324 522690 215326
rect 618897 215323 618963 215326
rect 676262 215310 676322 215356
rect 673637 215252 673703 215253
rect 673637 215248 673684 215252
rect 673748 215250 673754 215252
rect 673637 215192 673642 215248
rect 673637 215188 673684 215192
rect 673748 215190 673794 215250
rect 673748 215188 673754 215190
rect 675886 215188 675892 215252
rect 675956 215250 675962 215252
rect 676078 215250 676322 215310
rect 675956 215190 676138 215250
rect 675956 215188 675962 215190
rect 673637 215187 673703 215188
rect 663750 215054 669330 215114
rect 47761 214978 47827 214981
rect 41492 214976 47827 214978
rect 41492 214920 47766 214976
rect 47822 214920 47827 214976
rect 41492 214918 47827 214920
rect 47761 214915 47827 214918
rect 35801 214706 35867 214709
rect 35758 214704 35867 214706
rect 35758 214648 35806 214704
rect 35862 214648 35867 214704
rect 35758 214643 35867 214648
rect 35758 214540 35818 214643
rect 658733 214570 658799 214573
rect 663750 214570 663810 215054
rect 669270 214706 669330 215054
rect 673637 214978 673703 214981
rect 673637 214976 676292 214978
rect 673637 214920 673642 214976
rect 673698 214920 676292 214976
rect 673637 214918 676292 214920
rect 673637 214915 673703 214918
rect 675937 214706 676003 214709
rect 669270 214704 676003 214706
rect 669270 214648 675942 214704
rect 675998 214648 676003 214704
rect 669270 214646 676003 214648
rect 675937 214643 676003 214646
rect 658733 214568 663810 214570
rect 658733 214512 658738 214568
rect 658794 214512 663810 214568
rect 658733 214510 663810 214512
rect 676170 214510 676292 214570
rect 658733 214507 658799 214510
rect 35801 214298 35867 214301
rect 35758 214296 35867 214298
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214235 35867 214240
rect 35758 214132 35818 214235
rect 575982 214026 576042 214404
rect 675886 214372 675892 214436
rect 675956 214434 675962 214436
rect 676170 214434 676230 214510
rect 675956 214374 676230 214434
rect 675956 214372 675962 214374
rect 674465 214162 674531 214165
rect 674465 214160 676292 214162
rect 674465 214104 674470 214160
rect 674526 214104 676292 214160
rect 674465 214102 676292 214104
rect 674465 214099 674531 214102
rect 578877 214026 578943 214029
rect 674097 214026 674163 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 666510 214024 674163 214026
rect 666510 213968 674102 214024
rect 674158 213968 674163 214024
rect 666510 213966 674163 213968
rect 44817 213754 44883 213757
rect 666510 213754 666570 213966
rect 674097 213963 674163 213966
rect 41492 213752 44883 213754
rect 41492 213696 44822 213752
rect 44878 213696 44883 213752
rect 41492 213694 44883 213696
rect 44817 213691 44883 213694
rect 663750 213694 666570 213754
rect 672533 213754 672599 213757
rect 672533 213752 676292 213754
rect 672533 213696 672538 213752
rect 672594 213696 676292 213752
rect 672533 213694 676292 213696
rect 661493 213482 661559 213485
rect 663750 213482 663810 213694
rect 672533 213691 672599 213694
rect 661493 213480 663810 213482
rect 661493 213424 661498 213480
rect 661554 213424 663810 213480
rect 661493 213422 663810 213424
rect 661493 213419 661559 213422
rect 47761 213346 47827 213349
rect 41492 213344 47827 213346
rect 41492 213288 47766 213344
rect 47822 213288 47827 213344
rect 41492 213286 47827 213288
rect 47761 213283 47827 213286
rect 672717 213346 672783 213349
rect 672717 213344 676292 213346
rect 672717 213288 672722 213344
rect 672778 213288 676292 213344
rect 672717 213286 676292 213288
rect 672717 213283 672783 213286
rect 656525 213210 656591 213213
rect 668025 213210 668091 213213
rect 656525 213208 668091 213210
rect 656525 213152 656530 213208
rect 656586 213152 668030 213208
rect 668086 213152 668091 213208
rect 656525 213150 668091 213152
rect 656525 213147 656591 213150
rect 668025 213147 668091 213150
rect 45553 212938 45619 212941
rect 683113 212938 683179 212941
rect 41492 212936 45619 212938
rect 41492 212880 45558 212936
rect 45614 212880 45619 212936
rect 682916 212936 683179 212938
rect 682916 212908 683118 212936
rect 41492 212878 45619 212880
rect 45553 212875 45619 212878
rect 682886 212880 683118 212908
rect 683174 212880 683179 212936
rect 682886 212878 683179 212880
rect 674005 212802 674071 212805
rect 674230 212802 674236 212804
rect 674005 212800 674236 212802
rect 674005 212744 674010 212800
rect 674066 212744 674236 212800
rect 674005 212742 674236 212744
rect 674005 212739 674071 212742
rect 674230 212740 674236 212742
rect 674300 212740 674306 212804
rect 682886 212500 682946 212878
rect 683113 212875 683179 212878
rect 35390 212261 35450 212500
rect 35390 212256 35499 212261
rect 35390 212200 35438 212256
rect 35494 212200 35499 212256
rect 35390 212198 35499 212200
rect 35433 212195 35499 212198
rect 44633 212122 44699 212125
rect 41492 212120 44699 212122
rect 41492 212064 44638 212120
rect 44694 212064 44699 212120
rect 41492 212062 44699 212064
rect 44633 212059 44699 212062
rect 35617 211850 35683 211853
rect 35574 211848 35683 211850
rect 35574 211792 35622 211848
rect 35678 211792 35683 211848
rect 35574 211787 35683 211792
rect 39573 211850 39639 211853
rect 42793 211850 42859 211853
rect 39573 211848 42859 211850
rect 39573 211792 39578 211848
rect 39634 211792 42798 211848
rect 42854 211792 42859 211848
rect 39573 211790 42859 211792
rect 39573 211787 39639 211790
rect 42793 211787 42859 211790
rect 35574 211684 35634 211787
rect 575982 211714 576042 212228
rect 675845 212122 675911 212125
rect 675845 212120 676292 212122
rect 675845 212064 675850 212120
rect 675906 212064 676292 212120
rect 675845 212062 676292 212064
rect 675845 212059 675911 212062
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 679022 211445 679082 211684
rect 35801 211442 35867 211445
rect 35758 211440 35867 211442
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211379 35867 211384
rect 678973 211440 679082 211445
rect 678973 211384 678978 211440
rect 679034 211384 679082 211440
rect 678973 211382 679082 211384
rect 678973 211379 679039 211382
rect 35758 211276 35818 211379
rect 47945 210898 48011 210901
rect 41492 210896 48011 210898
rect 41492 210840 47950 210896
rect 48006 210840 48011 210896
rect 41492 210838 48011 210840
rect 47945 210835 48011 210838
rect 676254 210836 676260 210900
rect 676324 210898 676330 210900
rect 676622 210898 676628 210900
rect 676324 210838 676628 210898
rect 676324 210836 676330 210838
rect 676622 210836 676628 210838
rect 676692 210836 676698 210900
rect 675886 210564 675892 210628
rect 675956 210626 675962 210628
rect 680353 210626 680419 210629
rect 675956 210624 680419 210626
rect 675956 210568 680358 210624
rect 680414 210568 680419 210624
rect 675956 210566 680419 210568
rect 675956 210564 675962 210566
rect 680353 210563 680419 210566
rect 670785 210492 670851 210493
rect 670734 210490 670740 210492
rect 35758 210221 35818 210460
rect 670694 210430 670740 210490
rect 670804 210488 670851 210492
rect 670846 210432 670851 210488
rect 670734 210428 670740 210430
rect 670804 210428 670851 210432
rect 670785 210427 670851 210428
rect 683297 210354 683363 210357
rect 678930 210352 683363 210354
rect 678930 210296 683302 210352
rect 683358 210296 683363 210352
rect 678930 210294 683363 210296
rect 35758 210216 35867 210221
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35758 210158 35867 210160
rect 35801 210155 35867 210158
rect 41822 210082 41828 210084
rect 41492 210022 41828 210082
rect 41822 210020 41828 210022
rect 41892 210020 41898 210084
rect 575982 209810 576042 210052
rect 670785 209946 670851 209949
rect 678930 209946 678990 210294
rect 683297 210291 683363 210294
rect 670785 209944 678990 209946
rect 670785 209888 670790 209944
rect 670846 209888 678990 209944
rect 670785 209886 678990 209888
rect 670785 209883 670851 209886
rect 579521 209810 579587 209813
rect 575982 209808 579587 209810
rect 575982 209752 579526 209808
rect 579582 209752 579587 209808
rect 575982 209750 579587 209752
rect 579521 209747 579587 209750
rect 46933 209674 46999 209677
rect 41492 209672 46999 209674
rect 41492 209616 46938 209672
rect 46994 209616 46999 209672
rect 41492 209614 46999 209616
rect 46933 209611 46999 209614
rect 674097 209674 674163 209677
rect 675845 209674 675911 209677
rect 674097 209672 675911 209674
rect 674097 209616 674102 209672
rect 674158 209616 675850 209672
rect 675906 209616 675911 209672
rect 674097 209614 675911 209616
rect 674097 209611 674163 209614
rect 675845 209611 675911 209614
rect 35574 208997 35634 209236
rect 35574 208992 35683 208997
rect 35574 208936 35622 208992
rect 35678 208936 35683 208992
rect 35574 208934 35683 208936
rect 35617 208931 35683 208934
rect 35758 208589 35818 208828
rect 35758 208584 35867 208589
rect 35758 208528 35806 208584
rect 35862 208528 35867 208584
rect 35758 208526 35867 208528
rect 35801 208523 35867 208526
rect 44357 208450 44423 208453
rect 41492 208448 44423 208450
rect 41492 208392 44362 208448
rect 44418 208392 44423 208448
rect 41492 208390 44423 208392
rect 44357 208387 44423 208390
rect 40033 208178 40099 208181
rect 41454 208178 41460 208180
rect 40033 208176 41460 208178
rect 40033 208120 40038 208176
rect 40094 208120 41460 208176
rect 40033 208118 41460 208120
rect 40033 208115 40099 208118
rect 41454 208116 41460 208118
rect 41524 208116 41530 208180
rect 41689 208178 41755 208181
rect 49509 208178 49575 208181
rect 41689 208176 49575 208178
rect 41689 208120 41694 208176
rect 41750 208120 49514 208176
rect 49570 208120 49575 208176
rect 41689 208118 49575 208120
rect 41689 208115 41755 208118
rect 49509 208115 49575 208118
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 35758 207773 35818 208012
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 35758 207768 35867 207773
rect 35758 207712 35806 207768
rect 35862 207712 35867 207768
rect 35758 207710 35867 207712
rect 35801 207707 35867 207710
rect 40493 207770 40559 207773
rect 42977 207770 43043 207773
rect 40493 207768 43043 207770
rect 40493 207712 40498 207768
rect 40554 207712 42982 207768
rect 43038 207712 43043 207768
rect 40493 207710 43043 207712
rect 40493 207707 40559 207710
rect 42977 207707 43043 207710
rect 40542 207364 40602 207604
rect 575982 207498 576042 207876
rect 668025 207634 668091 207637
rect 678973 207634 679039 207637
rect 668025 207632 679039 207634
rect 668025 207576 668030 207632
rect 668086 207576 678978 207632
rect 679034 207576 679039 207632
rect 668025 207574 679039 207576
rect 668025 207571 668091 207574
rect 678973 207571 679039 207574
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40534 207300 40540 207364
rect 40604 207300 40610 207364
rect 44173 207226 44239 207229
rect 41492 207224 44239 207226
rect 41492 207168 44178 207224
rect 44234 207168 44239 207224
rect 41492 207166 44239 207168
rect 44173 207163 44239 207166
rect 676070 206892 676076 206956
rect 676140 206954 676146 206956
rect 676857 206954 676923 206957
rect 676140 206952 676923 206954
rect 676140 206896 676862 206952
rect 676918 206896 676923 206952
rect 676140 206894 676923 206896
rect 676140 206892 676146 206894
rect 676857 206891 676923 206894
rect 40726 206548 40786 206788
rect 40718 206484 40724 206548
rect 40788 206484 40794 206548
rect 41321 206546 41387 206549
rect 48773 206546 48839 206549
rect 41321 206544 48839 206546
rect 41321 206488 41326 206544
rect 41382 206488 48778 206544
rect 48834 206488 48839 206544
rect 41321 206486 48839 206488
rect 41321 206483 41387 206486
rect 48773 206483 48839 206486
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 35801 206138 35867 206141
rect 40910 206140 40970 206380
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 35758 206136 35867 206138
rect 35758 206080 35806 206136
rect 35862 206080 35867 206136
rect 35758 206075 35867 206080
rect 40902 206076 40908 206140
rect 40972 206076 40978 206140
rect 35758 205972 35818 206075
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 40217 205730 40283 205733
rect 41638 205730 41644 205732
rect 40217 205728 41644 205730
rect 40217 205672 40222 205728
rect 40278 205672 41644 205728
rect 40217 205670 41644 205672
rect 40217 205667 40283 205670
rect 41638 205668 41644 205670
rect 41708 205668 41714 205732
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 675753 205594 675819 205597
rect 676438 205594 676444 205596
rect 675753 205592 676444 205594
rect 41462 205322 41522 205564
rect 675753 205536 675758 205592
rect 675814 205536 676444 205592
rect 675753 205534 676444 205536
rect 675753 205531 675819 205534
rect 676438 205532 676444 205534
rect 676508 205532 676514 205596
rect 44633 205322 44699 205325
rect 41462 205320 44699 205322
rect 41462 205264 44638 205320
rect 44694 205264 44699 205320
rect 41462 205262 44699 205264
rect 44633 205259 44699 205262
rect 35574 204917 35634 205156
rect 35574 204912 35683 204917
rect 44817 204914 44883 204917
rect 35574 204856 35622 204912
rect 35678 204856 35683 204912
rect 35574 204854 35683 204856
rect 35617 204851 35683 204854
rect 41462 204912 44883 204914
rect 41462 204856 44822 204912
rect 44878 204856 44883 204912
rect 41462 204854 44883 204856
rect 41462 204748 41522 204854
rect 44817 204851 44883 204854
rect 589457 204778 589523 204781
rect 589457 204776 592572 204778
rect 589457 204720 589462 204776
rect 589518 204720 592572 204776
rect 589457 204718 592572 204720
rect 589457 204715 589523 204718
rect 40953 204506 41019 204509
rect 43161 204506 43227 204509
rect 40953 204504 43227 204506
rect 40953 204448 40958 204504
rect 41014 204448 43166 204504
rect 43222 204448 43227 204504
rect 40953 204446 43227 204448
rect 40953 204443 41019 204446
rect 43161 204443 43227 204446
rect 671889 204506 671955 204509
rect 675109 204506 675175 204509
rect 671889 204504 675175 204506
rect 671889 204448 671894 204504
rect 671950 204448 675114 204504
rect 675170 204448 675175 204504
rect 671889 204446 675175 204448
rect 671889 204443 671955 204446
rect 675109 204443 675175 204446
rect 43345 204370 43411 204373
rect 43989 204370 44055 204373
rect 43345 204368 44055 204370
rect 35758 204101 35818 204340
rect 43345 204312 43350 204368
rect 43406 204312 43994 204368
rect 44050 204312 44055 204368
rect 43345 204310 44055 204312
rect 43345 204307 43411 204310
rect 43989 204307 44055 204310
rect 675753 204234 675819 204237
rect 676070 204234 676076 204236
rect 675753 204232 676076 204234
rect 675753 204176 675758 204232
rect 675814 204176 676076 204232
rect 675753 204174 676076 204176
rect 675753 204171 675819 204174
rect 676070 204172 676076 204174
rect 676140 204172 676146 204236
rect 35758 204096 35867 204101
rect 35758 204040 35806 204096
rect 35862 204040 35867 204096
rect 35758 204038 35867 204040
rect 35801 204035 35867 204038
rect 40401 204098 40467 204101
rect 43805 204098 43871 204101
rect 668025 204098 668091 204101
rect 40401 204096 43871 204098
rect 40401 204040 40406 204096
rect 40462 204040 43810 204096
rect 43866 204040 43871 204096
rect 40401 204038 43871 204040
rect 40401 204035 40467 204038
rect 43805 204035 43871 204038
rect 666694 204096 668091 204098
rect 666694 204040 668030 204096
rect 668086 204040 668091 204096
rect 666694 204038 668091 204040
rect 666694 204030 666754 204038
rect 668025 204035 668091 204038
rect 666356 203970 666754 204030
rect 28582 203693 28642 203932
rect 28533 203688 28642 203693
rect 28533 203632 28538 203688
rect 28594 203632 28642 203688
rect 28533 203630 28642 203632
rect 28533 203627 28599 203630
rect 46197 203554 46263 203557
rect 41492 203552 46263 203554
rect 41492 203496 46202 203552
rect 46258 203496 46263 203552
rect 41492 203494 46263 203496
rect 46197 203491 46263 203494
rect 40769 203282 40835 203285
rect 42793 203282 42859 203285
rect 40769 203280 42859 203282
rect 40769 203224 40774 203280
rect 40830 203224 42798 203280
rect 42854 203224 42859 203280
rect 40769 203222 42859 203224
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 40769 203219 40835 203222
rect 42793 203219 42859 203222
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 673085 201378 673151 201381
rect 675109 201378 675175 201381
rect 673085 201376 675175 201378
rect 575982 200834 576042 201348
rect 673085 201320 673090 201376
rect 673146 201320 675114 201376
rect 675170 201320 675175 201376
rect 673085 201318 675175 201320
rect 673085 201315 673151 201318
rect 675109 201315 675175 201318
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 674465 200834 674531 200837
rect 675293 200834 675359 200837
rect 674465 200832 675359 200834
rect 674465 200776 674470 200832
rect 674526 200776 675298 200832
rect 675354 200776 675359 200832
rect 674465 200774 675359 200776
rect 674465 200771 674531 200774
rect 675293 200771 675359 200774
rect 675753 200698 675819 200701
rect 676254 200698 676260 200700
rect 675753 200696 676260 200698
rect 675753 200640 675758 200696
rect 675814 200640 676260 200696
rect 675753 200638 676260 200640
rect 675753 200635 675819 200638
rect 676254 200636 676260 200638
rect 676324 200636 676330 200700
rect 673637 200562 673703 200565
rect 675109 200562 675175 200565
rect 673637 200560 675175 200562
rect 673637 200504 673642 200560
rect 673698 200504 675114 200560
rect 675170 200504 675175 200560
rect 673637 200502 675175 200504
rect 673637 200499 673703 200502
rect 675109 200499 675175 200502
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 28533 199338 28599 199341
rect 42241 199338 42307 199341
rect 28533 199336 42307 199338
rect 28533 199280 28538 199336
rect 28594 199280 42246 199336
rect 42302 199280 42307 199336
rect 28533 199278 42307 199280
rect 28533 199275 28599 199278
rect 42241 199275 42307 199278
rect 667933 199202 667999 199205
rect 666694 199200 667999 199202
rect 575982 198930 576042 199172
rect 666694 199144 667938 199200
rect 667994 199144 667999 199200
rect 666694 199142 667999 199144
rect 666694 199134 666754 199142
rect 667933 199139 667999 199142
rect 666356 199074 666754 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 675753 198388 675819 198389
rect 675702 198386 675708 198388
rect 675662 198326 675708 198386
rect 675772 198384 675819 198388
rect 675814 198328 675819 198384
rect 675702 198324 675708 198326
rect 675772 198324 675819 198328
rect 675753 198323 675819 198324
rect 590377 198250 590443 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 590377 198187 590443 198190
rect 42057 197026 42123 197029
rect 44357 197026 44423 197029
rect 42057 197024 44423 197026
rect 42057 196968 42062 197024
rect 42118 196968 44362 197024
rect 44418 196968 44423 197024
rect 42057 196966 44423 196968
rect 42057 196963 42123 196966
rect 44357 196963 44423 196966
rect 49509 196482 49575 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49509 196480 52164 196482
rect 49509 196424 49514 196480
rect 49570 196424 52164 196480
rect 49509 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49509 196419 49575 196422
rect 578509 196419 578575 196422
rect 672533 196346 672599 196349
rect 675109 196346 675175 196349
rect 672533 196344 675175 196346
rect 672533 196288 672538 196344
rect 672594 196288 675114 196344
rect 675170 196288 675175 196344
rect 672533 196286 675175 196288
rect 672533 196283 672599 196286
rect 675109 196283 675175 196286
rect 676622 196074 676628 196076
rect 675296 196014 676628 196074
rect 675296 195805 675356 196014
rect 676622 196012 676628 196014
rect 676692 196012 676698 196076
rect 675293 195800 675359 195805
rect 675293 195744 675298 195800
rect 675354 195744 675359 195800
rect 675293 195739 675359 195744
rect 41873 195260 41939 195261
rect 41822 195258 41828 195260
rect 41782 195198 41828 195258
rect 41892 195256 41939 195260
rect 41934 195200 41939 195256
rect 41822 195196 41828 195198
rect 41892 195196 41939 195200
rect 41873 195195 41939 195196
rect 40902 194924 40908 194988
rect 40972 194986 40978 194988
rect 42241 194986 42307 194989
rect 579521 194986 579587 194989
rect 40972 194984 42307 194986
rect 40972 194928 42246 194984
rect 42302 194928 42307 194984
rect 40972 194926 42307 194928
rect 40972 194924 40978 194926
rect 42241 194923 42307 194926
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 48313 194442 48379 194445
rect 48313 194440 52164 194442
rect 48313 194384 48318 194440
rect 48374 194384 52164 194440
rect 48313 194382 52164 194384
rect 48313 194379 48379 194382
rect 666356 194178 666754 194238
rect 666694 194170 666754 194178
rect 667933 194170 667999 194173
rect 666694 194168 667999 194170
rect 666694 194112 667938 194168
rect 667994 194112 667999 194168
rect 666694 194110 667999 194112
rect 667933 194107 667999 194110
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 40718 193156 40724 193220
rect 40788 193218 40794 193220
rect 41781 193218 41847 193221
rect 40788 193216 41847 193218
rect 40788 193160 41786 193216
rect 41842 193160 41847 193216
rect 40788 193158 41847 193160
rect 40788 193156 40794 193158
rect 41781 193155 41847 193158
rect 670785 193218 670851 193221
rect 675109 193218 675175 193221
rect 670785 193216 675175 193218
rect 670785 193160 670790 193216
rect 670846 193160 675114 193216
rect 675170 193160 675175 193216
rect 670785 193158 675175 193160
rect 670785 193155 670851 193158
rect 675109 193155 675175 193158
rect 675661 192674 675727 192677
rect 675886 192674 675892 192676
rect 675661 192672 675892 192674
rect 48773 192402 48839 192405
rect 48773 192400 52164 192402
rect 48773 192344 48778 192400
rect 48834 192344 52164 192400
rect 48773 192342 52164 192344
rect 48773 192339 48839 192342
rect 575982 192266 576042 192644
rect 675661 192616 675666 192672
rect 675722 192616 675892 192672
rect 675661 192614 675892 192616
rect 675661 192611 675727 192614
rect 675886 192612 675892 192614
rect 675956 192612 675962 192676
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 42057 191586 42123 191589
rect 43989 191586 44055 191589
rect 42057 191584 44055 191586
rect 42057 191528 42062 191584
rect 42118 191528 43994 191584
rect 44050 191528 44055 191584
rect 42057 191526 44055 191528
rect 42057 191523 42123 191526
rect 43989 191523 44055 191526
rect 42241 190906 42307 190909
rect 44633 190906 44699 190909
rect 42241 190904 44699 190906
rect 42241 190848 42246 190904
rect 42302 190848 44638 190904
rect 44694 190848 44699 190904
rect 42241 190846 44699 190848
rect 42241 190843 42307 190846
rect 44633 190843 44699 190846
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 47761 190498 47827 190501
rect 47761 190496 52164 190498
rect 47761 190440 47766 190496
rect 47822 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 47761 190438 52164 190440
rect 47761 190435 47827 190438
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 667933 189682 667999 189685
rect 676857 189682 676923 189685
rect 666878 189680 676923 189682
rect 666878 189624 667938 189680
rect 667994 189624 676862 189680
rect 676918 189624 676923 189680
rect 666878 189622 676923 189624
rect 666878 189342 666938 189622
rect 667933 189619 667999 189622
rect 676857 189619 676923 189622
rect 666356 189282 666938 189342
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 186826 42491 186829
rect 44173 186826 44239 186829
rect 42425 186824 44239 186826
rect 42425 186768 42430 186824
rect 42486 186768 44178 186824
rect 44234 186768 44239 186824
rect 42425 186766 44239 186768
rect 42425 186763 42491 186766
rect 44173 186763 44239 186766
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 40534 186356 40540 186420
rect 40604 186418 40610 186420
rect 41781 186418 41847 186421
rect 40604 186416 41847 186418
rect 40604 186360 41786 186416
rect 41842 186360 41847 186416
rect 40604 186358 41847 186360
rect 40604 186356 40610 186358
rect 41781 186355 41847 186358
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 41454 185948 41460 186012
rect 41524 186010 41530 186012
rect 41781 186010 41847 186013
rect 41524 186008 41847 186010
rect 41524 185952 41786 186008
rect 41842 185952 41847 186008
rect 41524 185950 41847 185952
rect 41524 185948 41530 185950
rect 41781 185947 41847 185950
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 666694 184378 666754 184386
rect 668025 184378 668091 184381
rect 666694 184376 668091 184378
rect 666694 184320 668030 184376
rect 668086 184320 668091 184376
rect 666694 184318 668091 184320
rect 41781 184108 41847 184109
rect 41781 184104 41828 184108
rect 41892 184106 41898 184108
rect 41781 184048 41786 184104
rect 41781 184044 41828 184048
rect 41892 184046 41938 184106
rect 41892 184044 41898 184046
rect 41781 184043 41847 184044
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 668025 184315 668091 184318
rect 589457 183562 589523 183565
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 589457 183499 589523 183502
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 42425 180706 42491 180709
rect 46933 180706 46999 180709
rect 42425 180704 46999 180706
rect 42425 180648 42430 180704
rect 42486 180648 46938 180704
rect 46994 180648 46999 180704
rect 42425 180646 46999 180648
rect 42425 180643 42491 180646
rect 46933 180643 46999 180646
rect 589641 180298 589707 180301
rect 672257 180298 672323 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 672257 180296 676322 180298
rect 672257 180240 672262 180296
rect 672318 180240 676322 180296
rect 672257 180238 676322 180240
rect 589641 180235 589707 180238
rect 672257 180235 672323 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 666356 179490 666754 179550
rect 666694 179482 666754 179490
rect 668025 179482 668091 179485
rect 666694 179480 668091 179482
rect 666694 179424 668030 179480
rect 668086 179424 668091 179480
rect 666694 179422 668091 179424
rect 668025 179419 668091 179422
rect 42057 179346 42123 179349
rect 50705 179346 50771 179349
rect 42057 179344 50771 179346
rect 42057 179288 42062 179344
rect 42118 179288 50710 179344
rect 50766 179288 50771 179344
rect 42057 179286 50771 179288
rect 42057 179283 42123 179286
rect 50705 179283 50771 179286
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 676262 178500 676322 180238
rect 674281 178122 674347 178125
rect 674281 178120 676292 178122
rect 674281 178064 674286 178120
rect 674342 178064 676292 178120
rect 674281 178062 676292 178064
rect 674281 178059 674347 178062
rect 671153 177986 671219 177989
rect 666694 177984 671219 177986
rect 666694 177928 671158 177984
rect 671214 177928 671219 177984
rect 666694 177926 671219 177928
rect 666694 177918 666754 177926
rect 671153 177923 671219 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 672901 177714 672967 177717
rect 672901 177712 676292 177714
rect 672901 177656 672906 177712
rect 672962 177656 676292 177712
rect 672901 177654 676292 177656
rect 672901 177651 672967 177654
rect 673913 177306 673979 177309
rect 673913 177304 676292 177306
rect 673913 177248 673918 177304
rect 673974 177248 676292 177304
rect 673913 177246 676292 177248
rect 673913 177243 673979 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 673361 176898 673427 176901
rect 673361 176896 676292 176898
rect 673361 176840 673366 176896
rect 673422 176840 676292 176896
rect 673361 176838 676292 176840
rect 673361 176835 673427 176838
rect 667013 176490 667079 176493
rect 667013 176488 676292 176490
rect 667013 176432 667018 176488
rect 667074 176432 676292 176488
rect 667013 176430 676292 176432
rect 667013 176427 667079 176430
rect 672349 176082 672415 176085
rect 672349 176080 676292 176082
rect 672349 176024 672354 176080
rect 672410 176024 676292 176080
rect 672349 176022 676292 176024
rect 672349 176019 672415 176022
rect 672533 175674 672599 175677
rect 672533 175672 676292 175674
rect 672533 175616 672538 175672
rect 672594 175616 676292 175672
rect 672533 175614 676292 175616
rect 672533 175611 672599 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 674649 175266 674715 175269
rect 674649 175264 676292 175266
rect 575982 175130 576042 175236
rect 674649 175208 674654 175264
rect 674710 175208 676292 175264
rect 674649 175206 676292 175208
rect 674649 175203 674715 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 667749 174994 667815 174997
rect 667749 174992 672826 174994
rect 667749 174936 667754 174992
rect 667810 174936 672826 174992
rect 667749 174934 672826 174936
rect 667749 174931 667815 174934
rect 672766 174858 672826 174934
rect 672766 174798 676292 174858
rect 669405 174722 669471 174725
rect 666694 174720 669471 174722
rect 666694 174664 669410 174720
rect 669466 174664 669471 174720
rect 666694 174662 669471 174664
rect 666694 174654 666754 174662
rect 669405 174659 669471 174662
rect 666356 174594 666754 174654
rect 674373 174450 674439 174453
rect 674373 174448 676292 174450
rect 674373 174392 674378 174448
rect 674434 174392 676292 174448
rect 674373 174390 676292 174392
rect 674373 174387 674439 174390
rect 675201 174042 675267 174045
rect 675201 174040 676292 174042
rect 675201 173984 675206 174040
rect 675262 173984 676292 174040
rect 675201 173982 676292 173984
rect 675201 173979 675267 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675518 173572 675524 173636
rect 675588 173634 675594 173636
rect 675588 173574 676292 173634
rect 675588 173572 675594 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 668209 173090 668275 173093
rect 666694 173088 668275 173090
rect 666694 173032 668214 173088
rect 668270 173032 668275 173088
rect 666694 173030 668275 173032
rect 666694 173022 666754 173030
rect 668209 173027 668275 173030
rect 666356 172962 666754 173022
rect 675886 172756 675892 172820
rect 675956 172818 675962 172820
rect 675956 172758 676292 172818
rect 675956 172756 675962 172758
rect 675702 172348 675708 172412
rect 675772 172410 675778 172412
rect 675772 172350 676292 172410
rect 675772 172348 675778 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 669405 172002 669471 172005
rect 669405 172000 676292 172002
rect 669405 171944 669410 172000
rect 669466 171944 676292 172000
rect 669405 171942 676292 171944
rect 669405 171939 669471 171942
rect 678237 171594 678303 171597
rect 678237 171592 678316 171594
rect 678237 171536 678242 171592
rect 678298 171536 678316 171592
rect 678237 171534 678316 171536
rect 678237 171531 678303 171534
rect 675385 171186 675451 171189
rect 675385 171184 676292 171186
rect 675385 171128 675390 171184
rect 675446 171128 676292 171184
rect 675385 171126 676292 171128
rect 675385 171123 675451 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 669446 170988 669452 171052
rect 669516 171050 669522 171052
rect 670601 171050 670667 171053
rect 669516 171048 670667 171050
rect 669516 170992 670606 171048
rect 670662 170992 670667 171048
rect 669516 170990 670667 170992
rect 669516 170988 669522 170990
rect 670601 170987 670667 170990
rect 671981 170778 672047 170781
rect 671981 170776 676292 170778
rect 671981 170720 671986 170776
rect 672042 170720 676292 170776
rect 671981 170718 676292 170720
rect 671981 170715 672047 170718
rect 589641 170506 589707 170509
rect 589641 170504 592572 170506
rect 589641 170448 589646 170504
rect 589702 170448 592572 170504
rect 589641 170446 592572 170448
rect 589641 170443 589707 170446
rect 670601 170370 670667 170373
rect 670601 170368 676292 170370
rect 670601 170312 670606 170368
rect 670662 170312 676292 170368
rect 670601 170310 676292 170312
rect 670601 170307 670667 170310
rect 676581 169962 676647 169965
rect 676581 169960 676660 169962
rect 676581 169904 676586 169960
rect 676642 169904 676660 169960
rect 676581 169902 676660 169904
rect 676581 169899 676647 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 675940 169698 676230 169758
rect 668393 169690 668459 169693
rect 675940 169692 676000 169698
rect 666694 169688 668459 169690
rect 666694 169632 668398 169688
rect 668454 169632 668459 169688
rect 666694 169630 668459 169632
rect 668393 169627 668459 169630
rect 675886 169628 675892 169692
rect 675956 169630 676000 169692
rect 675956 169628 675962 169630
rect 676170 169554 676230 169698
rect 676170 169494 676292 169554
rect 674833 169418 674899 169421
rect 675937 169418 676003 169421
rect 674833 169416 676003 169418
rect 674833 169360 674838 169416
rect 674894 169360 675942 169416
rect 675998 169360 676003 169416
rect 674833 169358 676003 169360
rect 674833 169355 674899 169358
rect 675937 169355 676003 169358
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 672165 169146 672231 169149
rect 672165 169144 676292 169146
rect 672165 169088 672170 169144
rect 672226 169088 676292 169144
rect 672165 169086 676292 169088
rect 672165 169083 672231 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673913 168738 673979 168741
rect 673913 168736 676292 168738
rect 673913 168680 673918 168736
rect 673974 168680 676292 168736
rect 673913 168678 676292 168680
rect 673913 168675 673979 168678
rect 672533 168330 672599 168333
rect 672533 168328 676292 168330
rect 672533 168272 672538 168328
rect 672594 168272 676292 168328
rect 672533 168270 676292 168272
rect 672533 168267 672599 168270
rect 666356 168066 666938 168126
rect 666878 167922 666938 168066
rect 673177 167922 673243 167925
rect 666878 167920 673243 167922
rect 666878 167864 673182 167920
rect 673238 167864 673243 167920
rect 666878 167862 673243 167864
rect 673177 167859 673243 167862
rect 675845 167922 675911 167925
rect 675845 167920 676292 167922
rect 675845 167864 675850 167920
rect 675906 167864 676292 167920
rect 675845 167862 676292 167864
rect 675845 167859 675911 167862
rect 675702 167452 675708 167516
rect 675772 167514 675778 167516
rect 675772 167454 676292 167514
rect 675772 167452 675778 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676029 167106 676095 167109
rect 676029 167104 676292 167106
rect 676029 167048 676034 167104
rect 676090 167048 676292 167104
rect 676029 167046 676292 167048
rect 676029 167043 676095 167046
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 673085 166970 673151 166973
rect 675845 166970 675911 166973
rect 673085 166968 675911 166970
rect 673085 166912 673090 166968
rect 673146 166912 675850 166968
rect 675906 166912 675911 166968
rect 673085 166910 675911 166912
rect 673085 166907 673151 166910
rect 675845 166907 675911 166910
rect 676814 166429 676874 166668
rect 676581 166428 676647 166429
rect 676581 166426 676628 166428
rect 676536 166424 676628 166426
rect 676536 166368 676586 166424
rect 676536 166366 676628 166368
rect 676581 166364 676628 166366
rect 676692 166364 676698 166428
rect 676814 166424 676923 166429
rect 676814 166368 676862 166424
rect 676918 166368 676923 166424
rect 676814 166366 676923 166368
rect 676581 166363 676647 166364
rect 676857 166363 676923 166366
rect 589457 165610 589523 165613
rect 672901 165610 672967 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 672901 165608 676095 165610
rect 672901 165552 672906 165608
rect 672962 165552 676034 165608
rect 676090 165552 676095 165608
rect 672901 165550 676095 165552
rect 589457 165547 589523 165550
rect 672901 165547 672967 165550
rect 676029 165547 676095 165550
rect 668209 164930 668275 164933
rect 666694 164928 668275 164930
rect 666694 164872 668214 164928
rect 668270 164872 668275 164928
rect 666694 164870 668275 164872
rect 666694 164862 666754 164870
rect 668209 164867 668275 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668209 163298 668275 163301
rect 666694 163296 668275 163298
rect 666694 163240 668214 163296
rect 668270 163240 668275 163296
rect 666694 163238 668275 163240
rect 666694 163230 666754 163238
rect 668209 163235 668275 163238
rect 666356 163170 666754 163230
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675518 162148 675524 162212
rect 675588 162210 675594 162212
rect 676070 162210 676076 162212
rect 675588 162150 676076 162210
rect 675588 162148 675594 162150
rect 676070 162148 676076 162150
rect 676140 162148 676146 162212
rect 673310 161332 673316 161396
rect 673380 161394 673386 161396
rect 675477 161394 675543 161397
rect 673380 161392 675543 161394
rect 673380 161336 675482 161392
rect 675538 161336 675543 161392
rect 673380 161334 675543 161336
rect 673380 161332 673386 161334
rect 675477 161331 675543 161334
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 674833 160578 674899 160581
rect 675477 160578 675543 160581
rect 674833 160576 675543 160578
rect 674833 160520 674838 160576
rect 674894 160520 675482 160576
rect 675538 160520 675543 160576
rect 674833 160518 675543 160520
rect 674833 160515 674899 160518
rect 675477 160515 675543 160518
rect 668209 160034 668275 160037
rect 666694 160032 668275 160034
rect 575982 159898 576042 160004
rect 666694 159976 668214 160032
rect 668270 159976 668275 160032
rect 666694 159974 668275 159976
rect 666694 159966 666754 159974
rect 668209 159971 668275 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 675017 159490 675083 159493
rect 675477 159490 675543 159493
rect 675017 159488 675543 159490
rect 675017 159432 675022 159488
rect 675078 159432 675482 159488
rect 675538 159432 675543 159488
rect 675017 159430 675543 159432
rect 675017 159427 675083 159430
rect 675477 159427 675543 159430
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 578417 158402 578483 158405
rect 668577 158402 668643 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 668643 158402
rect 666694 158344 668582 158400
rect 668638 158344 668643 158400
rect 666694 158342 668643 158344
rect 666694 158334 666754 158342
rect 668577 158339 668643 158342
rect 666356 158274 666754 158334
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 675753 157042 675819 157045
rect 676438 157042 676444 157044
rect 675753 157040 676444 157042
rect 675753 156984 675758 157040
rect 675814 156984 676444 157040
rect 675753 156982 676444 156984
rect 675753 156979 675819 156982
rect 676438 156980 676444 156982
rect 676508 156980 676514 157044
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 675753 155682 675819 155685
rect 676254 155682 676260 155684
rect 675753 155680 676260 155682
rect 675753 155624 675758 155680
rect 675814 155624 676260 155680
rect 675753 155622 676260 155624
rect 675753 155619 675819 155622
rect 676254 155620 676260 155622
rect 676324 155620 676330 155684
rect 668301 155138 668367 155141
rect 666694 155136 668367 155138
rect 666694 155080 668306 155136
rect 668362 155080 668367 155136
rect 666694 155078 668367 155080
rect 666694 155070 666754 155078
rect 668301 155075 668367 155078
rect 666356 155010 666754 155070
rect 671981 154458 672047 154461
rect 675109 154458 675175 154461
rect 671981 154456 675175 154458
rect 671981 154400 671986 154456
rect 672042 154400 675114 154456
rect 675170 154400 675175 154456
rect 671981 154398 675175 154400
rect 671981 154395 672047 154398
rect 675109 154395 675175 154398
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 154050 578391 154053
rect 575798 154048 578391 154050
rect 575798 153992 578330 154048
rect 578386 153992 578391 154048
rect 575798 153990 578391 153992
rect 575798 153476 575858 153990
rect 578325 153987 578391 153990
rect 666356 153378 666938 153438
rect 666878 153370 666938 153378
rect 673729 153370 673795 153373
rect 666878 153368 673795 153370
rect 666878 153312 673734 153368
rect 673790 153312 673795 153368
rect 666878 153310 673795 153312
rect 673729 153307 673795 153310
rect 672165 153098 672231 153101
rect 675109 153098 675175 153101
rect 672165 153096 675175 153098
rect 672165 153040 672170 153096
rect 672226 153040 675114 153096
rect 675170 153040 675175 153096
rect 672165 153038 675175 153040
rect 672165 153035 672231 153038
rect 675109 153035 675175 153038
rect 675661 153098 675727 153101
rect 675886 153098 675892 153100
rect 675661 153096 675892 153098
rect 675661 153040 675666 153096
rect 675722 153040 675892 153096
rect 675661 153038 675892 153040
rect 675661 153035 675727 153038
rect 675886 153036 675892 153038
rect 675956 153036 675962 153100
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 675753 151466 675819 151469
rect 676622 151466 676628 151468
rect 675753 151464 676628 151466
rect 675753 151408 675758 151464
rect 675814 151408 676628 151464
rect 675753 151406 676628 151408
rect 675753 151403 675819 151406
rect 676622 151404 676628 151406
rect 676692 151404 676698 151468
rect 673913 151058 673979 151061
rect 675109 151058 675175 151061
rect 673913 151056 675175 151058
rect 673913 151000 673918 151056
rect 673974 151000 675114 151056
rect 675170 151000 675175 151056
rect 673913 150998 675175 151000
rect 673913 150995 673979 150998
rect 675109 150995 675175 150998
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 671705 150242 671771 150245
rect 666694 150240 671771 150242
rect 666694 150184 671710 150240
rect 671766 150184 671771 150240
rect 666694 150182 671771 150184
rect 666694 150174 666754 150182
rect 671705 150179 671771 150182
rect 666356 150114 666754 150174
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 669405 149018 669471 149021
rect 675293 149018 675359 149021
rect 669405 149016 675359 149018
rect 669405 148960 669410 149016
rect 669466 148960 675298 149016
rect 675354 148960 675359 149016
rect 669405 148958 675359 148960
rect 669405 148955 669471 148958
rect 675293 148955 675359 148958
rect 668209 148610 668275 148613
rect 666694 148608 668275 148610
rect 666694 148552 668214 148608
rect 668270 148552 668275 148608
rect 666694 148550 668275 148552
rect 666694 148542 666754 148550
rect 668209 148547 668275 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 588537 147658 588603 147661
rect 670601 147658 670667 147661
rect 675109 147658 675175 147661
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 670601 147656 675175 147658
rect 670601 147600 670606 147656
rect 670662 147600 675114 147656
rect 675170 147600 675175 147656
rect 670601 147598 675175 147600
rect 588537 147595 588603 147598
rect 670601 147595 670667 147598
rect 675109 147595 675175 147598
rect 675661 147660 675727 147661
rect 675661 147656 675708 147660
rect 675772 147658 675778 147660
rect 675661 147600 675666 147656
rect 675661 147596 675708 147600
rect 675772 147598 675818 147658
rect 675772 147596 675778 147598
rect 675661 147595 675727 147596
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 671521 145346 671587 145349
rect 666694 145344 671587 145346
rect 666694 145288 671526 145344
rect 671582 145288 671587 145344
rect 666694 145286 671587 145288
rect 666694 145278 666754 145286
rect 671521 145283 671587 145286
rect 666356 145218 666754 145278
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 669221 143714 669287 143717
rect 666694 143712 669287 143714
rect 666694 143656 669226 143712
rect 669282 143656 669287 143712
rect 666694 143654 669287 143656
rect 666694 143646 666754 143654
rect 669221 143651 669287 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 669262 140450 669268 140452
rect 666694 140390 669268 140450
rect 666694 140382 666754 140390
rect 669262 140388 669268 140390
rect 669332 140388 669338 140452
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 668945 138818 669011 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 669011 138818
rect 666694 138760 668950 138816
rect 669006 138760 669011 138816
rect 666694 138758 669011 138760
rect 666694 138750 666754 138758
rect 668945 138755 669011 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 668209 135554 668275 135557
rect 666694 135552 668275 135554
rect 666694 135496 668214 135552
rect 668270 135496 668275 135552
rect 666694 135494 668275 135496
rect 666694 135486 666754 135494
rect 668209 135491 668275 135494
rect 666356 135426 666754 135486
rect 590377 134602 590443 134605
rect 667381 134602 667447 134605
rect 676029 134602 676095 134605
rect 590377 134600 592572 134602
rect 590377 134544 590382 134600
rect 590438 134544 592572 134600
rect 590377 134542 592572 134544
rect 667381 134600 676095 134602
rect 667381 134544 667386 134600
rect 667442 134544 676034 134600
rect 676090 134544 676095 134600
rect 667381 134542 676095 134544
rect 590377 134539 590443 134542
rect 667381 134539 667447 134542
rect 676029 134539 676095 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 669221 133786 669287 133789
rect 666694 133784 669287 133786
rect 666694 133728 669226 133784
rect 669282 133728 669287 133784
rect 666694 133726 669287 133728
rect 669221 133723 669287 133726
rect 667565 133378 667631 133381
rect 667565 133376 676292 133378
rect 667565 133320 667570 133376
rect 667626 133320 676292 133376
rect 667565 133318 676292 133320
rect 667565 133315 667631 133318
rect 589457 132970 589523 132973
rect 589457 132968 592572 132970
rect 589457 132912 589462 132968
rect 589518 132912 592572 132968
rect 589457 132910 592572 132912
rect 589457 132907 589523 132910
rect 674046 132908 674052 132972
rect 674116 132970 674122 132972
rect 674116 132910 676292 132970
rect 674116 132908 674122 132910
rect 669221 132698 669287 132701
rect 673494 132698 673500 132700
rect 669221 132696 673500 132698
rect 669221 132640 669226 132696
rect 669282 132640 673500 132696
rect 669221 132638 673500 132640
rect 669221 132635 669287 132638
rect 673494 132636 673500 132638
rect 673564 132636 673570 132700
rect 676029 132562 676095 132565
rect 676029 132560 676292 132562
rect 676029 132504 676034 132560
rect 676090 132504 676292 132560
rect 676029 132502 676292 132504
rect 676029 132499 676095 132502
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 673361 132154 673427 132157
rect 673361 132152 676292 132154
rect 673361 132096 673366 132152
rect 673422 132096 676292 132152
rect 673361 132094 676292 132096
rect 673361 132091 673427 132094
rect 672165 131746 672231 131749
rect 672165 131744 676292 131746
rect 672165 131688 672170 131744
rect 672226 131688 676292 131744
rect 672165 131686 676292 131688
rect 672165 131683 672231 131686
rect 672349 131474 672415 131477
rect 672349 131472 676322 131474
rect 672349 131416 672354 131472
rect 672410 131416 676322 131472
rect 672349 131414 676322 131416
rect 672349 131411 672415 131414
rect 589457 131338 589523 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 676262 131308 676322 131414
rect 589457 131278 592572 131280
rect 589457 131275 589523 131278
rect 668945 131202 669011 131205
rect 672533 131202 672599 131205
rect 668945 131200 672599 131202
rect 668945 131144 668950 131200
rect 669006 131144 672538 131200
rect 672594 131144 672599 131200
rect 668945 131142 672599 131144
rect 668945 131139 669011 131142
rect 672533 131139 672599 131142
rect 669957 130930 670023 130933
rect 669957 130928 676292 130930
rect 669957 130872 669962 130928
rect 670018 130872 676292 130928
rect 669957 130870 676292 130872
rect 669957 130867 670023 130870
rect 668761 130658 668827 130661
rect 666694 130656 668827 130658
rect 666694 130600 668766 130656
rect 668822 130600 668827 130656
rect 666694 130598 668827 130600
rect 666694 130590 666754 130598
rect 668761 130595 668827 130598
rect 666356 130530 666754 130590
rect 674649 130522 674715 130525
rect 674649 130520 676292 130522
rect 674649 130464 674654 130520
rect 674710 130464 676292 130520
rect 674649 130462 676292 130464
rect 674649 130459 674715 130462
rect 676213 130250 676279 130253
rect 676213 130248 676322 130250
rect 676213 130192 676218 130248
rect 676274 130192 676322 130248
rect 676213 130187 676322 130192
rect 676262 130084 676322 130187
rect 578877 129706 578943 129709
rect 575798 129704 578943 129706
rect 575798 129648 578882 129704
rect 578938 129648 578943 129704
rect 575798 129646 578943 129648
rect 575798 129540 575858 129646
rect 578877 129643 578943 129646
rect 588721 129706 588787 129709
rect 674373 129706 674439 129709
rect 588721 129704 592572 129706
rect 588721 129648 588726 129704
rect 588782 129648 592572 129704
rect 588721 129646 592572 129648
rect 674373 129704 676292 129706
rect 674373 129648 674378 129704
rect 674434 129648 676292 129704
rect 674373 129646 676292 129648
rect 588721 129643 588787 129646
rect 674373 129643 674439 129646
rect 674281 129298 674347 129301
rect 674281 129296 676292 129298
rect 674281 129240 674286 129296
rect 674342 129240 676292 129296
rect 674281 129238 676292 129240
rect 674281 129235 674347 129238
rect 668577 129026 668643 129029
rect 666694 129024 668643 129026
rect 666694 128968 668582 129024
rect 668638 128968 668643 129024
rect 666694 128966 668643 128968
rect 666694 128958 666754 128966
rect 668577 128963 668643 128966
rect 666356 128898 666754 128958
rect 675201 128890 675267 128893
rect 675201 128888 676292 128890
rect 675201 128832 675206 128888
rect 675262 128832 676292 128888
rect 675201 128830 676292 128832
rect 675201 128827 675267 128830
rect 676446 128210 676506 128452
rect 676673 128210 676739 128213
rect 676446 128208 676739 128210
rect 676446 128152 676678 128208
rect 676734 128152 676739 128208
rect 676446 128150 676739 128152
rect 676673 128147 676739 128150
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 579521 127938 579587 127941
rect 575798 127936 579587 127938
rect 575798 127880 579526 127936
rect 579582 127880 579587 127936
rect 575798 127878 579587 127880
rect 575798 127364 575858 127878
rect 579521 127875 579587 127878
rect 676446 127805 676506 128044
rect 668577 127802 668643 127805
rect 676213 127802 676279 127805
rect 668577 127800 676279 127802
rect 668577 127744 668582 127800
rect 668638 127744 676218 127800
rect 676274 127744 676279 127800
rect 668577 127742 676279 127744
rect 668577 127739 668643 127742
rect 676213 127739 676279 127742
rect 676397 127800 676506 127805
rect 676397 127744 676402 127800
rect 676458 127744 676506 127800
rect 676397 127742 676506 127744
rect 676397 127739 676463 127742
rect 676446 127396 676506 127636
rect 676438 127332 676444 127396
rect 676508 127332 676514 127396
rect 675886 127196 675892 127260
rect 675956 127258 675962 127260
rect 675956 127198 676292 127258
rect 675956 127196 675962 127198
rect 671981 126850 672047 126853
rect 671981 126848 676292 126850
rect 671981 126792 671986 126848
rect 672042 126792 676292 126848
rect 671981 126790 676292 126792
rect 671981 126787 672047 126790
rect 590101 126442 590167 126445
rect 590101 126440 592572 126442
rect 590101 126384 590106 126440
rect 590162 126384 592572 126440
rect 590101 126382 592572 126384
rect 590101 126379 590167 126382
rect 676070 126108 676076 126172
rect 676140 126170 676146 126172
rect 676673 126170 676739 126173
rect 676140 126168 676739 126170
rect 676140 126112 676678 126168
rect 676734 126112 676739 126168
rect 676140 126110 676739 126112
rect 682886 126170 682946 126412
rect 683113 126170 683179 126173
rect 682886 126168 683179 126170
rect 682886 126112 683118 126168
rect 683174 126112 683179 126168
rect 682886 126110 683179 126112
rect 676140 126108 676146 126110
rect 676673 126107 676739 126110
rect 683113 126107 683179 126110
rect 669221 126034 669287 126037
rect 672717 126034 672783 126037
rect 669221 126032 672783 126034
rect 669221 125976 669226 126032
rect 669282 125976 672722 126032
rect 672778 125976 672783 126032
rect 669221 125974 672783 125976
rect 669221 125971 669287 125974
rect 672717 125971 672783 125974
rect 676814 125765 676874 126004
rect 670734 125762 670740 125764
rect 666694 125702 670740 125762
rect 666694 125694 666754 125702
rect 670734 125700 670740 125702
rect 670804 125700 670810 125764
rect 676814 125760 676923 125765
rect 676814 125704 676862 125760
rect 676918 125704 676923 125760
rect 676814 125702 676923 125704
rect 676857 125699 676923 125702
rect 666356 125634 666754 125694
rect 674465 125626 674531 125629
rect 674465 125624 676292 125626
rect 674465 125568 674470 125624
rect 674526 125568 676292 125624
rect 674465 125566 676292 125568
rect 674465 125563 674531 125566
rect 578325 125354 578391 125357
rect 575798 125352 578391 125354
rect 575798 125296 578330 125352
rect 578386 125296 578391 125352
rect 575798 125294 578391 125296
rect 575798 125188 575858 125294
rect 578325 125291 578391 125294
rect 668025 125354 668091 125357
rect 675937 125354 676003 125357
rect 668025 125352 676003 125354
rect 668025 125296 668030 125352
rect 668086 125296 675942 125352
rect 675998 125296 676003 125352
rect 668025 125294 676003 125296
rect 668025 125291 668091 125294
rect 675937 125291 676003 125294
rect 676121 125354 676187 125357
rect 676581 125354 676647 125357
rect 678973 125354 679039 125357
rect 676121 125352 676230 125354
rect 676121 125296 676126 125352
rect 676182 125296 676230 125352
rect 676121 125291 676230 125296
rect 676581 125352 679039 125354
rect 676581 125296 676586 125352
rect 676642 125296 678978 125352
rect 679034 125296 679039 125352
rect 676581 125294 679039 125296
rect 676581 125291 676647 125294
rect 678973 125291 679039 125294
rect 676170 125218 676230 125291
rect 676170 125158 676292 125218
rect 590561 124810 590627 124813
rect 674649 124810 674715 124813
rect 590561 124808 592572 124810
rect 590561 124752 590566 124808
rect 590622 124752 592572 124808
rect 590561 124750 592572 124752
rect 674649 124808 676292 124810
rect 674649 124752 674654 124808
rect 674710 124752 676292 124808
rect 674649 124750 676292 124752
rect 590561 124747 590627 124750
rect 674649 124747 674715 124750
rect 676254 124476 676260 124540
rect 676324 124476 676330 124540
rect 676262 124372 676322 124476
rect 669221 124130 669287 124133
rect 666694 124128 669287 124130
rect 666694 124072 669226 124128
rect 669282 124072 669287 124128
rect 666694 124070 669287 124072
rect 666694 124062 666754 124070
rect 669221 124067 669287 124070
rect 666356 124002 666754 124062
rect 672717 123994 672783 123997
rect 672717 123992 676292 123994
rect 672717 123936 672722 123992
rect 672778 123936 676292 123992
rect 672717 123934 676292 123936
rect 672717 123931 672783 123934
rect 578693 123586 578759 123589
rect 575798 123584 578759 123586
rect 575798 123528 578698 123584
rect 578754 123528 578759 123584
rect 575798 123526 578759 123528
rect 575798 123012 575858 123526
rect 578693 123523 578759 123526
rect 673729 123586 673795 123589
rect 673729 123584 676292 123586
rect 673729 123528 673734 123584
rect 673790 123528 676292 123584
rect 673729 123526 676292 123528
rect 673729 123523 673795 123526
rect 589457 123178 589523 123181
rect 673545 123178 673611 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 673545 123176 676292 123178
rect 673545 123120 673550 123176
rect 673606 123120 676292 123176
rect 673545 123118 676292 123120
rect 589457 123115 589523 123118
rect 673545 123115 673611 123118
rect 676806 122844 676812 122908
rect 676876 122906 676882 122908
rect 683113 122906 683179 122909
rect 676876 122904 683179 122906
rect 676876 122848 683118 122904
rect 683174 122848 683179 122904
rect 676876 122846 683179 122848
rect 676876 122844 676882 122846
rect 683113 122843 683179 122846
rect 671521 122770 671587 122773
rect 671521 122768 676292 122770
rect 671521 122712 671526 122768
rect 671582 122712 676292 122768
rect 671521 122710 676292 122712
rect 671521 122707 671587 122710
rect 677550 122093 677610 122332
rect 677550 122088 677659 122093
rect 677550 122032 677598 122088
rect 677654 122032 677659 122088
rect 677550 122030 677659 122032
rect 677593 122027 677659 122030
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 678973 121682 679039 121685
rect 678973 121680 679082 121682
rect 678973 121624 678978 121680
rect 679034 121624 679082 121680
rect 589273 121546 589339 121549
rect 589273 121544 592572 121546
rect 589273 121488 589278 121544
rect 589334 121488 592572 121544
rect 589273 121486 592572 121488
rect 589273 121483 589339 121486
rect 578877 121410 578943 121413
rect 575798 121408 578943 121410
rect 575798 121352 578882 121408
rect 578938 121352 578943 121408
rect 575798 121350 578943 121352
rect 575798 120836 575858 121350
rect 578877 121347 578943 121350
rect 670693 121410 670759 121413
rect 675894 121410 675954 121622
rect 678973 121619 679082 121624
rect 679022 121516 679082 121619
rect 670693 121408 675954 121410
rect 670693 121352 670698 121408
rect 670754 121352 675954 121408
rect 670693 121350 675954 121352
rect 670693 121347 670759 121350
rect 666356 120738 666938 120798
rect 666878 120458 666938 120738
rect 673361 120730 673427 120733
rect 676121 120730 676187 120733
rect 673361 120728 676187 120730
rect 673361 120672 673366 120728
rect 673422 120672 676126 120728
rect 676182 120672 676187 120728
rect 673361 120670 676187 120672
rect 673361 120667 673427 120670
rect 676121 120667 676187 120670
rect 674097 120458 674163 120461
rect 666878 120456 674163 120458
rect 666878 120400 674102 120456
rect 674158 120400 674163 120456
rect 666878 120398 674163 120400
rect 674097 120395 674163 120398
rect 668761 120050 668827 120053
rect 674281 120050 674347 120053
rect 668761 120048 674347 120050
rect 668761 119992 668766 120048
rect 668822 119992 674286 120048
rect 674342 119992 674347 120048
rect 668761 119990 674347 119992
rect 668761 119987 668827 119990
rect 674281 119987 674347 119990
rect 589641 119914 589707 119917
rect 589641 119912 592572 119914
rect 589641 119856 589646 119912
rect 589702 119856 592572 119912
rect 589641 119854 592572 119856
rect 589641 119851 589707 119854
rect 668945 119234 669011 119237
rect 666694 119232 669011 119234
rect 666694 119176 668950 119232
rect 669006 119176 669011 119232
rect 666694 119174 669011 119176
rect 666694 119166 666754 119174
rect 668945 119171 669011 119174
rect 666356 119106 666754 119166
rect 575982 118418 576042 118660
rect 675293 118554 675359 118557
rect 675845 118554 675911 118557
rect 675293 118552 675911 118554
rect 675293 118496 675298 118552
rect 675354 118496 675850 118552
rect 675906 118496 675911 118552
rect 675293 118494 675911 118496
rect 675293 118491 675359 118494
rect 675845 118491 675911 118494
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 590101 118282 590167 118285
rect 590101 118280 592572 118282
rect 590101 118224 590106 118280
rect 590162 118224 592572 118280
rect 590101 118222 592572 118224
rect 590101 118219 590167 118222
rect 673085 117602 673151 117605
rect 666694 117600 673151 117602
rect 666694 117544 673090 117600
rect 673146 117544 673151 117600
rect 666694 117542 673151 117544
rect 666694 117534 666754 117542
rect 673085 117539 673151 117542
rect 666356 117474 666754 117534
rect 669221 117058 669287 117061
rect 673545 117058 673611 117061
rect 669221 117056 673611 117058
rect 669221 117000 669226 117056
rect 669282 117000 673550 117056
rect 673606 117000 673611 117056
rect 669221 116998 673611 117000
rect 669221 116995 669287 116998
rect 673545 116995 673611 116998
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 675017 116378 675083 116381
rect 675845 116378 675911 116381
rect 675017 116376 675911 116378
rect 675017 116320 675022 116376
rect 675078 116320 675850 116376
rect 675906 116320 675911 116376
rect 675017 116318 675911 116320
rect 675017 116315 675083 116318
rect 675845 116315 675911 116318
rect 667197 116106 667263 116109
rect 675477 116106 675543 116109
rect 667197 116104 675543 116106
rect 667197 116048 667202 116104
rect 667258 116048 675482 116104
rect 675538 116048 675543 116104
rect 667197 116046 675543 116048
rect 667197 116043 667263 116046
rect 675477 116043 675543 116046
rect 675702 116044 675708 116108
rect 675772 116106 675778 116108
rect 677593 116106 677659 116109
rect 675772 116104 677659 116106
rect 675772 116048 677598 116104
rect 677654 116048 677659 116104
rect 675772 116046 677659 116048
rect 675772 116044 675778 116046
rect 677593 116043 677659 116046
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 672901 115834 672967 115837
rect 666694 115832 672967 115834
rect 666694 115776 672906 115832
rect 672962 115776 672967 115832
rect 666694 115774 672967 115776
rect 672901 115771 672967 115774
rect 590285 115018 590351 115021
rect 590285 115016 592572 115018
rect 590285 114960 590290 115016
rect 590346 114960 592572 115016
rect 590285 114958 592572 114960
rect 590285 114955 590351 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 669221 114338 669287 114341
rect 666694 114336 669287 114338
rect 666694 114280 669226 114336
rect 669282 114280 669287 114336
rect 666694 114278 669287 114280
rect 666694 114270 666754 114278
rect 669221 114275 669287 114278
rect 674833 114338 674899 114341
rect 675385 114338 675451 114341
rect 674833 114336 675451 114338
rect 674833 114280 674838 114336
rect 674894 114280 675390 114336
rect 675446 114280 675451 114336
rect 674833 114278 675451 114280
rect 674833 114275 674899 114278
rect 675385 114275 675451 114278
rect 675753 114338 675819 114341
rect 676806 114338 676812 114340
rect 675753 114336 676812 114338
rect 675753 114280 675758 114336
rect 675814 114280 676812 114336
rect 675753 114278 676812 114280
rect 675753 114275 675819 114278
rect 676806 114276 676812 114278
rect 676876 114276 676882 114340
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 671521 112706 671587 112709
rect 666694 112704 671587 112706
rect 666694 112648 671526 112704
rect 671582 112648 671587 112704
rect 666694 112646 671587 112648
rect 666694 112638 666754 112646
rect 671521 112643 671587 112646
rect 666356 112578 666754 112638
rect 579521 112570 579587 112573
rect 575798 112568 579587 112570
rect 575798 112512 579526 112568
rect 579582 112512 579587 112568
rect 575798 112510 579587 112512
rect 575798 112132 575858 112510
rect 579521 112507 579587 112510
rect 675753 112434 675819 112437
rect 676438 112434 676444 112436
rect 675753 112432 676444 112434
rect 675753 112376 675758 112432
rect 675814 112376 676444 112432
rect 675753 112374 676444 112376
rect 675753 112371 675819 112374
rect 676438 112372 676444 112374
rect 676508 112372 676514 112436
rect 589457 111754 589523 111757
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 589457 111691 589523 111694
rect 674465 111346 674531 111349
rect 675385 111346 675451 111349
rect 674465 111344 675451 111346
rect 674465 111288 674470 111344
rect 674526 111288 675390 111344
rect 675446 111288 675451 111344
rect 674465 111286 675451 111288
rect 674465 111283 674531 111286
rect 675385 111283 675451 111286
rect 668209 111074 668275 111077
rect 666694 111072 668275 111074
rect 666694 111016 668214 111072
rect 668270 111016 668275 111072
rect 666694 111014 668275 111016
rect 666694 111006 666754 111014
rect 668209 111011 668275 111014
rect 666356 110946 666754 111006
rect 675753 110394 675819 110397
rect 676254 110394 676260 110396
rect 675753 110392 676260 110394
rect 675753 110336 675758 110392
rect 675814 110336 676260 110392
rect 675753 110334 676260 110336
rect 675753 110331 675819 110334
rect 676254 110332 676260 110334
rect 676324 110332 676330 110396
rect 579337 110122 579403 110125
rect 575798 110120 579403 110122
rect 575798 110064 579342 110120
rect 579398 110064 579403 110120
rect 575798 110062 579403 110064
rect 575798 109956 575858 110062
rect 579337 110059 579403 110062
rect 589457 110122 589523 110125
rect 589457 110120 592572 110122
rect 589457 110064 589462 110120
rect 589518 110064 592572 110120
rect 589457 110062 592572 110064
rect 589457 110059 589523 110062
rect 666645 109374 666711 109377
rect 666356 109372 666711 109374
rect 666356 109316 666650 109372
rect 666706 109316 666711 109372
rect 666356 109314 666711 109316
rect 666645 109311 666711 109314
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 667933 107810 667999 107813
rect 666694 107808 667999 107810
rect 666694 107752 667938 107808
rect 667994 107752 667999 107808
rect 666694 107750 667999 107752
rect 666694 107742 666754 107750
rect 667933 107747 667999 107750
rect 666356 107682 666754 107742
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 672717 106586 672783 106589
rect 675109 106586 675175 106589
rect 672717 106584 675175 106586
rect 672717 106528 672722 106584
rect 672778 106528 675114 106584
rect 675170 106528 675175 106584
rect 672717 106526 675175 106528
rect 672717 106523 672783 106526
rect 675109 106523 675175 106526
rect 668117 106178 668183 106181
rect 672349 106178 672415 106181
rect 666694 106176 672415 106178
rect 666694 106120 668122 106176
rect 668178 106120 672354 106176
rect 672410 106120 672415 106176
rect 666694 106118 672415 106120
rect 666694 106110 666754 106118
rect 668117 106115 668183 106118
rect 672349 106115 672415 106118
rect 666356 106050 666754 106110
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 589825 105226 589891 105229
rect 589825 105224 592572 105226
rect 589825 105168 589830 105224
rect 589886 105168 592572 105224
rect 589825 105166 592572 105168
rect 589825 105163 589891 105166
rect 668301 104818 668367 104821
rect 668761 104818 668827 104821
rect 668301 104816 668827 104818
rect 668301 104760 668306 104816
rect 668362 104760 668766 104816
rect 668822 104760 668827 104816
rect 668301 104758 668827 104760
rect 668301 104755 668367 104758
rect 668761 104755 668827 104758
rect 673361 104546 673427 104549
rect 675109 104546 675175 104549
rect 673361 104544 675175 104546
rect 673361 104488 673366 104544
rect 673422 104488 675114 104544
rect 675170 104488 675175 104544
rect 673361 104486 675175 104488
rect 673361 104483 673427 104486
rect 675109 104483 675175 104486
rect 666356 104418 666754 104478
rect 666694 104410 666754 104418
rect 668301 104410 668367 104413
rect 666694 104408 668367 104410
rect 666694 104352 668306 104408
rect 668362 104352 668367 104408
rect 666694 104350 668367 104352
rect 668301 104347 668367 104350
rect 588537 103594 588603 103597
rect 588537 103592 592572 103594
rect 588537 103536 588542 103592
rect 588598 103536 592572 103592
rect 588537 103534 592572 103536
rect 588537 103531 588603 103534
rect 575982 103186 576042 103428
rect 578509 103186 578575 103189
rect 575982 103184 578575 103186
rect 575982 103128 578514 103184
rect 578570 103128 578575 103184
rect 575982 103126 578575 103128
rect 578509 103123 578575 103126
rect 675753 103186 675819 103189
rect 676070 103186 676076 103188
rect 675753 103184 676076 103186
rect 675753 103128 675758 103184
rect 675814 103128 676076 103184
rect 675753 103126 676076 103128
rect 675753 103123 675819 103126
rect 676070 103124 676076 103126
rect 676140 103124 676146 103188
rect 666356 102786 666754 102846
rect 666694 102778 666754 102786
rect 667933 102778 667999 102781
rect 668577 102778 668643 102781
rect 666694 102776 668643 102778
rect 666694 102720 667938 102776
rect 667994 102720 668582 102776
rect 668638 102720 668643 102776
rect 666694 102718 668643 102720
rect 667933 102715 667999 102718
rect 668577 102715 668643 102718
rect 675661 102644 675727 102645
rect 675661 102640 675708 102644
rect 675772 102642 675778 102644
rect 675661 102584 675666 102640
rect 675661 102580 675708 102584
rect 675772 102582 675818 102642
rect 675772 102580 675778 102582
rect 675661 102579 675727 102580
rect 589457 101962 589523 101965
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 589457 101899 589523 101902
rect 579153 101690 579219 101693
rect 575798 101688 579219 101690
rect 575798 101632 579158 101688
rect 579214 101632 579219 101688
rect 575798 101630 579219 101632
rect 575798 101252 575858 101630
rect 579153 101627 579219 101630
rect 671981 99378 672047 99381
rect 675293 99378 675359 99381
rect 671981 99376 675359 99378
rect 671981 99320 671986 99376
rect 672042 99320 675298 99376
rect 675354 99320 675359 99376
rect 671981 99318 675359 99320
rect 671981 99315 672047 99318
rect 675293 99315 675359 99318
rect 579521 99242 579587 99245
rect 575798 99240 579587 99242
rect 575798 99184 579526 99240
rect 579582 99184 579587 99240
rect 575798 99182 579587 99184
rect 575798 99076 575858 99182
rect 579521 99179 579587 99182
rect 578601 97474 578667 97477
rect 575798 97472 578667 97474
rect 575798 97416 578606 97472
rect 578662 97416 578667 97472
rect 575798 97414 578667 97416
rect 575798 96900 575858 97414
rect 578601 97411 578667 97414
rect 635549 96930 635615 96933
rect 635774 96930 635780 96932
rect 635549 96928 635780 96930
rect 635549 96872 635554 96928
rect 635610 96872 635780 96928
rect 635549 96870 635780 96872
rect 635549 96867 635615 96870
rect 635774 96868 635780 96870
rect 635844 96868 635850 96932
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 641989 96522 642055 96525
rect 647182 96522 647188 96524
rect 641989 96520 647188 96522
rect 641989 96464 641994 96520
rect 642050 96464 647188 96520
rect 641989 96462 647188 96464
rect 641989 96459 642055 96462
rect 647182 96460 647188 96462
rect 647252 96460 647258 96524
rect 645577 96114 645643 96117
rect 647509 96114 647575 96117
rect 645577 96112 647575 96114
rect 645577 96056 645582 96112
rect 645638 96056 647514 96112
rect 647570 96056 647575 96112
rect 645577 96054 647575 96056
rect 645577 96051 645643 96054
rect 647509 96051 647575 96054
rect 633934 95916 633940 95980
rect 634004 95978 634010 95980
rect 635733 95978 635799 95981
rect 634004 95976 635799 95978
rect 634004 95920 635738 95976
rect 635794 95920 635799 95976
rect 634004 95918 635799 95920
rect 634004 95916 634010 95918
rect 635733 95915 635799 95918
rect 645761 95570 645827 95573
rect 647509 95570 647575 95573
rect 645761 95568 647575 95570
rect 645761 95512 645766 95568
rect 645822 95512 647514 95568
rect 647570 95512 647575 95568
rect 645761 95510 647575 95512
rect 645761 95507 645827 95510
rect 647509 95507 647575 95510
rect 578325 95026 578391 95029
rect 575798 95024 578391 95026
rect 575798 94968 578330 95024
rect 578386 94968 578391 95024
rect 575798 94966 578391 94968
rect 575798 94724 575858 94966
rect 578325 94963 578391 94966
rect 647325 95026 647391 95029
rect 647325 95024 647434 95026
rect 647325 94968 647330 95024
rect 647386 94968 647434 95024
rect 647325 94963 647434 94968
rect 625429 94482 625495 94485
rect 625429 94480 628268 94482
rect 625429 94424 625434 94480
rect 625490 94424 628268 94480
rect 647374 94452 647434 94963
rect 625429 94422 628268 94424
rect 625429 94419 625495 94422
rect 654317 94210 654383 94213
rect 654317 94208 656788 94210
rect 654317 94152 654322 94208
rect 654378 94152 656788 94208
rect 654317 94150 656788 94152
rect 654317 94147 654383 94150
rect 626349 93666 626415 93669
rect 626349 93664 628268 93666
rect 626349 93608 626354 93664
rect 626410 93608 628268 93664
rect 626349 93606 628268 93608
rect 626349 93603 626415 93606
rect 654685 93394 654751 93397
rect 665357 93394 665423 93397
rect 654685 93392 656788 93394
rect 654685 93336 654690 93392
rect 654746 93336 656788 93392
rect 654685 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 654685 93331 654751 93334
rect 665357 93331 665423 93334
rect 579245 93122 579311 93125
rect 575798 93120 579311 93122
rect 575798 93064 579250 93120
rect 579306 93064 579311 93120
rect 575798 93062 579311 93064
rect 575798 92548 575858 93062
rect 579245 93059 579311 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 663793 93122 663859 93125
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626165 92850 626231 92853
rect 626165 92848 628268 92850
rect 626165 92792 626170 92848
rect 626226 92792 628268 92848
rect 626165 92790 628268 92792
rect 626165 92787 626231 92790
rect 656758 92548 656818 93062
rect 663566 93120 663859 93122
rect 663566 93064 663798 93120
rect 663854 93064 663859 93120
rect 663566 93062 663859 93064
rect 663566 92548 663626 93062
rect 663793 93059 663859 93062
rect 625797 92034 625863 92037
rect 648797 92034 648863 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 625797 91974 628268 91976
rect 648140 92032 648863 92034
rect 648140 91976 648802 92032
rect 648858 91976 648863 92032
rect 648140 91974 648863 91976
rect 625797 91971 625863 91974
rect 648797 91971 648863 91974
rect 663977 91762 664043 91765
rect 663596 91760 664043 91762
rect 663596 91704 663982 91760
rect 664038 91704 664043 91760
rect 663596 91702 664043 91704
rect 663977 91699 664043 91702
rect 655421 91490 655487 91493
rect 655421 91488 656788 91490
rect 655421 91432 655426 91488
rect 655482 91432 656788 91488
rect 655421 91430 656788 91432
rect 655421 91427 655487 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 578601 90946 578667 90949
rect 575798 90944 578667 90946
rect 575798 90888 578606 90944
rect 578662 90888 578667 90944
rect 575798 90886 578667 90888
rect 575798 90372 575858 90886
rect 578601 90883 578667 90886
rect 655421 90674 655487 90677
rect 664345 90674 664411 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 655421 90614 656788 90616
rect 663596 90672 664411 90674
rect 663596 90616 664350 90672
rect 664406 90616 664411 90672
rect 663596 90614 664411 90616
rect 655421 90611 655487 90614
rect 664345 90611 664411 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 647693 89858 647759 89861
rect 655789 89858 655855 89861
rect 664529 89858 664595 89861
rect 647693 89856 648170 89858
rect 647693 89800 647698 89856
rect 647754 89800 648170 89856
rect 647693 89798 648170 89800
rect 647693 89795 647759 89798
rect 626257 89586 626323 89589
rect 626257 89584 628268 89586
rect 626257 89528 626262 89584
rect 626318 89528 628268 89584
rect 648110 89556 648170 89798
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664595 89858
rect 663596 89800 664534 89856
rect 664590 89800 664595 89856
rect 663596 89798 664595 89800
rect 655789 89795 655855 89798
rect 664529 89795 664595 89798
rect 626257 89526 628268 89528
rect 626257 89523 626323 89526
rect 665173 89042 665239 89045
rect 663596 89040 665239 89042
rect 663596 88984 665178 89040
rect 665234 88984 665239 89040
rect 663596 88982 665239 88984
rect 665173 88979 665239 88982
rect 626441 88770 626507 88773
rect 626441 88768 628268 88770
rect 626441 88712 626446 88768
rect 626502 88712 628268 88768
rect 626441 88710 628268 88712
rect 626441 88707 626507 88710
rect 624969 88362 625035 88365
rect 626257 88362 626323 88365
rect 624969 88360 626323 88362
rect 624969 88304 624974 88360
rect 625030 88304 626262 88360
rect 626318 88304 626323 88360
rect 624969 88302 626323 88304
rect 624969 88299 625035 88302
rect 626257 88299 626323 88302
rect 575982 88090 576042 88196
rect 579245 88090 579311 88093
rect 575982 88088 579311 88090
rect 575982 88032 579250 88088
rect 579306 88032 579311 88088
rect 575982 88030 579311 88032
rect 579245 88027 579311 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 626257 87138 626323 87141
rect 650545 87138 650611 87141
rect 626257 87136 628268 87138
rect 626257 87080 626262 87136
rect 626318 87080 628268 87136
rect 626257 87078 628268 87080
rect 648140 87136 650611 87138
rect 648140 87080 650550 87136
rect 650606 87080 650611 87136
rect 648140 87078 650611 87080
rect 626257 87075 626323 87078
rect 650545 87075 650611 87078
rect 578325 86458 578391 86461
rect 575798 86456 578391 86458
rect 575798 86400 578330 86456
rect 578386 86400 578391 86456
rect 575798 86398 578391 86400
rect 575798 86020 575858 86398
rect 578325 86395 578391 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 626441 85506 626507 85509
rect 626441 85504 628268 85506
rect 626441 85448 626446 85504
rect 626502 85448 628268 85504
rect 626441 85446 628268 85448
rect 626441 85443 626507 85446
rect 625245 84690 625311 84693
rect 648613 84690 648679 84693
rect 625245 84688 628268 84690
rect 625245 84632 625250 84688
rect 625306 84632 628268 84688
rect 625245 84630 628268 84632
rect 648140 84688 648679 84690
rect 648140 84632 648618 84688
rect 648674 84632 648679 84688
rect 648140 84630 648679 84632
rect 625245 84627 625311 84630
rect 648613 84627 648679 84630
rect 579245 84010 579311 84013
rect 575798 84008 579311 84010
rect 575798 83952 579250 84008
rect 579306 83952 579311 84008
rect 575798 83950 579311 83952
rect 575798 83844 575858 83950
rect 579245 83947 579311 83950
rect 626441 83874 626507 83877
rect 626441 83872 628268 83874
rect 626441 83816 626446 83872
rect 626502 83816 628268 83872
rect 626441 83814 628268 83816
rect 626441 83811 626507 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 578877 82242 578943 82245
rect 650269 82242 650335 82245
rect 575798 82240 578943 82242
rect 575798 82184 578882 82240
rect 578938 82184 578943 82240
rect 648140 82240 650335 82242
rect 575798 82182 578943 82184
rect 575798 81668 575858 82182
rect 578877 82179 578943 82182
rect 628790 81698 628850 82212
rect 648140 82184 650274 82240
rect 650330 82184 650335 82240
rect 648140 82182 650335 82184
rect 650269 82179 650335 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 579429 80066 579495 80069
rect 575798 80064 579495 80066
rect 575798 80008 579434 80064
rect 579490 80008 579495 80064
rect 575798 80006 579495 80008
rect 575798 79492 575858 80006
rect 579429 80003 579495 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 635774 78100 635780 78164
rect 635844 78162 635850 78164
rect 647509 78162 647575 78165
rect 635844 78160 647575 78162
rect 635844 78104 647514 78160
rect 647570 78104 647575 78160
rect 635844 78102 647575 78104
rect 635844 78100 635850 78102
rect 647509 78099 647575 78102
rect 578233 77890 578299 77893
rect 575798 77888 578299 77890
rect 575798 77832 578238 77888
rect 578294 77832 578299 77888
rect 575798 77830 578299 77832
rect 575798 77316 575858 77830
rect 578233 77827 578299 77830
rect 580441 77890 580507 77893
rect 580441 77888 625170 77890
rect 580441 77832 580446 77888
rect 580502 77832 625170 77888
rect 580441 77830 625170 77832
rect 580441 77827 580507 77830
rect 625110 77618 625170 77830
rect 637062 77618 637068 77620
rect 625110 77558 637068 77618
rect 637062 77556 637068 77558
rect 637132 77618 637138 77620
rect 639597 77618 639663 77621
rect 637132 77616 639663 77618
rect 637132 77560 639602 77616
rect 639658 77560 639663 77616
rect 637132 77558 639663 77560
rect 637132 77556 637138 77558
rect 639597 77555 639663 77558
rect 623037 77346 623103 77349
rect 633893 77346 633959 77349
rect 623037 77344 633959 77346
rect 623037 77288 623042 77344
rect 623098 77288 633898 77344
rect 633954 77288 633959 77344
rect 623037 77286 633959 77288
rect 623037 77283 623103 77286
rect 633893 77283 633959 77286
rect 579245 75714 579311 75717
rect 575798 75712 579311 75714
rect 575798 75656 579250 75712
rect 579306 75656 579311 75712
rect 575798 75654 579311 75656
rect 575798 75140 575858 75654
rect 579245 75651 579311 75654
rect 646497 74218 646563 74221
rect 646454 74216 646563 74218
rect 646454 74160 646502 74216
rect 646558 74160 646563 74216
rect 646454 74155 646563 74160
rect 646454 73848 646514 74155
rect 579521 73130 579587 73133
rect 575798 73128 579587 73130
rect 575798 73072 579526 73128
rect 579582 73072 579587 73128
rect 575798 73070 579587 73072
rect 575798 72964 575858 73070
rect 579521 73067 579587 73070
rect 646681 71770 646747 71773
rect 646638 71768 646747 71770
rect 646638 71712 646686 71768
rect 646742 71712 646747 71768
rect 646638 71707 646747 71712
rect 646638 71400 646698 71707
rect 578509 71226 578575 71229
rect 575798 71224 578575 71226
rect 575798 71168 578514 71224
rect 578570 71168 578575 71224
rect 575798 71166 578575 71168
rect 575798 70788 575858 71166
rect 578509 71163 578575 71166
rect 646313 69186 646379 69189
rect 646270 69184 646379 69186
rect 646270 69128 646318 69184
rect 646374 69128 646379 69184
rect 646270 69123 646379 69128
rect 646270 68952 646330 69123
rect 575798 66874 575858 68612
rect 646129 67146 646195 67149
rect 646086 67144 646195 67146
rect 646086 67088 646134 67144
rect 646190 67088 646195 67144
rect 646086 67083 646195 67088
rect 579521 66874 579587 66877
rect 575798 66872 579587 66874
rect 575798 66816 579526 66872
rect 579582 66816 579587 66872
rect 575798 66814 579587 66816
rect 575798 66436 575858 66814
rect 579521 66811 579587 66814
rect 646086 66504 646146 67083
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 647325 64426 647391 64429
rect 646638 64424 647391 64426
rect 646638 64368 647330 64424
rect 647386 64368 647391 64424
rect 646638 64366 647391 64368
rect 646638 64056 646698 64366
rect 647325 64363 647391 64366
rect 648981 62114 649047 62117
rect 646638 62112 649047 62114
rect 575982 61842 576042 62084
rect 646638 62056 648986 62112
rect 649042 62056 649047 62112
rect 646638 62054 649047 62056
rect 579521 61842 579587 61845
rect 575982 61840 579587 61842
rect 575982 61784 579526 61840
rect 579582 61784 579587 61840
rect 575982 61782 579587 61784
rect 579521 61779 579587 61782
rect 646638 61608 646698 62054
rect 648981 62051 649047 62054
rect 578877 60482 578943 60485
rect 575798 60480 578943 60482
rect 575798 60424 578882 60480
rect 578938 60424 578943 60480
rect 575798 60422 578943 60424
rect 575798 59908 575858 60422
rect 578877 60419 578943 60422
rect 648613 59258 648679 59261
rect 646638 59256 648679 59258
rect 646638 59200 648618 59256
rect 648674 59200 648679 59256
rect 646638 59198 648679 59200
rect 646638 59160 646698 59198
rect 648613 59195 648679 59198
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 647509 57354 647575 57357
rect 646638 57352 647575 57354
rect 646638 57296 647514 57352
rect 647570 57296 647575 57352
rect 646638 57294 647575 57296
rect 646638 56712 646698 57294
rect 647509 57291 647575 57294
rect 578325 56130 578391 56133
rect 575798 56128 578391 56130
rect 575798 56072 578330 56128
rect 578386 56072 578391 56128
rect 575798 56070 578391 56072
rect 575798 55556 575858 56070
rect 578325 56067 578391 56070
rect 461710 54980 461716 55044
rect 461780 55042 461786 55044
rect 576117 55042 576183 55045
rect 461780 55040 576183 55042
rect 461780 54984 576122 55040
rect 576178 54984 576183 55040
rect 461780 54982 576183 54984
rect 461780 54980 461786 54982
rect 576117 54979 576183 54982
rect 574461 54770 574527 54773
rect 459878 54768 574527 54770
rect 459878 54712 574466 54768
rect 574522 54712 574527 54768
rect 459878 54710 574527 54712
rect 459878 53685 459938 54710
rect 574461 54707 574527 54710
rect 591297 54498 591363 54501
rect 466410 54496 591363 54498
rect 466410 54440 591302 54496
rect 591358 54440 591363 54496
rect 466410 54438 591363 54440
rect 466410 54226 466470 54438
rect 591297 54435 591363 54438
rect 577497 54226 577563 54229
rect 460798 54166 466470 54226
rect 469170 54224 577563 54226
rect 469170 54168 577502 54224
rect 577558 54168 577563 54224
rect 469170 54166 577563 54168
rect 460798 53685 460858 54166
rect 461710 53892 461716 53956
rect 461780 53892 461786 53956
rect 469170 53954 469230 54166
rect 577497 54163 577563 54166
rect 462638 53894 469230 53954
rect 461718 53685 461778 53892
rect 462638 53685 462698 53894
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462589 53680 462698 53685
rect 462589 53624 462594 53680
rect 462650 53624 462698 53680
rect 462589 53622 462698 53624
rect 470317 53682 470383 53685
rect 471973 53682 472039 53685
rect 470317 53680 472039 53682
rect 470317 53624 470322 53680
rect 470378 53624 471978 53680
rect 472034 53624 472039 53680
rect 470317 53622 472039 53624
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53619 462655 53622
rect 470317 53619 470383 53622
rect 471973 53619 472039 53622
rect 470961 53410 471027 53413
rect 476757 53410 476823 53413
rect 470961 53408 476823 53410
rect 470961 53352 470966 53408
rect 471022 53352 476762 53408
rect 476818 53352 476823 53408
rect 470961 53350 476823 53352
rect 470961 53347 471027 53350
rect 476757 53347 476823 53350
rect 463877 53138 463943 53141
rect 471145 53138 471211 53141
rect 463877 53136 471211 53138
rect 463877 53080 463882 53136
rect 463938 53080 471150 53136
rect 471206 53080 471211 53136
rect 463877 53078 471211 53080
rect 463877 53075 463943 53078
rect 471145 53075 471211 53078
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 661585 48512 661651 48515
rect 661480 48510 661651 48512
rect 661480 48454 661590 48510
rect 661646 48454 661651 48510
rect 661480 48452 661651 48454
rect 661585 48449 661651 48452
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 661769 47791 661835 47794
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 661388 47789 661835 47791
rect 661388 47733 661774 47789
rect 661830 47733 661835 47789
rect 661388 47731 661835 47733
rect 661769 47728 661835 47731
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 465073 46746 465139 46749
rect 458357 46744 465139 46746
rect 458357 46688 458362 46744
rect 458418 46688 465078 46744
rect 465134 46688 465139 46744
rect 458357 46686 465139 46688
rect 458357 46683 458423 46686
rect 465073 46683 465139 46686
rect 463918 44508 463924 44572
rect 463988 44570 463994 44572
rect 464705 44570 464771 44573
rect 463988 44568 464771 44570
rect 463988 44512 464710 44568
rect 464766 44512 464771 44568
rect 463988 44510 464771 44512
rect 463988 44508 463994 44510
rect 464705 44507 464771 44510
rect 458173 44434 458239 44437
rect 461025 44434 461091 44437
rect 458173 44432 461091 44434
rect 458173 44376 458178 44432
rect 458234 44376 461030 44432
rect 461086 44376 461091 44432
rect 458173 44374 461091 44376
rect 458173 44371 458239 44374
rect 461025 44371 461091 44374
rect 463693 44436 463759 44437
rect 463693 44432 463740 44436
rect 463804 44434 463810 44436
rect 463693 44376 463698 44432
rect 463693 44372 463740 44376
rect 463804 44374 463850 44434
rect 463804 44372 463810 44374
rect 463693 44371 463759 44372
rect 129089 44298 129155 44301
rect 131941 44298 132007 44301
rect 142613 44298 142679 44301
rect 129089 44296 132007 44298
rect 129089 44240 129094 44296
rect 129150 44240 131946 44296
rect 132002 44240 132007 44296
rect 129089 44238 132007 44240
rect 129089 44235 129155 44238
rect 131941 44235 132007 44238
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 307293 44162 307359 44165
rect 463877 44162 463943 44165
rect 307293 44160 463943 44162
rect 307293 44104 307298 44160
rect 307354 44104 463882 44160
rect 463938 44104 463943 44160
rect 307293 44102 463943 44104
rect 307293 44099 307359 44102
rect 463877 44099 463943 44102
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 460841 43890 460907 43893
rect 471053 43890 471119 43893
rect 460841 43888 471119 43890
rect 460841 43832 460846 43888
rect 460902 43832 471058 43888
rect 471114 43832 471119 43888
rect 460841 43830 471119 43832
rect 460841 43827 460907 43830
rect 471053 43827 471119 43830
rect 419717 43618 419783 43621
rect 440233 43618 440299 43621
rect 419717 43616 440299 43618
rect 419717 43560 419722 43616
rect 419778 43560 440238 43616
rect 440294 43560 440299 43616
rect 419717 43558 440299 43560
rect 419717 43555 419783 43558
rect 440233 43555 440299 43558
rect 441061 43618 441127 43621
rect 462865 43618 462931 43621
rect 441061 43616 462931 43618
rect 441061 43560 441066 43616
rect 441122 43560 462870 43616
rect 462926 43560 462931 43616
rect 441061 43558 462931 43560
rect 441061 43555 441127 43558
rect 462865 43555 462931 43558
rect 462681 43210 462747 43213
rect 465809 43210 465875 43213
rect 462681 43208 465875 43210
rect 462681 43152 462686 43208
rect 462742 43152 465814 43208
rect 465870 43152 465875 43208
rect 462681 43150 465875 43152
rect 462681 43147 462747 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463969 42938 464035 42941
rect 461761 42936 464035 42938
rect 461761 42880 461766 42936
rect 461822 42880 463974 42936
rect 464030 42880 464035 42936
rect 461761 42878 464035 42880
rect 461761 42875 461827 42878
rect 463969 42875 464035 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 416589 42396 416655 42397
rect 416589 42392 416636 42396
rect 416700 42394 416706 42396
rect 416589 42336 416594 42392
rect 416589 42332 416636 42336
rect 416700 42334 416746 42394
rect 416700 42332 416706 42334
rect 416589 42331 416655 42332
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 404629 42122 404695 42125
rect 405181 42122 405247 42125
rect 404629 42120 405247 42122
rect 404629 42064 404634 42120
rect 404690 42064 405186 42120
rect 405242 42064 405247 42120
rect 404629 42062 405247 42064
rect 194317 42059 194383 42060
rect 404629 42059 404695 42062
rect 405181 42059 405247 42062
rect 415577 42122 415643 42125
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 415577 42120 422310 42122
rect 415577 42064 415582 42120
rect 415638 42064 422310 42120
rect 415577 42062 422310 42064
rect 415577 42059 415643 42062
rect 310421 41850 310487 41853
rect 311065 41850 311131 41853
rect 310421 41848 311131 41850
rect 310421 41792 310426 41848
rect 310482 41792 311070 41848
rect 311126 41792 311131 41848
rect 310421 41790 311131 41792
rect 310421 41787 310487 41790
rect 311065 41787 311131 41790
rect 361941 41852 362007 41853
rect 361941 41848 361988 41852
rect 362052 41850 362058 41852
rect 365161 41850 365227 41853
rect 365662 41850 365668 41852
rect 361941 41792 361946 41848
rect 361941 41788 361988 41792
rect 362052 41790 362098 41850
rect 365161 41848 365668 41850
rect 365161 41792 365166 41848
rect 365222 41792 365668 41848
rect 365161 41790 365668 41792
rect 362052 41788 362058 41790
rect 361941 41787 362007 41788
rect 365161 41787 365227 41790
rect 365662 41788 365668 41790
rect 365732 41788 365738 41852
rect 402830 41788 402836 41852
rect 402900 41850 402906 41852
rect 421966 41850 421972 41852
rect 402900 41790 421972 41850
rect 402900 41788 402906 41790
rect 421966 41788 421972 41790
rect 422036 41788 422042 41852
rect 422250 41578 422310 42062
rect 460974 42060 460980 42124
rect 461044 42122 461050 42124
rect 463918 42122 463924 42124
rect 461044 42062 463924 42122
rect 461044 42060 461050 42062
rect 463918 42060 463924 42062
rect 463988 42060 463994 42124
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 451222 41788 451228 41852
rect 451292 41850 451298 41852
rect 460606 41850 460612 41852
rect 451292 41790 460612 41850
rect 451292 41788 451298 41790
rect 460606 41788 460612 41790
rect 460676 41788 460682 41852
rect 461945 41850 462011 41853
rect 460890 41848 462011 41850
rect 460890 41792 461950 41848
rect 462006 41792 462011 41848
rect 460890 41790 462011 41792
rect 422250 41518 441630 41578
rect 441570 41442 441630 41518
rect 460890 41442 460950 41790
rect 461945 41787 462011 41790
rect 441570 41382 460950 41442
rect 425838 41246 431970 41306
rect 416630 40428 416636 40492
rect 416700 40490 416706 40492
rect 425838 40490 425898 41246
rect 431910 41170 431970 41246
rect 458173 41170 458239 41173
rect 431910 41168 458239 41170
rect 431910 41112 458178 41168
rect 458234 41112 458239 41168
rect 431910 41110 458239 41112
rect 458173 41107 458239 41110
rect 416700 40430 425898 40490
rect 416700 40428 416706 40430
rect 141693 40356 141759 40357
rect 141693 40352 141740 40356
rect 141804 40354 141810 40356
rect 141693 40296 141698 40352
rect 141693 40292 141740 40296
rect 141804 40294 141850 40354
rect 141804 40292 141810 40294
rect 141693 40291 141759 40292
<< via3 >>
rect 675892 892196 675956 892260
rect 675892 887708 675956 887772
rect 675708 885804 675772 885868
rect 675524 880636 675588 880700
rect 676260 880364 676324 880428
rect 675340 878460 675404 878524
rect 675340 874108 675404 874172
rect 676444 873020 676508 873084
rect 676260 872748 676324 872812
rect 675708 865676 675772 865740
rect 676076 865404 676140 865468
rect 675892 864996 675956 865060
rect 41828 813180 41892 813244
rect 41828 811956 41892 812020
rect 41644 805564 41708 805628
rect 40908 805156 40972 805220
rect 40724 804884 40788 804948
rect 40540 804612 40604 804676
rect 40356 800804 40420 800868
rect 41092 800532 41156 800596
rect 42012 800320 42076 800324
rect 42012 800264 42026 800320
rect 42026 800264 42076 800320
rect 42012 800260 42076 800264
rect 40356 796180 40420 796244
rect 41092 794412 41156 794476
rect 42012 792976 42076 792980
rect 42012 792920 42062 792976
rect 42062 792920 42076 792976
rect 42012 792916 42076 792920
rect 41828 791556 41892 791620
rect 40724 791284 40788 791348
rect 40908 790604 40972 790668
rect 41644 788156 41708 788220
rect 41460 786796 41524 786860
rect 676076 786660 676140 786724
rect 40540 786116 40604 786180
rect 674236 783804 674300 783868
rect 674604 782444 674668 782508
rect 41460 769796 41524 769860
rect 40724 766532 40788 766596
rect 40540 765308 40604 765372
rect 40908 764900 40972 764964
rect 42012 759052 42076 759116
rect 42196 758976 42260 758980
rect 42196 758920 42210 758976
rect 42210 758920 42260 758976
rect 42196 758916 42260 758920
rect 41644 757692 41708 757756
rect 41828 757072 41892 757076
rect 41828 757016 41842 757072
rect 41842 757016 41892 757072
rect 41828 757012 41892 757016
rect 41828 755440 41892 755444
rect 41828 755384 41878 755440
rect 41878 755384 41892 755440
rect 41828 755380 41892 755384
rect 40908 754836 40972 754900
rect 41828 754836 41892 754900
rect 42196 754896 42260 754900
rect 42196 754840 42210 754896
rect 42210 754840 42260 754896
rect 42196 754836 42260 754840
rect 41828 750408 41892 750412
rect 41828 750352 41842 750408
rect 41842 750352 41892 750408
rect 41828 750348 41892 750352
rect 40540 749532 40604 749596
rect 40724 746676 40788 746740
rect 41644 745044 41708 745108
rect 42012 744832 42076 744836
rect 42012 744776 42062 744832
rect 42062 744776 42076 744832
rect 42012 744772 42076 744776
rect 41460 743684 41524 743748
rect 676812 739740 676876 739804
rect 674420 738108 674484 738172
rect 676076 726820 676140 726884
rect 674236 726412 674300 726476
rect 41828 725792 41892 725796
rect 41828 725736 41842 725792
rect 41842 725736 41892 725792
rect 41828 725732 41892 725736
rect 674788 722256 674852 722260
rect 674788 722200 674838 722256
rect 674838 722200 674852 722256
rect 674788 722196 674852 722200
rect 676076 721516 676140 721580
rect 40724 718524 40788 718588
rect 41644 718252 41708 718316
rect 40540 717980 40604 718044
rect 41828 716076 41892 716140
rect 41276 714232 41340 714236
rect 41276 714176 41290 714232
rect 41290 714176 41340 714232
rect 41276 714172 41340 714176
rect 41276 712132 41340 712196
rect 674604 707508 674668 707572
rect 40724 707372 40788 707436
rect 674604 706284 674668 706348
rect 40540 706148 40604 706212
rect 41828 702068 41892 702132
rect 41644 701796 41708 701860
rect 41460 700436 41524 700500
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 675340 687108 675404 687172
rect 676996 686156 677060 686220
rect 41828 683572 41892 683636
rect 675892 682076 675956 682140
rect 676076 681804 676140 681868
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 41828 678872 41892 678876
rect 41828 678816 41842 678872
rect 41842 678816 41892 678872
rect 41828 678812 41892 678816
rect 40908 677750 40972 677754
rect 40908 677694 40958 677750
rect 40958 677694 40972 677750
rect 40908 677690 40972 677694
rect 676076 676364 676140 676428
rect 41092 672964 41156 673028
rect 41828 672692 41892 672756
rect 43300 671936 43364 671940
rect 43300 671880 43314 671936
rect 43314 671880 43364 671936
rect 43300 671876 43364 671880
rect 40356 670924 40420 670988
rect 41092 669020 41156 669084
rect 42196 667388 42260 667452
rect 43300 666844 43364 666908
rect 42196 666632 42260 666636
rect 42196 666576 42210 666632
rect 42210 666576 42260 666632
rect 42196 666572 42260 666576
rect 40356 665484 40420 665548
rect 40908 665212 40972 665276
rect 676812 664124 676876 664188
rect 40724 663988 40788 664052
rect 40540 662628 40604 662692
rect 674420 662356 674484 662420
rect 41460 660860 41524 660924
rect 41644 658548 41708 658612
rect 41828 658336 41892 658340
rect 41828 658280 41842 658336
rect 41842 658280 41892 658336
rect 41828 658276 41892 658280
rect 674236 649708 674300 649772
rect 676812 648620 676876 648684
rect 674788 643996 674852 644060
rect 44220 642228 44284 642292
rect 41644 640596 41708 640660
rect 674788 640188 674852 640252
rect 41460 639372 41524 639436
rect 40540 637332 40604 637396
rect 676076 636108 676140 636172
rect 40724 635292 40788 635356
rect 40908 634884 40972 634948
rect 42380 632844 42444 632908
rect 41828 629852 41892 629916
rect 42196 625696 42260 625700
rect 42196 625640 42246 625696
rect 42246 625640 42260 625696
rect 42196 625636 42260 625640
rect 42380 624548 42444 624612
rect 40908 623732 40972 623796
rect 676996 621556 677060 621620
rect 40724 620876 40788 620940
rect 42196 619788 42260 619852
rect 40540 616388 40604 616452
rect 41828 616116 41892 616180
rect 674420 616116 674484 616180
rect 41644 615708 41708 615772
rect 41460 615164 41524 615228
rect 675340 608288 675404 608292
rect 675340 608232 675390 608288
rect 675390 608232 675404 608288
rect 675340 608228 675404 608232
rect 675524 604616 675588 604620
rect 675524 604560 675538 604616
rect 675538 604560 675588 604616
rect 675524 604556 675588 604560
rect 44220 599660 44284 599724
rect 43116 599252 43180 599316
rect 676996 598844 677060 598908
rect 42012 597212 42076 597276
rect 43116 597000 43180 597004
rect 43116 596944 43166 597000
rect 43166 596944 43180 597000
rect 43116 596940 43180 596944
rect 42196 596396 42260 596460
rect 675524 596260 675588 596324
rect 41828 593948 41892 594012
rect 40724 592894 40788 592958
rect 674236 592588 674300 592652
rect 41460 592078 41524 592142
rect 675524 592104 675588 592108
rect 675524 592048 675538 592104
rect 675538 592048 675588 592104
rect 675524 592044 675588 592048
rect 40356 590854 40420 590918
rect 40356 589596 40420 589660
rect 42196 587556 42260 587620
rect 675156 586256 675220 586260
rect 675156 586200 675170 586256
rect 675170 586200 675220 586256
rect 675156 586196 675220 586200
rect 676076 586196 676140 586260
rect 40356 585924 40420 585988
rect 41828 585108 41892 585172
rect 42196 581904 42260 581908
rect 42196 581848 42210 581904
rect 42210 581848 42260 581904
rect 42196 581844 42260 581848
rect 40356 580212 40420 580276
rect 40908 577764 40972 577828
rect 40540 575588 40604 575652
rect 676996 575180 677060 575244
rect 40724 574636 40788 574700
rect 676812 573548 676876 573612
rect 41460 572732 41524 572796
rect 41644 571508 41708 571572
rect 671476 570692 671540 570756
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 673868 565524 673932 565588
rect 676444 562668 676508 562732
rect 675340 561912 675404 561916
rect 675340 561856 675390 561912
rect 675390 561856 675404 561912
rect 675340 561852 675404 561856
rect 41092 558724 41156 558788
rect 41092 557488 41156 557552
rect 41828 553964 41892 554028
rect 676812 553828 676876 553892
rect 41828 552740 41892 552804
rect 676996 552060 677060 552124
rect 676444 547572 676508 547636
rect 675892 547300 675956 547364
rect 676076 547028 676140 547092
rect 41644 546348 41708 546412
rect 40724 545668 40788 545732
rect 40540 545396 40604 545460
rect 675340 544504 675404 544508
rect 675340 544448 675354 544504
rect 675354 544448 675404 544504
rect 675340 544444 675404 544448
rect 40540 537372 40604 537436
rect 40724 536964 40788 537028
rect 41460 530708 41524 530772
rect 41644 529484 41708 529548
rect 41828 529000 41892 529004
rect 41828 528944 41842 529000
rect 41842 528944 41892 529000
rect 41828 528940 41892 528944
rect 675708 488820 675772 488884
rect 675892 483924 675956 483988
rect 675524 483516 675588 483580
rect 674604 477396 674668 477460
rect 673684 475356 673748 475420
rect 674420 475356 674484 475420
rect 671476 474812 671540 474876
rect 673684 464748 673748 464812
rect 673868 454956 673932 455020
rect 675340 447748 675404 447812
rect 676812 440268 676876 440332
rect 41828 426396 41892 426460
rect 42012 424764 42076 424828
rect 42196 424220 42260 424284
rect 41828 422724 41892 422788
rect 41828 421908 41892 421972
rect 41460 418780 41524 418844
rect 41644 413340 41708 413404
rect 42196 413340 42260 413404
rect 675340 410484 675404 410548
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40908 405588 40972 405652
rect 41828 401840 41892 401844
rect 41828 401784 41842 401840
rect 41842 401784 41892 401840
rect 41828 401780 41892 401784
rect 677180 401236 677244 401300
rect 676812 400420 676876 400484
rect 40540 400012 40604 400076
rect 41460 398788 41524 398852
rect 676076 398788 676140 398852
rect 676260 396748 676324 396812
rect 676444 395932 676508 395996
rect 676628 395116 676692 395180
rect 675892 389812 675956 389876
rect 675708 388452 675772 388516
rect 676260 385324 676324 385388
rect 676444 381652 676508 381716
rect 40540 380564 40604 380628
rect 41460 379748 41524 379812
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40724 378116 40788 378180
rect 676628 377300 676692 377364
rect 41276 374580 41340 374644
rect 676076 373628 676140 373692
rect 41644 372676 41708 372740
rect 675892 372948 675956 373012
rect 41828 371860 41892 371924
rect 41276 368460 41340 368524
rect 40724 363700 40788 363764
rect 41828 360088 41892 360092
rect 41828 360032 41842 360088
rect 41842 360032 41892 360088
rect 41828 360028 41892 360032
rect 41644 359484 41708 359548
rect 41460 358668 41524 358732
rect 40540 356084 40604 356148
rect 675524 353364 675588 353428
rect 675708 352956 675772 353020
rect 675938 352140 676002 352204
rect 675892 351928 675956 351932
rect 675892 351872 675906 351928
rect 675906 351872 675956 351928
rect 675892 351868 675956 351872
rect 676444 346624 676508 346628
rect 676444 346568 676494 346624
rect 676494 346568 676508 346624
rect 676444 346564 676508 346568
rect 676812 346156 676876 346220
rect 44404 342892 44468 342956
rect 44220 341532 44284 341596
rect 675524 340776 675588 340780
rect 675524 340720 675574 340776
rect 675574 340720 675588 340776
rect 675524 340716 675588 340720
rect 42748 340444 42812 340508
rect 44588 340172 44652 340236
rect 676444 340172 676508 340236
rect 41644 338132 41708 338196
rect 675892 337724 675956 337788
rect 42932 337588 42996 337652
rect 43116 337180 43180 337244
rect 40724 336908 40788 336972
rect 42012 336500 42076 336564
rect 41828 335684 41892 335748
rect 40540 335276 40604 335340
rect 40908 333644 40972 333708
rect 676076 328340 676140 328404
rect 676260 325484 676324 325548
rect 40908 325348 40972 325412
rect 676812 325212 676876 325276
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 41828 319968 41892 319972
rect 41828 319912 41878 319968
rect 41878 319912 41892 319968
rect 41828 319908 41892 319912
rect 40724 318956 40788 319020
rect 40540 317324 40604 317388
rect 43116 315964 43180 316028
rect 42012 313712 42076 313716
rect 42012 313656 42062 313712
rect 42062 313656 42076 313712
rect 42012 313652 42076 313656
rect 42932 312700 42996 312764
rect 675708 309028 675772 309092
rect 675708 308756 675772 308820
rect 675892 307124 675956 307188
rect 676444 301608 676508 301612
rect 676444 301552 676494 301608
rect 676494 301552 676508 301608
rect 676444 301548 676508 301552
rect 676260 300596 676324 300660
rect 44404 300052 44468 300116
rect 675708 299372 675772 299436
rect 44588 299236 44652 299300
rect 44220 298420 44284 298484
rect 42748 297604 42812 297668
rect 42012 296788 42076 296852
rect 675340 296788 675404 296852
rect 675524 296516 675588 296580
rect 675340 295292 675404 295356
rect 676628 294476 676692 294540
rect 41368 292528 41432 292592
rect 675524 292224 675588 292228
rect 675524 292168 675574 292224
rect 675574 292168 675588 292224
rect 675524 292164 675588 292168
rect 41828 291484 41892 291548
rect 676444 291484 676508 291548
rect 676260 290804 676324 290868
rect 40724 289172 40788 289236
rect 41644 284820 41708 284884
rect 42012 284276 42076 284340
rect 675892 283596 675956 283660
rect 675708 282840 675772 282844
rect 675708 282784 675722 282840
rect 675722 282784 675772 282840
rect 675708 282780 675772 282784
rect 676076 281148 676140 281212
rect 40908 278428 40972 278492
rect 40724 277068 40788 277132
rect 40540 274212 40604 274276
rect 42012 272368 42076 272372
rect 42012 272312 42026 272368
rect 42026 272312 42076 272368
rect 42012 272308 42076 272312
rect 41460 270404 41524 270468
rect 41828 270056 41892 270060
rect 41828 270000 41878 270056
rect 41878 270000 41892 270056
rect 41828 269996 41892 270000
rect 674972 264148 675036 264212
rect 676076 263604 676140 263668
rect 676812 261564 676876 261628
rect 676996 259932 677060 259996
rect 40540 250140 40604 250204
rect 676812 250140 676876 250204
rect 40724 249732 40788 249796
rect 674972 249732 675036 249796
rect 676076 249596 676140 249660
rect 673316 246196 673380 246260
rect 676996 242252 677060 242316
rect 676812 241844 676876 241908
rect 674972 241572 675036 241636
rect 42012 237356 42076 237420
rect 40724 236540 40788 236604
rect 40540 233004 40604 233068
rect 674972 230148 675036 230212
rect 674052 229740 674116 229804
rect 42012 228984 42076 228988
rect 42012 228928 42026 228984
rect 42026 228928 42076 228984
rect 42012 228924 42076 228928
rect 671108 224768 671172 224772
rect 671108 224712 671158 224768
rect 671158 224712 671172 224768
rect 671108 224708 671172 224712
rect 671108 223136 671172 223140
rect 671108 223080 671158 223136
rect 671158 223080 671172 223136
rect 671108 223076 671172 223080
rect 674236 221852 674300 221916
rect 675892 220628 675956 220692
rect 675892 218180 675956 218244
rect 509188 217772 509252 217836
rect 510108 217832 510172 217836
rect 510108 217776 510158 217832
rect 510158 217776 510172 217832
rect 510108 217772 510172 217776
rect 522620 217832 522684 217836
rect 522620 217776 522634 217832
rect 522634 217776 522684 217832
rect 522620 217772 522684 217776
rect 566964 217832 567028 217836
rect 566964 217776 566978 217832
rect 566978 217776 567028 217832
rect 566964 217772 567028 217776
rect 574324 217772 574388 217836
rect 675708 217364 675772 217428
rect 493732 217288 493796 217292
rect 493732 217232 493782 217288
rect 493782 217232 493796 217288
rect 493732 217228 493796 217232
rect 574324 216684 574388 216748
rect 566964 216140 567028 216204
rect 509188 215868 509252 215932
rect 522620 215324 522684 215388
rect 673684 215248 673748 215252
rect 673684 215192 673698 215248
rect 673698 215192 673748 215248
rect 673684 215188 673748 215192
rect 675892 215188 675956 215252
rect 675892 214372 675956 214436
rect 674236 212740 674300 212804
rect 676260 210836 676324 210900
rect 676628 210836 676692 210900
rect 675892 210564 675956 210628
rect 670740 210488 670804 210492
rect 670740 210432 670790 210488
rect 670790 210432 670804 210488
rect 670740 210428 670804 210432
rect 41828 210020 41892 210084
rect 41460 208116 41524 208180
rect 40540 207300 40604 207364
rect 676076 206892 676140 206956
rect 40724 206484 40788 206548
rect 40908 206076 40972 206140
rect 41644 205668 41708 205732
rect 676444 205532 676508 205596
rect 676076 204172 676140 204236
rect 676260 200636 676324 200700
rect 675708 198384 675772 198388
rect 675708 198328 675758 198384
rect 675758 198328 675772 198384
rect 675708 198324 675772 198328
rect 676628 196012 676692 196076
rect 41828 195256 41892 195260
rect 41828 195200 41878 195256
rect 41878 195200 41892 195256
rect 41828 195196 41892 195200
rect 40908 194924 40972 194988
rect 40724 193156 40788 193220
rect 675892 192612 675956 192676
rect 40540 186356 40604 186420
rect 41460 185948 41524 186012
rect 41828 184104 41892 184108
rect 41828 184048 41842 184104
rect 41842 184048 41892 184104
rect 41828 184044 41892 184048
rect 675524 173572 675588 173636
rect 675892 172756 675956 172820
rect 675708 172348 675772 172412
rect 669452 170988 669516 171052
rect 675892 169628 675956 169692
rect 675708 167452 675772 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 675524 162148 675588 162212
rect 676076 162148 676140 162212
rect 673316 161332 673380 161396
rect 676444 156980 676508 157044
rect 676260 155620 676324 155684
rect 675892 153036 675956 153100
rect 676628 151404 676692 151468
rect 676076 148412 676140 148476
rect 675708 147656 675772 147660
rect 675708 147600 675722 147656
rect 675722 147600 675772 147656
rect 675708 147596 675772 147600
rect 669268 140388 669332 140452
rect 674052 132908 674116 132972
rect 673500 132636 673564 132700
rect 676444 127332 676508 127396
rect 675892 127196 675956 127260
rect 676076 126108 676140 126172
rect 670740 125700 670804 125764
rect 676260 124476 676324 124540
rect 676812 122844 676876 122908
rect 675708 116044 675772 116108
rect 676812 114276 676876 114340
rect 676444 112372 676508 112436
rect 676260 110332 676324 110396
rect 675892 108020 675956 108084
rect 676076 103124 676140 103188
rect 675708 102640 675772 102644
rect 675708 102584 675722 102640
rect 675722 102584 675772 102640
rect 675708 102580 675772 102584
rect 635780 96868 635844 96932
rect 637252 96868 637316 96932
rect 647188 96460 647252 96524
rect 633940 95916 634004 95980
rect 650316 93060 650380 93124
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 635780 78100 635844 78164
rect 637068 77556 637132 77620
rect 461716 54980 461780 55044
rect 461716 53892 461780 53956
rect 194364 50220 194428 50284
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 463924 44508 463988 44572
rect 463740 44432 463804 44436
rect 463740 44376 463754 44432
rect 463754 44376 463804 44432
rect 463740 44372 463804 44376
rect 141740 43964 141804 44028
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 416636 42392 416700 42396
rect 416636 42336 416650 42392
rect 416650 42336 416700 42392
rect 416636 42332 416700 42336
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 361988 41848 362052 41852
rect 361988 41792 362002 41848
rect 362002 41792 362052 41848
rect 361988 41788 362052 41792
rect 365668 41788 365732 41852
rect 402836 41788 402900 41852
rect 421972 41788 422036 41852
rect 460980 42060 461044 42124
rect 463924 42060 463988 42124
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 451228 41788 451292 41852
rect 460612 41788 460676 41852
rect 416636 40428 416700 40492
rect 141740 40352 141804 40356
rect 141740 40296 141754 40352
rect 141754 40296 141804 40352
rect 141740 40292 141804 40296
<< metal4 >>
rect 675891 892260 675957 892261
rect 675891 892196 675892 892260
rect 675956 892196 675957 892260
rect 675891 892195 675957 892196
rect 675894 891510 675954 892195
rect 675710 891450 675954 891510
rect 675710 887090 675770 891450
rect 675891 887772 675957 887773
rect 675891 887708 675892 887772
rect 675956 887770 675957 887772
rect 675956 887710 676322 887770
rect 675956 887708 675957 887710
rect 675891 887707 675957 887708
rect 675710 887030 675954 887090
rect 675707 885868 675773 885869
rect 675707 885804 675708 885868
rect 675772 885804 675773 885868
rect 675707 885803 675773 885804
rect 675523 880700 675589 880701
rect 675523 880636 675524 880700
rect 675588 880636 675589 880700
rect 675523 880635 675589 880636
rect 675339 878524 675405 878525
rect 675339 878460 675340 878524
rect 675404 878460 675405 878524
rect 675339 878459 675405 878460
rect 675342 874173 675402 878459
rect 675339 874172 675405 874173
rect 675339 874108 675340 874172
rect 675404 874108 675405 874172
rect 675339 874107 675405 874108
rect 675526 872190 675586 880635
rect 675710 876890 675770 885803
rect 675894 881850 675954 887030
rect 676262 881850 676322 887710
rect 675894 881790 676138 881850
rect 676262 881790 676506 881850
rect 675710 876830 675954 876890
rect 675526 872130 675770 872190
rect 675710 865741 675770 872130
rect 675707 865740 675773 865741
rect 675707 865676 675708 865740
rect 675772 865676 675773 865740
rect 675707 865675 675773 865676
rect 675894 865061 675954 876830
rect 676078 865469 676138 881790
rect 676259 880428 676325 880429
rect 676259 880364 676260 880428
rect 676324 880364 676325 880428
rect 676259 880363 676325 880364
rect 676262 872813 676322 880363
rect 676446 873085 676506 881790
rect 676443 873084 676509 873085
rect 676443 873020 676444 873084
rect 676508 873020 676509 873084
rect 676443 873019 676509 873020
rect 676259 872812 676325 872813
rect 676259 872748 676260 872812
rect 676324 872748 676325 872812
rect 676259 872747 676325 872748
rect 676075 865468 676141 865469
rect 676075 865404 676076 865468
rect 676140 865404 676141 865468
rect 676075 865403 676141 865404
rect 675891 865060 675957 865061
rect 675891 864996 675892 865060
rect 675956 864996 675957 865060
rect 675891 864995 675957 864996
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40907 805220 40973 805221
rect 40907 805156 40908 805220
rect 40972 805156 40973 805220
rect 40907 805155 40973 805156
rect 40723 804948 40789 804949
rect 40723 804884 40724 804948
rect 40788 804884 40789 804948
rect 40723 804883 40789 804884
rect 40539 804676 40605 804677
rect 40539 804612 40540 804676
rect 40604 804612 40605 804676
rect 40539 804611 40605 804612
rect 40355 800868 40421 800869
rect 40355 800804 40356 800868
rect 40420 800804 40421 800868
rect 40355 800803 40421 800804
rect 40358 796245 40418 800803
rect 40355 796244 40421 796245
rect 40355 796180 40356 796244
rect 40420 796180 40421 796244
rect 40355 796179 40421 796180
rect 40542 786181 40602 804611
rect 40726 791349 40786 804883
rect 40723 791348 40789 791349
rect 40723 791284 40724 791348
rect 40788 791284 40789 791348
rect 40723 791283 40789 791284
rect 40910 790669 40970 805155
rect 41091 800596 41157 800597
rect 41091 800532 41092 800596
rect 41156 800532 41157 800596
rect 41091 800531 41157 800532
rect 41094 794477 41154 800531
rect 41091 794476 41157 794477
rect 41091 794412 41092 794476
rect 41156 794412 41157 794476
rect 41091 794411 41157 794412
rect 40907 790668 40973 790669
rect 40907 790604 40908 790668
rect 40972 790604 40973 790668
rect 40907 790603 40973 790604
rect 41462 786861 41522 812910
rect 41827 812020 41893 812021
rect 41827 811956 41828 812020
rect 41892 811956 41893 812020
rect 41827 811955 41893 811956
rect 41643 805628 41709 805629
rect 41643 805564 41644 805628
rect 41708 805564 41709 805628
rect 41643 805563 41709 805564
rect 41646 788221 41706 805563
rect 41830 791621 41890 811955
rect 42011 800324 42077 800325
rect 42011 800260 42012 800324
rect 42076 800260 42077 800324
rect 42011 800259 42077 800260
rect 42014 792981 42074 800259
rect 42011 792980 42077 792981
rect 42011 792916 42012 792980
rect 42076 792916 42077 792980
rect 42011 792915 42077 792916
rect 41827 791620 41893 791621
rect 41827 791556 41828 791620
rect 41892 791556 41893 791620
rect 41827 791555 41893 791556
rect 41643 788220 41709 788221
rect 41643 788156 41644 788220
rect 41708 788156 41709 788220
rect 41643 788155 41709 788156
rect 41459 786860 41525 786861
rect 41459 786796 41460 786860
rect 41524 786796 41525 786860
rect 41459 786795 41525 786796
rect 676075 786724 676141 786725
rect 676075 786660 676076 786724
rect 676140 786660 676141 786724
rect 676075 786659 676141 786660
rect 40539 786180 40605 786181
rect 40539 786116 40540 786180
rect 40604 786116 40605 786180
rect 40539 786115 40605 786116
rect 674235 783868 674301 783869
rect 674235 783804 674236 783868
rect 674300 783804 674301 783868
rect 674235 783803 674301 783804
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40723 766596 40789 766597
rect 40723 766532 40724 766596
rect 40788 766532 40789 766596
rect 40723 766531 40789 766532
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40542 749597 40602 765307
rect 40539 749596 40605 749597
rect 40539 749532 40540 749596
rect 40604 749532 40605 749596
rect 40539 749531 40605 749532
rect 40726 746741 40786 766531
rect 40907 764964 40973 764965
rect 40907 764900 40908 764964
rect 40972 764900 40973 764964
rect 40907 764899 40973 764900
rect 40910 754901 40970 764899
rect 40907 754900 40973 754901
rect 40907 754836 40908 754900
rect 40972 754836 40973 754900
rect 40907 754835 40973 754836
rect 40723 746740 40789 746741
rect 40723 746676 40724 746740
rect 40788 746676 40789 746740
rect 40723 746675 40789 746676
rect 41462 743749 41522 769795
rect 42011 759116 42077 759117
rect 42011 759052 42012 759116
rect 42076 759052 42077 759116
rect 42011 759051 42077 759052
rect 41643 757756 41709 757757
rect 41643 757692 41644 757756
rect 41708 757692 41709 757756
rect 41643 757691 41709 757692
rect 41646 745109 41706 757691
rect 41827 757076 41893 757077
rect 41827 757012 41828 757076
rect 41892 757012 41893 757076
rect 41827 757011 41893 757012
rect 41830 755445 41890 757011
rect 41827 755444 41893 755445
rect 41827 755380 41828 755444
rect 41892 755380 41893 755444
rect 41827 755379 41893 755380
rect 41827 754900 41893 754901
rect 41827 754836 41828 754900
rect 41892 754836 41893 754900
rect 41827 754835 41893 754836
rect 41830 750413 41890 754835
rect 41827 750412 41893 750413
rect 41827 750348 41828 750412
rect 41892 750348 41893 750412
rect 41827 750347 41893 750348
rect 41643 745108 41709 745109
rect 41643 745044 41644 745108
rect 41708 745044 41709 745108
rect 41643 745043 41709 745044
rect 42014 744837 42074 759051
rect 42195 758980 42261 758981
rect 42195 758916 42196 758980
rect 42260 758916 42261 758980
rect 42195 758915 42261 758916
rect 42198 754901 42258 758915
rect 42195 754900 42261 754901
rect 42195 754836 42196 754900
rect 42260 754836 42261 754900
rect 42195 754835 42261 754836
rect 42011 744836 42077 744837
rect 42011 744772 42012 744836
rect 42076 744772 42077 744836
rect 42011 744771 42077 744772
rect 41459 743748 41525 743749
rect 41459 743684 41460 743748
rect 41524 743684 41525 743748
rect 41459 743683 41525 743684
rect 674238 726477 674298 783803
rect 674603 782508 674669 782509
rect 674603 782444 674604 782508
rect 674668 782444 674669 782508
rect 674603 782443 674669 782444
rect 674419 738172 674485 738173
rect 674419 738108 674420 738172
rect 674484 738108 674485 738172
rect 674419 738107 674485 738108
rect 674235 726476 674301 726477
rect 674235 726412 674236 726476
rect 674300 726412 674301 726476
rect 674235 726411 674301 726412
rect 41827 725796 41893 725797
rect 41827 725732 41828 725796
rect 41892 725732 41893 725796
rect 41827 725731 41893 725732
rect 41830 725250 41890 725731
rect 41462 725190 41890 725250
rect 40723 718588 40789 718589
rect 40723 718524 40724 718588
rect 40788 718524 40789 718588
rect 40723 718523 40789 718524
rect 40539 718044 40605 718045
rect 40539 717980 40540 718044
rect 40604 717980 40605 718044
rect 40539 717979 40605 717980
rect 40542 706213 40602 717979
rect 40726 707437 40786 718523
rect 41275 714236 41341 714237
rect 41275 714172 41276 714236
rect 41340 714172 41341 714236
rect 41275 714171 41341 714172
rect 41278 712197 41338 714171
rect 41275 712196 41341 712197
rect 41275 712132 41276 712196
rect 41340 712132 41341 712196
rect 41275 712131 41341 712132
rect 40723 707436 40789 707437
rect 40723 707372 40724 707436
rect 40788 707372 40789 707436
rect 40723 707371 40789 707372
rect 40539 706212 40605 706213
rect 40539 706148 40540 706212
rect 40604 706148 40605 706212
rect 40539 706147 40605 706148
rect 41462 700501 41522 725190
rect 41643 718316 41709 718317
rect 41643 718252 41644 718316
rect 41708 718252 41709 718316
rect 41643 718251 41709 718252
rect 41646 701861 41706 718251
rect 41827 716140 41893 716141
rect 41827 716076 41828 716140
rect 41892 716076 41893 716140
rect 41827 716075 41893 716076
rect 41830 702133 41890 716075
rect 41827 702132 41893 702133
rect 41827 702068 41828 702132
rect 41892 702068 41893 702132
rect 41827 702067 41893 702068
rect 41643 701860 41709 701861
rect 41643 701796 41644 701860
rect 41708 701796 41709 701860
rect 41643 701795 41709 701796
rect 41459 700500 41525 700501
rect 41459 700436 41460 700500
rect 41524 700436 41525 700500
rect 41459 700435 41525 700436
rect 41827 683636 41893 683637
rect 41827 683572 41828 683636
rect 41892 683572 41893 683636
rect 41827 683571 41893 683572
rect 41830 683090 41890 683571
rect 41646 683030 41890 683090
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 41646 678990 41706 683030
rect 40723 678927 40789 678928
rect 41462 678930 41706 678990
rect 40355 670988 40421 670989
rect 40355 670924 40356 670988
rect 40420 670924 40421 670988
rect 40355 670923 40421 670924
rect 40358 665549 40418 670923
rect 40355 665548 40421 665549
rect 40355 665484 40356 665548
rect 40420 665484 40421 665548
rect 40355 665483 40421 665484
rect 40542 662693 40602 678927
rect 40726 664053 40786 678927
rect 40907 677754 40973 677755
rect 40907 677690 40908 677754
rect 40972 677690 40973 677754
rect 40907 677689 40973 677690
rect 40910 665277 40970 677689
rect 41091 673028 41157 673029
rect 41091 672964 41092 673028
rect 41156 672964 41157 673028
rect 41091 672963 41157 672964
rect 41094 669085 41154 672963
rect 41091 669084 41157 669085
rect 41091 669020 41092 669084
rect 41156 669020 41157 669084
rect 41091 669019 41157 669020
rect 40907 665276 40973 665277
rect 40907 665212 40908 665276
rect 40972 665212 40973 665276
rect 40907 665211 40973 665212
rect 40723 664052 40789 664053
rect 40723 663988 40724 664052
rect 40788 663988 40789 664052
rect 40723 663987 40789 663988
rect 40539 662692 40605 662693
rect 40539 662628 40540 662692
rect 40604 662628 40605 662692
rect 40539 662627 40605 662628
rect 41462 660925 41522 678930
rect 41827 678876 41893 678877
rect 41827 678812 41828 678876
rect 41892 678812 41893 678876
rect 41827 678811 41893 678812
rect 41830 678330 41890 678811
rect 41646 678270 41890 678330
rect 41459 660924 41525 660925
rect 41459 660860 41460 660924
rect 41524 660860 41525 660924
rect 41459 660859 41525 660860
rect 41646 658613 41706 678270
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 672691
rect 43299 671940 43365 671941
rect 43299 671876 43300 671940
rect 43364 671876 43365 671940
rect 43299 671875 43365 671876
rect 42195 667452 42261 667453
rect 42195 667388 42196 667452
rect 42260 667388 42261 667452
rect 42195 667387 42261 667388
rect 42198 666637 42258 667387
rect 43302 666909 43362 671875
rect 43299 666908 43365 666909
rect 43299 666844 43300 666908
rect 43364 666844 43365 666908
rect 43299 666843 43365 666844
rect 42195 666636 42261 666637
rect 42195 666572 42196 666636
rect 42260 666572 42261 666636
rect 42195 666571 42261 666572
rect 674422 662421 674482 738107
rect 674606 707573 674666 782443
rect 676078 726885 676138 786659
rect 676811 739804 676877 739805
rect 676811 739740 676812 739804
rect 676876 739740 676877 739804
rect 676811 739739 676877 739740
rect 676075 726884 676141 726885
rect 676075 726820 676076 726884
rect 676140 726820 676141 726884
rect 676075 726819 676141 726820
rect 674787 722260 674853 722261
rect 674787 722196 674788 722260
rect 674852 722196 674853 722260
rect 674787 722195 674853 722196
rect 674790 707970 674850 722195
rect 676075 721580 676141 721581
rect 676075 721516 676076 721580
rect 676140 721516 676141 721580
rect 676075 721515 676141 721516
rect 674790 707910 675954 707970
rect 674603 707572 674669 707573
rect 674603 707508 674604 707572
rect 674668 707508 674669 707572
rect 674603 707507 674669 707508
rect 674603 706348 674669 706349
rect 674603 706284 674604 706348
rect 674668 706284 674669 706348
rect 674603 706283 674669 706284
rect 674419 662420 674485 662421
rect 674419 662356 674420 662420
rect 674484 662356 674485 662420
rect 674419 662355 674485 662356
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 674235 649772 674301 649773
rect 674235 649708 674236 649772
rect 674300 649708 674301 649772
rect 674235 649707 674301 649708
rect 44219 642292 44285 642293
rect 44219 642228 44220 642292
rect 44284 642228 44285 642292
rect 44219 642227 44285 642228
rect 41643 640660 41709 640661
rect 41643 640596 41644 640660
rect 41708 640596 41709 640660
rect 41643 640595 41709 640596
rect 41459 639436 41525 639437
rect 41459 639372 41460 639436
rect 41524 639372 41525 639436
rect 41459 639371 41525 639372
rect 40539 637396 40605 637397
rect 40539 637332 40540 637396
rect 40604 637332 40605 637396
rect 40539 637331 40605 637332
rect 40542 616453 40602 637331
rect 40723 635356 40789 635357
rect 40723 635292 40724 635356
rect 40788 635292 40789 635356
rect 40723 635291 40789 635292
rect 40726 620941 40786 635291
rect 40907 634948 40973 634949
rect 40907 634884 40908 634948
rect 40972 634884 40973 634948
rect 40907 634883 40973 634884
rect 40910 623797 40970 634883
rect 40907 623796 40973 623797
rect 40907 623732 40908 623796
rect 40972 623732 40973 623796
rect 40907 623731 40973 623732
rect 40723 620940 40789 620941
rect 40723 620876 40724 620940
rect 40788 620876 40789 620940
rect 40723 620875 40789 620876
rect 40539 616452 40605 616453
rect 40539 616388 40540 616452
rect 40604 616388 40605 616452
rect 40539 616387 40605 616388
rect 41462 615229 41522 639371
rect 41646 615773 41706 640595
rect 42379 632908 42445 632909
rect 42379 632844 42380 632908
rect 42444 632844 42445 632908
rect 42379 632843 42445 632844
rect 41827 629916 41893 629917
rect 41827 629852 41828 629916
rect 41892 629852 41893 629916
rect 41827 629851 41893 629852
rect 41830 616181 41890 629851
rect 42195 625700 42261 625701
rect 42195 625636 42196 625700
rect 42260 625636 42261 625700
rect 42195 625635 42261 625636
rect 42198 619853 42258 625635
rect 42382 624613 42442 632843
rect 42379 624612 42445 624613
rect 42379 624548 42380 624612
rect 42444 624548 42445 624612
rect 42379 624547 42445 624548
rect 42195 619852 42261 619853
rect 42195 619788 42196 619852
rect 42260 619788 42261 619852
rect 42195 619787 42261 619788
rect 41827 616180 41893 616181
rect 41827 616116 41828 616180
rect 41892 616116 41893 616180
rect 41827 616115 41893 616116
rect 41643 615772 41709 615773
rect 41643 615708 41644 615772
rect 41708 615708 41709 615772
rect 41643 615707 41709 615708
rect 41459 615228 41525 615229
rect 41459 615164 41460 615228
rect 41524 615164 41525 615228
rect 41459 615163 41525 615164
rect 44222 599725 44282 642227
rect 44219 599724 44285 599725
rect 44219 599660 44220 599724
rect 44284 599660 44285 599724
rect 44219 599659 44285 599660
rect 43115 599316 43181 599317
rect 43115 599252 43116 599316
rect 43180 599252 43181 599316
rect 43115 599251 43181 599252
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 41827 594012 41893 594013
rect 41827 594010 41828 594012
rect 40542 593950 41828 594010
rect 40355 590918 40421 590919
rect 40355 590854 40356 590918
rect 40420 590854 40421 590918
rect 40355 590853 40421 590854
rect 40358 589661 40418 590853
rect 40355 589660 40421 589661
rect 40355 589596 40356 589660
rect 40420 589596 40421 589660
rect 40355 589595 40421 589596
rect 40355 585988 40421 585989
rect 40355 585924 40356 585988
rect 40420 585924 40421 585988
rect 40355 585923 40421 585924
rect 40358 580277 40418 585923
rect 40355 580276 40421 580277
rect 40355 580212 40356 580276
rect 40420 580212 40421 580276
rect 40355 580211 40421 580212
rect 40542 575653 40602 593950
rect 41827 593948 41828 593950
rect 41892 593948 41893 594012
rect 41827 593947 41893 593948
rect 42014 593330 42074 597211
rect 43118 597005 43178 599251
rect 43115 597004 43181 597005
rect 43115 596940 43116 597004
rect 43180 596940 43181 597004
rect 43115 596939 43181 596940
rect 42195 596460 42261 596461
rect 42195 596396 42196 596460
rect 42260 596396 42261 596460
rect 42195 596395 42261 596396
rect 41646 593270 42074 593330
rect 40723 592958 40789 592959
rect 40723 592894 40724 592958
rect 40788 592894 40789 592958
rect 40723 592893 40789 592894
rect 40539 575652 40605 575653
rect 40539 575588 40540 575652
rect 40604 575588 40605 575652
rect 40539 575587 40605 575588
rect 40726 574701 40786 592893
rect 40910 592590 41522 592650
rect 40910 577829 40970 592590
rect 41462 592143 41522 592590
rect 41459 592142 41525 592143
rect 41459 592078 41460 592142
rect 41524 592078 41525 592142
rect 41459 592077 41525 592078
rect 41646 587210 41706 593270
rect 42198 589290 42258 596395
rect 674238 592653 674298 649707
rect 674419 616180 674485 616181
rect 674419 616116 674420 616180
rect 674484 616116 674485 616180
rect 674419 616115 674485 616116
rect 674235 592652 674301 592653
rect 674235 592588 674236 592652
rect 674300 592588 674301 592652
rect 674235 592587 674301 592588
rect 41462 587150 41706 587210
rect 41830 589230 42258 589290
rect 40907 577828 40973 577829
rect 40907 577764 40908 577828
rect 40972 577764 40973 577828
rect 40907 577763 40973 577764
rect 40723 574700 40789 574701
rect 40723 574636 40724 574700
rect 40788 574636 40789 574700
rect 40723 574635 40789 574636
rect 41462 572797 41522 587150
rect 41830 586530 41890 589230
rect 42195 587620 42261 587621
rect 42195 587556 42196 587620
rect 42260 587556 42261 587620
rect 42195 587555 42261 587556
rect 41646 586470 41890 586530
rect 41459 572796 41525 572797
rect 41459 572732 41460 572796
rect 41524 572732 41525 572796
rect 41459 572731 41525 572732
rect 41646 571573 41706 586470
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41643 571572 41709 571573
rect 41643 571508 41644 571572
rect 41708 571508 41709 571572
rect 41643 571507 41709 571508
rect 41830 570213 41890 585107
rect 42198 581909 42258 587555
rect 42195 581908 42261 581909
rect 42195 581844 42196 581908
rect 42260 581844 42261 581908
rect 42195 581843 42261 581844
rect 671475 570756 671541 570757
rect 671475 570692 671476 570756
rect 671540 570692 671541 570756
rect 671475 570691 671541 570692
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 41091 558788 41157 558789
rect 41091 558724 41092 558788
rect 41156 558724 41157 558788
rect 41091 558723 41157 558724
rect 41094 557553 41154 558723
rect 41091 557552 41157 557553
rect 41091 557488 41092 557552
rect 41156 557488 41157 557552
rect 41091 557487 41157 557488
rect 41827 554028 41893 554029
rect 41827 553964 41828 554028
rect 41892 553964 41893 554028
rect 41827 553963 41893 553964
rect 41830 553410 41890 553963
rect 41462 553350 41890 553410
rect 40723 545732 40789 545733
rect 40723 545668 40724 545732
rect 40788 545668 40789 545732
rect 40723 545667 40789 545668
rect 40539 545460 40605 545461
rect 40539 545396 40540 545460
rect 40604 545396 40605 545460
rect 40539 545395 40605 545396
rect 40542 537437 40602 545395
rect 40539 537436 40605 537437
rect 40539 537372 40540 537436
rect 40604 537372 40605 537436
rect 40539 537371 40605 537372
rect 40726 537029 40786 545667
rect 40723 537028 40789 537029
rect 40723 536964 40724 537028
rect 40788 536964 40789 537028
rect 40723 536963 40789 536964
rect 41462 530773 41522 553350
rect 41827 552804 41893 552805
rect 41827 552740 41828 552804
rect 41892 552740 41893 552804
rect 41827 552739 41893 552740
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 41459 530772 41525 530773
rect 41459 530708 41460 530772
rect 41524 530708 41525 530772
rect 41459 530707 41525 530708
rect 41646 529549 41706 546347
rect 41643 529548 41709 529549
rect 41643 529484 41644 529548
rect 41708 529484 41709 529548
rect 41643 529483 41709 529484
rect 41830 529005 41890 552739
rect 41827 529004 41893 529005
rect 41827 528940 41828 529004
rect 41892 528940 41893 529004
rect 41827 528939 41893 528940
rect 671478 474877 671538 570691
rect 673867 565588 673933 565589
rect 673867 565524 673868 565588
rect 673932 565524 673933 565588
rect 673867 565523 673933 565524
rect 673683 475420 673749 475421
rect 673683 475356 673684 475420
rect 673748 475356 673749 475420
rect 673683 475355 673749 475356
rect 671475 474876 671541 474877
rect 671475 474812 671476 474876
rect 671540 474812 671541 474876
rect 671475 474811 671541 474812
rect 673686 464813 673746 475355
rect 673683 464812 673749 464813
rect 673683 464748 673684 464812
rect 673748 464748 673749 464812
rect 673683 464747 673749 464748
rect 673870 455021 673930 565523
rect 674422 475421 674482 616115
rect 674606 477461 674666 706283
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 675342 687173 675402 696763
rect 675339 687172 675405 687173
rect 675339 687108 675340 687172
rect 675404 687108 675405 687172
rect 675339 687107 675405 687108
rect 675894 682141 675954 707910
rect 675891 682140 675957 682141
rect 675891 682076 675892 682140
rect 675956 682076 675957 682140
rect 675891 682075 675957 682076
rect 676078 681869 676138 721515
rect 676075 681868 676141 681869
rect 676075 681804 676076 681868
rect 676140 681804 676141 681868
rect 676075 681803 676141 681804
rect 676075 676428 676141 676429
rect 676075 676364 676076 676428
rect 676140 676364 676141 676428
rect 676075 676363 676141 676364
rect 674787 644060 674853 644061
rect 674787 643996 674788 644060
rect 674852 643996 674853 644060
rect 674787 643995 674853 643996
rect 674790 640253 674850 643995
rect 674787 640252 674853 640253
rect 674787 640188 674788 640252
rect 674852 640188 674853 640252
rect 674787 640187 674853 640188
rect 676078 636173 676138 676363
rect 676814 664189 676874 739739
rect 676995 686220 677061 686221
rect 676995 686156 676996 686220
rect 677060 686156 677061 686220
rect 676995 686155 677061 686156
rect 676811 664188 676877 664189
rect 676811 664124 676812 664188
rect 676876 664124 676877 664188
rect 676811 664123 676877 664124
rect 676811 648684 676877 648685
rect 676811 648620 676812 648684
rect 676876 648620 676877 648684
rect 676811 648619 676877 648620
rect 676075 636172 676141 636173
rect 676075 636108 676076 636172
rect 676140 636108 676141 636172
rect 676075 636107 676141 636108
rect 675339 608292 675405 608293
rect 675339 608228 675340 608292
rect 675404 608228 675405 608292
rect 675339 608227 675405 608228
rect 675342 592650 675402 608227
rect 675523 604620 675589 604621
rect 675523 604556 675524 604620
rect 675588 604556 675589 604620
rect 675523 604555 675589 604556
rect 675526 596325 675586 604555
rect 675523 596324 675589 596325
rect 675523 596260 675524 596324
rect 675588 596260 675589 596324
rect 675523 596259 675589 596260
rect 675342 592590 675586 592650
rect 675526 592109 675586 592590
rect 675523 592108 675589 592109
rect 675523 592044 675524 592108
rect 675588 592044 675589 592108
rect 675523 592043 675589 592044
rect 675155 586260 675221 586261
rect 675155 586196 675156 586260
rect 675220 586196 675221 586260
rect 675155 586195 675221 586196
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675158 576870 675218 586195
rect 675158 576810 675954 576870
rect 675339 561916 675405 561917
rect 675339 561852 675340 561916
rect 675404 561852 675405 561916
rect 675339 561851 675405 561852
rect 675342 544509 675402 561851
rect 675894 547365 675954 576810
rect 675891 547364 675957 547365
rect 675891 547300 675892 547364
rect 675956 547300 675957 547364
rect 675891 547299 675957 547300
rect 676078 547093 676138 586195
rect 676814 573613 676874 648619
rect 676998 621621 677058 686155
rect 676995 621620 677061 621621
rect 676995 621556 676996 621620
rect 677060 621556 677061 621620
rect 676995 621555 677061 621556
rect 676995 598908 677061 598909
rect 676995 598844 676996 598908
rect 677060 598844 677061 598908
rect 676995 598843 677061 598844
rect 676998 575245 677058 598843
rect 676995 575244 677061 575245
rect 676995 575180 676996 575244
rect 677060 575180 677061 575244
rect 676995 575179 677061 575180
rect 676811 573612 676877 573613
rect 676811 573548 676812 573612
rect 676876 573548 676877 573612
rect 676811 573547 676877 573548
rect 676443 562732 676509 562733
rect 676443 562668 676444 562732
rect 676508 562668 676509 562732
rect 676443 562667 676509 562668
rect 676446 547637 676506 562667
rect 676811 553892 676877 553893
rect 676811 553828 676812 553892
rect 676876 553828 676877 553892
rect 676811 553827 676877 553828
rect 676443 547636 676509 547637
rect 676443 547572 676444 547636
rect 676508 547572 676509 547636
rect 676443 547571 676509 547572
rect 676075 547092 676141 547093
rect 676075 547028 676076 547092
rect 676140 547028 676141 547092
rect 676075 547027 676141 547028
rect 675339 544508 675405 544509
rect 675339 544444 675340 544508
rect 675404 544444 675405 544508
rect 675339 544443 675405 544444
rect 676814 489290 676874 553827
rect 676995 552124 677061 552125
rect 676995 552060 676996 552124
rect 677060 552060 677061 552124
rect 676995 552059 677061 552060
rect 675526 489230 676874 489290
rect 675526 483581 675586 489230
rect 675707 488884 675773 488885
rect 675707 488820 675708 488884
rect 675772 488820 675773 488884
rect 675707 488819 675773 488820
rect 675523 483580 675589 483581
rect 675523 483516 675524 483580
rect 675588 483516 675589 483580
rect 675523 483515 675589 483516
rect 675710 481650 675770 488819
rect 676998 487930 677058 552059
rect 675894 487870 677058 487930
rect 675894 483989 675954 487870
rect 675891 483988 675957 483989
rect 675891 483924 675892 483988
rect 675956 483924 675957 483988
rect 675891 483923 675957 483924
rect 675710 481590 677242 481650
rect 674603 477460 674669 477461
rect 674603 477396 674604 477460
rect 674668 477396 674669 477460
rect 674603 477395 674669 477396
rect 674419 475420 674485 475421
rect 674419 475356 674420 475420
rect 674484 475356 674485 475420
rect 674419 475355 674485 475356
rect 673867 455020 673933 455021
rect 673867 454956 673868 455020
rect 673932 454956 673933 455020
rect 673867 454955 673933 454956
rect 675339 447812 675405 447813
rect 675339 447748 675340 447812
rect 675404 447748 675405 447812
rect 675339 447747 675405 447748
rect 41827 426460 41893 426461
rect 41827 426396 41828 426460
rect 41892 426396 41893 426460
rect 41827 426395 41893 426396
rect 41830 426050 41890 426395
rect 40542 425990 41890 426050
rect 40542 400077 40602 425990
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41827 422788 41893 422789
rect 41827 422724 41828 422788
rect 41892 422724 41893 422788
rect 41827 422723 41893 422724
rect 41830 422310 41890 422723
rect 40726 422250 41890 422310
rect 40726 409461 40786 422250
rect 41827 421972 41893 421973
rect 41827 421970 41828 421972
rect 40910 421910 41828 421970
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40910 405653 40970 421910
rect 41827 421908 41828 421910
rect 41892 421908 41893 421972
rect 41827 421907 41893 421908
rect 41459 418844 41525 418845
rect 41459 418780 41460 418844
rect 41524 418780 41525 418844
rect 41459 418779 41525 418780
rect 40907 405652 40973 405653
rect 40907 405588 40908 405652
rect 40972 405588 40973 405652
rect 40907 405587 40973 405588
rect 40539 400076 40605 400077
rect 40539 400012 40540 400076
rect 40604 400012 40605 400076
rect 40539 400011 40605 400012
rect 41462 398853 41522 418779
rect 41643 413404 41709 413405
rect 41643 413340 41644 413404
rect 41708 413340 41709 413404
rect 41643 413339 41709 413340
rect 41646 402990 41706 413339
rect 42014 408510 42074 424763
rect 42195 424284 42261 424285
rect 42195 424220 42196 424284
rect 42260 424220 42261 424284
rect 42195 424219 42261 424220
rect 42198 413405 42258 424219
rect 42195 413404 42261 413405
rect 42195 413340 42196 413404
rect 42260 413340 42261 413404
rect 42195 413339 42261 413340
rect 675342 410549 675402 447747
rect 676811 440332 676877 440333
rect 676811 440268 676812 440332
rect 676876 440268 676877 440332
rect 676811 440267 676877 440268
rect 675339 410548 675405 410549
rect 675339 410484 675340 410548
rect 675404 410484 675405 410548
rect 675339 410483 675405 410484
rect 41830 408450 42074 408510
rect 41830 406333 41890 408450
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41830 401845 41890 402930
rect 41827 401844 41893 401845
rect 41827 401780 41828 401844
rect 41892 401780 41893 401844
rect 41827 401779 41893 401780
rect 676814 400485 676874 440267
rect 677182 401301 677242 481590
rect 677179 401300 677245 401301
rect 677179 401236 677180 401300
rect 677244 401236 677245 401300
rect 677179 401235 677245 401236
rect 676811 400484 676877 400485
rect 676811 400420 676812 400484
rect 676876 400420 676877 400484
rect 676811 400419 676877 400420
rect 41459 398852 41525 398853
rect 41459 398788 41460 398852
rect 41524 398788 41525 398852
rect 41459 398787 41525 398788
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 389876 675957 389877
rect 675891 389812 675892 389876
rect 675956 389812 675957 389876
rect 675891 389811 675957 389812
rect 675707 388516 675773 388517
rect 675707 388452 675708 388516
rect 675772 388452 675773 388516
rect 675707 388451 675773 388452
rect 40539 380628 40605 380629
rect 40539 380564 40540 380628
rect 40604 380564 40605 380628
rect 40539 380563 40605 380564
rect 40542 356149 40602 380563
rect 41459 379812 41525 379813
rect 41459 379748 41460 379812
rect 41524 379748 41525 379812
rect 41459 379747 41525 379748
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363765 40786 378115
rect 41275 374644 41341 374645
rect 41275 374580 41276 374644
rect 41340 374580 41341 374644
rect 41275 374579 41341 374580
rect 41278 368525 41338 374579
rect 41275 368524 41341 368525
rect 41275 368460 41276 368524
rect 41340 368460 41341 368524
rect 41275 368459 41341 368460
rect 40723 363764 40789 363765
rect 40723 363700 40724 363764
rect 40788 363700 40789 363764
rect 40723 363699 40789 363700
rect 41462 358733 41522 379747
rect 675710 378725 675770 388451
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 675894 373013 675954 389811
rect 676078 373693 676138 398787
rect 676259 396812 676325 396813
rect 676259 396748 676260 396812
rect 676324 396748 676325 396812
rect 676259 396747 676325 396748
rect 676262 385389 676322 396747
rect 676443 395996 676509 395997
rect 676443 395932 676444 395996
rect 676508 395932 676509 395996
rect 676443 395931 676509 395932
rect 676259 385388 676325 385389
rect 676259 385324 676260 385388
rect 676324 385324 676325 385388
rect 676259 385323 676325 385324
rect 676446 381717 676506 395931
rect 676627 395180 676693 395181
rect 676627 395116 676628 395180
rect 676692 395116 676693 395180
rect 676627 395115 676693 395116
rect 676443 381716 676509 381717
rect 676443 381652 676444 381716
rect 676508 381652 676509 381716
rect 676443 381651 676509 381652
rect 676630 377365 676690 395115
rect 676627 377364 676693 377365
rect 676627 377300 676628 377364
rect 676692 377300 676693 377364
rect 676627 377299 676693 377300
rect 676075 373692 676141 373693
rect 676075 373628 676076 373692
rect 676140 373628 676141 373692
rect 676075 373627 676141 373628
rect 675891 373012 675957 373013
rect 675891 372948 675892 373012
rect 675956 372948 675957 373012
rect 675891 372947 675957 372948
rect 41643 372740 41709 372741
rect 41643 372676 41644 372740
rect 41708 372676 41709 372740
rect 41643 372675 41709 372676
rect 41646 359549 41706 372675
rect 41827 371924 41893 371925
rect 41827 371860 41828 371924
rect 41892 371860 41893 371924
rect 41827 371859 41893 371860
rect 41830 360093 41890 371859
rect 41827 360092 41893 360093
rect 41827 360028 41828 360092
rect 41892 360028 41893 360092
rect 41827 360027 41893 360028
rect 41643 359548 41709 359549
rect 41643 359484 41644 359548
rect 41708 359484 41709 359548
rect 41643 359483 41709 359484
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 40539 356148 40605 356149
rect 40539 356084 40540 356148
rect 40604 356084 40605 356148
rect 40539 356083 40605 356084
rect 675523 353428 675589 353429
rect 675523 353364 675524 353428
rect 675588 353364 675589 353428
rect 675523 353363 675589 353364
rect 44403 342956 44469 342957
rect 44403 342892 44404 342956
rect 44468 342892 44469 342956
rect 44403 342891 44469 342892
rect 44219 341596 44285 341597
rect 44219 341532 44220 341596
rect 44284 341532 44285 341596
rect 44219 341531 44285 341532
rect 42747 340508 42813 340509
rect 42747 340444 42748 340508
rect 42812 340444 42813 340508
rect 42747 340443 42813 340444
rect 41643 338196 41709 338197
rect 41643 338132 41644 338196
rect 41708 338132 41709 338196
rect 41643 338131 41709 338132
rect 40723 336972 40789 336973
rect 40723 336908 40724 336972
rect 40788 336908 40789 336972
rect 40723 336907 40789 336908
rect 40539 335340 40605 335341
rect 40539 335276 40540 335340
rect 40604 335276 40605 335340
rect 40539 335275 40605 335276
rect 40542 317389 40602 335275
rect 40726 319021 40786 336907
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40910 325413 40970 333643
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 41646 319970 41706 338131
rect 42011 336564 42077 336565
rect 42011 336500 42012 336564
rect 42076 336500 42077 336564
rect 42011 336499 42077 336500
rect 41827 335748 41893 335749
rect 41827 335684 41828 335748
rect 41892 335684 41893 335748
rect 41827 335683 41893 335684
rect 41830 324869 41890 335683
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41827 319972 41893 319973
rect 41827 319970 41828 319972
rect 41646 319910 41828 319970
rect 41827 319908 41828 319910
rect 41892 319908 41893 319972
rect 41827 319907 41893 319908
rect 40723 319020 40789 319021
rect 40723 318956 40724 319020
rect 40788 318956 40789 319020
rect 40723 318955 40789 318956
rect 40539 317388 40605 317389
rect 40539 317324 40540 317388
rect 40604 317324 40605 317388
rect 40539 317323 40605 317324
rect 42014 313717 42074 336499
rect 42011 313716 42077 313717
rect 42011 313652 42012 313716
rect 42076 313652 42077 313716
rect 42011 313651 42077 313652
rect 42750 297669 42810 340443
rect 42931 337652 42997 337653
rect 42931 337588 42932 337652
rect 42996 337588 42997 337652
rect 42931 337587 42997 337588
rect 42934 312765 42994 337587
rect 43115 337244 43181 337245
rect 43115 337180 43116 337244
rect 43180 337180 43181 337244
rect 43115 337179 43181 337180
rect 43118 316029 43178 337179
rect 43115 316028 43181 316029
rect 43115 315964 43116 316028
rect 43180 315964 43181 316028
rect 43115 315963 43181 315964
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 44222 298485 44282 341531
rect 44406 300117 44466 342891
rect 675526 340781 675586 353363
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 349210 675770 352955
rect 675937 352204 676003 352205
rect 675937 352140 675938 352204
rect 676002 352202 676003 352204
rect 676002 352142 676322 352202
rect 676002 352140 676003 352142
rect 675937 352139 676003 352140
rect 675891 351932 675957 351933
rect 675891 351868 675892 351932
rect 675956 351930 675957 351932
rect 675956 351870 676138 351930
rect 675956 351868 675957 351870
rect 675891 351867 675957 351868
rect 675710 349150 675954 349210
rect 675523 340780 675589 340781
rect 675523 340716 675524 340780
rect 675588 340716 675589 340780
rect 675523 340715 675589 340716
rect 44587 340236 44653 340237
rect 44587 340172 44588 340236
rect 44652 340172 44653 340236
rect 44587 340171 44653 340172
rect 44403 300116 44469 300117
rect 44403 300052 44404 300116
rect 44468 300052 44469 300116
rect 44403 300051 44469 300052
rect 44590 299301 44650 340171
rect 675894 337789 675954 349150
rect 675891 337788 675957 337789
rect 675891 337724 675892 337788
rect 675956 337724 675957 337788
rect 675891 337723 675957 337724
rect 676078 328405 676138 351870
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 676262 325549 676322 352142
rect 676443 346628 676509 346629
rect 676443 346564 676444 346628
rect 676508 346564 676509 346628
rect 676443 346563 676509 346564
rect 676446 340237 676506 346563
rect 676811 346220 676877 346221
rect 676811 346156 676812 346220
rect 676876 346156 676877 346220
rect 676811 346155 676877 346156
rect 676443 340236 676509 340237
rect 676443 340172 676444 340236
rect 676508 340172 676509 340236
rect 676443 340171 676509 340172
rect 676259 325548 676325 325549
rect 676259 325484 676260 325548
rect 676324 325484 676325 325548
rect 676259 325483 676325 325484
rect 676814 325277 676874 346155
rect 676811 325276 676877 325277
rect 676811 325212 676812 325276
rect 676876 325212 676877 325276
rect 676811 325211 676877 325212
rect 675707 309092 675773 309093
rect 675707 309028 675708 309092
rect 675772 309090 675773 309092
rect 675772 309030 675954 309090
rect 675772 309028 675773 309030
rect 675707 309027 675773 309028
rect 675707 308820 675773 308821
rect 675707 308756 675708 308820
rect 675772 308756 675773 308820
rect 675707 308755 675773 308756
rect 675710 302250 675770 308755
rect 675894 307730 675954 309030
rect 675894 307670 676690 307730
rect 675891 307188 675957 307189
rect 675891 307124 675892 307188
rect 675956 307124 675957 307188
rect 675891 307123 675957 307124
rect 675894 303650 675954 307123
rect 675894 303590 676138 303650
rect 675710 302190 675954 302250
rect 675707 299436 675773 299437
rect 675707 299372 675708 299436
rect 675772 299372 675773 299436
rect 675707 299371 675773 299372
rect 44587 299300 44653 299301
rect 44587 299236 44588 299300
rect 44652 299236 44653 299300
rect 44587 299235 44653 299236
rect 44219 298484 44285 298485
rect 44219 298420 44220 298484
rect 44284 298420 44285 298484
rect 44219 298419 44285 298420
rect 42747 297668 42813 297669
rect 42747 297604 42748 297668
rect 42812 297604 42813 297668
rect 42747 297603 42813 297604
rect 42011 296852 42077 296853
rect 42011 296788 42012 296852
rect 42076 296788 42077 296852
rect 42011 296787 42077 296788
rect 675339 296852 675405 296853
rect 675339 296788 675340 296852
rect 675404 296788 675405 296852
rect 675339 296787 675405 296788
rect 41367 292592 41433 292593
rect 41367 292528 41368 292592
rect 41432 292528 41433 292592
rect 41367 292527 41433 292528
rect 41370 292090 41430 292527
rect 40542 292030 41430 292090
rect 40542 274277 40602 292030
rect 41827 291548 41893 291549
rect 41827 291484 41828 291548
rect 41892 291484 41893 291548
rect 41827 291483 41893 291484
rect 41830 289830 41890 291483
rect 40910 289770 41890 289830
rect 40723 289236 40789 289237
rect 40723 289172 40724 289236
rect 40788 289172 40789 289236
rect 40723 289171 40789 289172
rect 40726 277133 40786 289171
rect 40910 278493 40970 289770
rect 42014 288010 42074 296787
rect 675342 295357 675402 296787
rect 675523 296580 675589 296581
rect 675523 296516 675524 296580
rect 675588 296516 675589 296580
rect 675523 296515 675589 296516
rect 675339 295356 675405 295357
rect 675339 295292 675340 295356
rect 675404 295292 675405 295356
rect 675339 295291 675405 295292
rect 675526 292229 675586 296515
rect 675523 292228 675589 292229
rect 675523 292164 675524 292228
rect 675588 292164 675589 292228
rect 675523 292163 675589 292164
rect 41462 287950 42074 288010
rect 40907 278492 40973 278493
rect 40907 278428 40908 278492
rect 40972 278428 40973 278492
rect 40907 278427 40973 278428
rect 40723 277132 40789 277133
rect 40723 277068 40724 277132
rect 40788 277068 40789 277132
rect 40723 277067 40789 277068
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 287950
rect 41643 284884 41709 284885
rect 41643 284820 41644 284884
rect 41708 284820 41709 284884
rect 41643 284819 41709 284820
rect 41646 282930 41706 284819
rect 42011 284340 42077 284341
rect 42011 284276 42012 284340
rect 42076 284276 42077 284340
rect 42011 284275 42077 284276
rect 41646 282870 41890 282930
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 270061 41890 282870
rect 42014 272373 42074 284275
rect 675710 282845 675770 299371
rect 675894 283661 675954 302190
rect 675891 283660 675957 283661
rect 675891 283596 675892 283660
rect 675956 283596 675957 283660
rect 675891 283595 675957 283596
rect 675707 282844 675773 282845
rect 675707 282780 675708 282844
rect 675772 282780 675773 282844
rect 675707 282779 675773 282780
rect 676078 281213 676138 303590
rect 676443 301612 676509 301613
rect 676443 301548 676444 301612
rect 676508 301548 676509 301612
rect 676443 301547 676509 301548
rect 676259 300660 676325 300661
rect 676259 300596 676260 300660
rect 676324 300596 676325 300660
rect 676259 300595 676325 300596
rect 676262 290869 676322 300595
rect 676446 291549 676506 301547
rect 676630 294541 676690 307670
rect 676627 294540 676693 294541
rect 676627 294476 676628 294540
rect 676692 294476 676693 294540
rect 676627 294475 676693 294476
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676259 290868 676325 290869
rect 676259 290804 676260 290868
rect 676324 290804 676325 290868
rect 676259 290803 676325 290804
rect 676075 281212 676141 281213
rect 676075 281148 676076 281212
rect 676140 281148 676141 281212
rect 676075 281147 676141 281148
rect 42011 272372 42077 272373
rect 42011 272308 42012 272372
rect 42076 272308 42077 272372
rect 42011 272307 42077 272308
rect 41827 270060 41893 270061
rect 41827 269996 41828 270060
rect 41892 269996 41893 270060
rect 41827 269995 41893 269996
rect 674971 264212 675037 264213
rect 674971 264148 674972 264212
rect 675036 264148 675037 264212
rect 674971 264147 675037 264148
rect 40539 250204 40605 250205
rect 40539 250140 40540 250204
rect 40604 250140 40605 250204
rect 40539 250139 40605 250140
rect 40542 233069 40602 250139
rect 674974 249797 675034 264147
rect 676075 263668 676141 263669
rect 676075 263604 676076 263668
rect 676140 263604 676141 263668
rect 676075 263603 676141 263604
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 674971 249796 675037 249797
rect 674971 249732 674972 249796
rect 675036 249732 675037 249796
rect 674971 249731 675037 249732
rect 40726 236605 40786 249731
rect 676078 249661 676138 263603
rect 676811 261628 676877 261629
rect 676811 261564 676812 261628
rect 676876 261564 676877 261628
rect 676811 261563 676877 261564
rect 676814 250205 676874 261563
rect 676995 259996 677061 259997
rect 676995 259932 676996 259996
rect 677060 259932 677061 259996
rect 676995 259931 677061 259932
rect 676811 250204 676877 250205
rect 676811 250140 676812 250204
rect 676876 250140 676877 250204
rect 676811 250139 676877 250140
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 673315 246260 673381 246261
rect 673315 246196 673316 246260
rect 673380 246196 673381 246260
rect 673315 246195 673381 246196
rect 42011 237420 42077 237421
rect 42011 237356 42012 237420
rect 42076 237356 42077 237420
rect 42011 237355 42077 237356
rect 40723 236604 40789 236605
rect 40723 236540 40724 236604
rect 40788 236540 40789 236604
rect 40723 236539 40789 236540
rect 40539 233068 40605 233069
rect 40539 233004 40540 233068
rect 40604 233004 40605 233068
rect 40539 233003 40605 233004
rect 42014 228989 42074 237355
rect 42011 228988 42077 228989
rect 42011 228924 42012 228988
rect 42076 228924 42077 228988
rect 42011 228923 42077 228924
rect 671107 224772 671173 224773
rect 671107 224708 671108 224772
rect 671172 224708 671173 224772
rect 671107 224707 671173 224708
rect 671110 223141 671170 224707
rect 671107 223140 671173 223141
rect 671107 223076 671108 223140
rect 671172 223076 671173 223140
rect 671107 223075 671173 223076
rect 509187 217836 509253 217837
rect 509187 217772 509188 217836
rect 509252 217772 509253 217836
rect 522619 217836 522685 217837
rect 509187 217771 509253 217772
rect 510107 217772 510108 217822
rect 510172 217772 510173 217822
rect 510107 217771 510173 217772
rect 522619 217772 522620 217836
rect 522684 217772 522685 217836
rect 522619 217771 522685 217772
rect 566963 217836 567029 217837
rect 566963 217772 566964 217836
rect 567028 217772 567029 217836
rect 566963 217771 567029 217772
rect 574323 217772 574324 217822
rect 574388 217772 574389 217822
rect 574323 217771 574389 217772
rect 509190 215933 509250 217771
rect 509187 215932 509253 215933
rect 509187 215868 509188 215932
rect 509252 215868 509253 215932
rect 509187 215867 509253 215868
rect 522622 215389 522682 217771
rect 566966 216205 567026 217771
rect 574326 216749 574386 217142
rect 574323 216748 574389 216749
rect 574323 216684 574324 216748
rect 574388 216684 574389 216748
rect 574323 216683 574389 216684
rect 566963 216204 567029 216205
rect 566963 216140 566964 216204
rect 567028 216140 567029 216204
rect 566963 216139 567029 216140
rect 522619 215388 522685 215389
rect 522619 215324 522620 215388
rect 522684 215324 522685 215388
rect 522619 215323 522685 215324
rect 670739 210492 670805 210493
rect 670739 210428 670740 210492
rect 670804 210428 670805 210492
rect 670739 210427 670805 210428
rect 41827 210084 41893 210085
rect 41827 210020 41828 210084
rect 41892 210020 41893 210084
rect 41827 210019 41893 210020
rect 41459 208180 41525 208181
rect 41459 208116 41460 208180
rect 41524 208116 41525 208180
rect 41459 208115 41525 208116
rect 40539 207364 40605 207365
rect 40539 207300 40540 207364
rect 40604 207300 40605 207364
rect 40539 207299 40605 207300
rect 40542 186421 40602 207299
rect 40723 206548 40789 206549
rect 40723 206484 40724 206548
rect 40788 206484 40789 206548
rect 40723 206483 40789 206484
rect 40726 193221 40786 206483
rect 40907 206140 40973 206141
rect 40907 206076 40908 206140
rect 40972 206076 40973 206140
rect 40907 206075 40973 206076
rect 40910 194989 40970 206075
rect 40907 194988 40973 194989
rect 40907 194924 40908 194988
rect 40972 194924 40973 194988
rect 40907 194923 40973 194924
rect 40723 193220 40789 193221
rect 40723 193156 40724 193220
rect 40788 193156 40789 193220
rect 40723 193155 40789 193156
rect 40539 186420 40605 186421
rect 40539 186356 40540 186420
rect 40604 186356 40605 186420
rect 40539 186355 40605 186356
rect 41462 186013 41522 208115
rect 41643 205732 41709 205733
rect 41643 205668 41644 205732
rect 41708 205668 41709 205732
rect 41643 205667 41709 205668
rect 41646 190470 41706 205667
rect 41830 195261 41890 210019
rect 41827 195260 41893 195261
rect 41827 195196 41828 195260
rect 41892 195196 41893 195260
rect 41827 195195 41893 195196
rect 41646 190410 41890 190470
rect 41459 186012 41525 186013
rect 41459 185948 41460 186012
rect 41524 185948 41525 186012
rect 41459 185947 41525 185948
rect 41830 184109 41890 190410
rect 41827 184108 41893 184109
rect 41827 184044 41828 184108
rect 41892 184044 41893 184108
rect 41827 184043 41893 184044
rect 669451 171052 669517 171053
rect 669451 170988 669452 171052
rect 669516 170988 669517 171052
rect 669451 170987 669517 170988
rect 669454 157350 669514 170987
rect 669270 157290 669514 157350
rect 669270 140453 669330 157290
rect 669267 140452 669333 140453
rect 669267 140388 669268 140452
rect 669332 140388 669333 140452
rect 669267 140387 669333 140388
rect 670742 125765 670802 210427
rect 673318 161397 673378 246195
rect 676998 242317 677058 259931
rect 676995 242316 677061 242317
rect 676995 242252 676996 242316
rect 677060 242252 677061 242316
rect 676995 242251 677061 242252
rect 676811 241908 676877 241909
rect 676811 241844 676812 241908
rect 676876 241844 676877 241908
rect 676811 241843 676877 241844
rect 674971 241636 675037 241637
rect 674971 241572 674972 241636
rect 675036 241572 675037 241636
rect 674971 241571 675037 241572
rect 674974 230213 675034 241571
rect 674971 230212 675037 230213
rect 674971 230148 674972 230212
rect 675036 230148 675037 230212
rect 674971 230147 675037 230148
rect 674051 229804 674117 229805
rect 674051 229740 674052 229804
rect 674116 229740 674117 229804
rect 674051 229739 674117 229740
rect 673683 215252 673749 215253
rect 673683 215188 673684 215252
rect 673748 215188 673749 215252
rect 673683 215187 673749 215188
rect 673686 212550 673746 215187
rect 673502 212490 673746 212550
rect 673315 161396 673381 161397
rect 673315 161332 673316 161396
rect 673380 161332 673381 161396
rect 673315 161331 673381 161332
rect 673502 132701 673562 212490
rect 674054 132973 674114 229739
rect 674235 221916 674301 221917
rect 674235 221852 674236 221916
rect 674300 221852 674301 221916
rect 674235 221851 674301 221852
rect 674238 212805 674298 221851
rect 675891 220692 675957 220693
rect 675891 220628 675892 220692
rect 675956 220690 675957 220692
rect 676814 220690 676874 241843
rect 675956 220630 676874 220690
rect 675956 220628 675957 220630
rect 675891 220627 675957 220628
rect 675891 218244 675957 218245
rect 675891 218180 675892 218244
rect 675956 218180 675957 218244
rect 675891 218179 675957 218180
rect 675894 217970 675954 218179
rect 675894 217910 676506 217970
rect 675707 217428 675773 217429
rect 675707 217364 675708 217428
rect 675772 217364 675773 217428
rect 675707 217363 675773 217364
rect 674235 212804 674301 212805
rect 674235 212740 674236 212804
rect 674300 212740 674301 212804
rect 674235 212739 674301 212740
rect 675710 198389 675770 217363
rect 675891 215252 675957 215253
rect 675891 215188 675892 215252
rect 675956 215250 675957 215252
rect 675956 215190 676322 215250
rect 675956 215188 675957 215190
rect 675891 215187 675957 215188
rect 675891 214436 675957 214437
rect 675891 214372 675892 214436
rect 675956 214372 675957 214436
rect 675891 214371 675957 214372
rect 675894 211170 675954 214371
rect 675894 211110 676138 211170
rect 675891 210628 675957 210629
rect 675891 210564 675892 210628
rect 675956 210564 675957 210628
rect 675891 210563 675957 210564
rect 675707 198388 675773 198389
rect 675707 198324 675708 198388
rect 675772 198324 675773 198388
rect 675707 198323 675773 198324
rect 675894 192677 675954 210563
rect 676078 210490 676138 211110
rect 676262 210901 676322 215190
rect 676259 210900 676325 210901
rect 676259 210836 676260 210900
rect 676324 210836 676325 210900
rect 676259 210835 676325 210836
rect 676078 210430 676322 210490
rect 676075 206956 676141 206957
rect 676075 206892 676076 206956
rect 676140 206892 676141 206956
rect 676075 206891 676141 206892
rect 676078 204237 676138 206891
rect 676075 204236 676141 204237
rect 676075 204172 676076 204236
rect 676140 204172 676141 204236
rect 676075 204171 676141 204172
rect 676262 200701 676322 210430
rect 676446 205597 676506 217910
rect 676627 210900 676693 210901
rect 676627 210836 676628 210900
rect 676692 210836 676693 210900
rect 676627 210835 676693 210836
rect 676443 205596 676509 205597
rect 676443 205532 676444 205596
rect 676508 205532 676509 205596
rect 676443 205531 676509 205532
rect 676259 200700 676325 200701
rect 676259 200636 676260 200700
rect 676324 200636 676325 200700
rect 676259 200635 676325 200636
rect 676630 196077 676690 210835
rect 676627 196076 676693 196077
rect 676627 196012 676628 196076
rect 676692 196012 676693 196076
rect 676627 196011 676693 196012
rect 675891 192676 675957 192677
rect 675891 192612 675892 192676
rect 675956 192612 675957 192676
rect 675891 192611 675957 192612
rect 675523 173636 675589 173637
rect 675523 173572 675524 173636
rect 675588 173572 675589 173636
rect 675523 173571 675589 173572
rect 675526 162213 675586 173571
rect 675891 172820 675957 172821
rect 675891 172756 675892 172820
rect 675956 172756 675957 172820
rect 675891 172755 675957 172756
rect 675707 172412 675773 172413
rect 675707 172348 675708 172412
rect 675772 172348 675773 172412
rect 675894 172410 675954 172755
rect 675894 172350 676506 172410
rect 675707 172347 675773 172348
rect 675710 169010 675770 172347
rect 675891 169692 675957 169693
rect 675891 169628 675892 169692
rect 675956 169690 675957 169692
rect 675956 169630 676322 169690
rect 675956 169628 675957 169630
rect 675891 169627 675957 169628
rect 675710 168950 675954 169010
rect 675707 167516 675773 167517
rect 675707 167452 675708 167516
rect 675772 167452 675773 167516
rect 675707 167451 675773 167452
rect 675523 162212 675589 162213
rect 675523 162148 675524 162212
rect 675588 162148 675589 162212
rect 675523 162147 675589 162148
rect 675710 147661 675770 167451
rect 675894 153101 675954 168950
rect 676075 162212 676141 162213
rect 676075 162148 676076 162212
rect 676140 162148 676141 162212
rect 676075 162147 676141 162148
rect 675891 153100 675957 153101
rect 675891 153036 675892 153100
rect 675956 153036 675957 153100
rect 675891 153035 675957 153036
rect 676078 148477 676138 162147
rect 676262 155685 676322 169630
rect 676446 157045 676506 172350
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 157044 676509 157045
rect 676443 156980 676444 157044
rect 676508 156980 676509 157044
rect 676443 156979 676509 156980
rect 676259 155684 676325 155685
rect 676259 155620 676260 155684
rect 676324 155620 676325 155684
rect 676259 155619 676325 155620
rect 676630 151469 676690 166363
rect 676627 151468 676693 151469
rect 676627 151404 676628 151468
rect 676692 151404 676693 151468
rect 676627 151403 676693 151404
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675707 147660 675773 147661
rect 675707 147596 675708 147660
rect 675772 147596 675773 147660
rect 675707 147595 675773 147596
rect 674051 132972 674117 132973
rect 674051 132908 674052 132972
rect 674116 132908 674117 132972
rect 674051 132907 674117 132908
rect 673499 132700 673565 132701
rect 673499 132636 673500 132700
rect 673564 132636 673565 132700
rect 673499 132635 673565 132636
rect 676443 127396 676509 127397
rect 676443 127332 676444 127396
rect 676508 127332 676509 127396
rect 676443 127331 676509 127332
rect 675891 127260 675957 127261
rect 675891 127196 675892 127260
rect 675956 127196 675957 127260
rect 675891 127195 675957 127196
rect 670739 125764 670805 125765
rect 670739 125700 670740 125764
rect 670804 125700 670805 125764
rect 670739 125699 670805 125700
rect 675707 116108 675773 116109
rect 675707 116044 675708 116108
rect 675772 116044 675773 116108
rect 675707 116043 675773 116044
rect 675710 102645 675770 116043
rect 675894 108085 675954 127195
rect 676075 126172 676141 126173
rect 676075 126108 676076 126172
rect 676140 126108 676141 126172
rect 676075 126107 676141 126108
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 676078 103189 676138 126107
rect 676259 124540 676325 124541
rect 676259 124476 676260 124540
rect 676324 124476 676325 124540
rect 676259 124475 676325 124476
rect 676262 110397 676322 124475
rect 676446 112437 676506 127331
rect 676811 122908 676877 122909
rect 676811 122844 676812 122908
rect 676876 122844 676877 122908
rect 676811 122843 676877 122844
rect 676814 114341 676874 122843
rect 676811 114340 676877 114341
rect 676811 114276 676812 114340
rect 676876 114276 676877 114340
rect 676811 114275 676877 114276
rect 676443 112436 676509 112437
rect 676443 112372 676444 112436
rect 676508 112372 676509 112436
rect 676443 112371 676509 112372
rect 676259 110396 676325 110397
rect 676259 110332 676260 110396
rect 676324 110332 676325 110396
rect 676259 110331 676325 110332
rect 676075 103188 676141 103189
rect 676075 103124 676076 103188
rect 676140 103124 676141 103188
rect 676075 103123 676141 103124
rect 675707 102644 675773 102645
rect 675707 102580 675708 102644
rect 675772 102580 675773 102644
rect 675707 102579 675773 102580
rect 635779 96932 635845 96933
rect 635779 96868 635780 96932
rect 635844 96868 635845 96932
rect 635779 96867 635845 96868
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 95980 634005 95981
rect 633939 95916 633940 95980
rect 634004 95916 634005 95980
rect 633939 95915 634005 95916
rect 633942 78573 634002 95915
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 635782 78165 635842 96867
rect 637254 84210 637314 96867
rect 647187 96524 647253 96525
rect 647187 96460 647188 96524
rect 647252 96460 647253 96524
rect 647187 96459 647253 96460
rect 647190 94298 647250 96459
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 635779 78164 635845 78165
rect 635779 78100 635780 78164
rect 635844 78100 635845 78164
rect 635779 78099 635845 78100
rect 637070 77621 637130 84150
rect 637067 77620 637133 77621
rect 637067 77556 637068 77620
rect 637132 77556 637133 77620
rect 637067 77555 637133 77556
rect 461715 55044 461781 55045
rect 461715 54980 461716 55044
rect 461780 54980 461781 55044
rect 461715 54979 461781 54980
rect 461718 53957 461778 54979
rect 461715 53956 461781 53957
rect 461715 53892 461716 53956
rect 461780 53892 461781 53956
rect 461715 53891 461781 53892
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40357 141802 43963
rect 194366 42125 194426 50219
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 463923 44572 463989 44573
rect 463923 44508 463924 44572
rect 463988 44508 463989 44572
rect 463923 44507 463989 44508
rect 463739 44436 463805 44437
rect 463739 44372 463740 44436
rect 463804 44372 463805 44436
rect 463739 44371 463805 44372
rect 416635 42396 416701 42397
rect 416635 42332 416636 42396
rect 416700 42332 416701 42396
rect 416635 42331 416701 42332
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 365667 41852 365733 41853
rect 365667 41788 365668 41852
rect 365732 41788 365733 41852
rect 365667 41787 365733 41788
rect 365670 41258 365730 41787
rect 416638 40493 416698 42331
rect 460979 42124 461045 42125
rect 460979 42060 460980 42124
rect 461044 42060 461045 42124
rect 460979 42059 461045 42060
rect 421971 41852 422037 41853
rect 421971 41788 421972 41852
rect 422036 41850 422037 41852
rect 422036 41790 422162 41850
rect 422036 41788 422037 41790
rect 421971 41787 422037 41788
rect 460611 41852 460677 41853
rect 460611 41788 460612 41852
rect 460676 41850 460677 41852
rect 460982 41850 461042 42059
rect 463742 41938 463802 44371
rect 463926 42125 463986 44507
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 463923 42124 463989 42125
rect 463923 42060 463924 42124
rect 463988 42060 463989 42124
rect 463923 42059 463989 42060
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 460676 41790 461042 41850
rect 460676 41788 460677 41790
rect 460611 41787 460677 41788
rect 416635 40492 416701 40493
rect 416635 40428 416636 40492
rect 416700 40428 416701 40492
rect 416635 40427 416701 40428
rect 141739 40356 141805 40357
rect 141739 40292 141740 40356
rect 141804 40292 141805 40356
rect 141739 40291 141805 40292
<< via4 >>
rect 510022 217836 510258 218058
rect 510022 217822 510108 217836
rect 510108 217822 510172 217836
rect 510172 217822 510258 217836
rect 574238 217836 574474 218058
rect 574238 217822 574324 217836
rect 574324 217822 574388 217836
rect 574388 217822 574474 217836
rect 493646 217292 493882 217378
rect 493646 217228 493732 217292
rect 493732 217228 493796 217292
rect 493796 217228 493882 217292
rect 493646 217142 493882 217228
rect 574238 217142 574474 217378
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 361902 41852 362138 41938
rect 361902 41788 361988 41852
rect 361988 41788 362052 41852
rect 362052 41788 362138 41852
rect 361902 41702 362138 41788
rect 402750 41852 402986 41938
rect 402750 41788 402836 41852
rect 402836 41788 402900 41852
rect 402900 41788 402986 41852
rect 402750 41702 402986 41788
rect 365582 41022 365818 41258
rect 422162 41702 422398 41938
rect 451142 41852 451378 41938
rect 451142 41788 451228 41852
rect 451228 41788 451292 41852
rect 451292 41788 451378 41852
rect 451142 41702 451378 41788
rect 463654 41702 463890 41938
<< metal5 >>
rect 78610 1018624 90778 1030789
rect 130010 1018624 142178 1030789
rect 181410 1018624 193578 1030789
rect 231810 1018624 243978 1030789
rect 284410 1018624 296578 1030789
rect 334810 1018624 346978 1030789
rect 386210 1018624 398378 1030789
rect 475210 1018624 487378 1030789
rect 526610 1018624 538778 1030789
rect 577010 1018624 589178 1030789
rect 628410 1018624 640578 1030789
rect 6811 956610 18976 968778
rect 698624 953022 710789 965190
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 509980 218058 574516 218100
rect 509980 217822 510022 218058
rect 510258 217822 574238 218058
rect 574474 217822 574516 218058
rect 509980 217780 574516 217822
rect 493604 217378 574516 217420
rect 493604 217142 493646 217378
rect 493882 217142 574238 217378
rect 574474 217142 574516 217378
rect 493604 217100 574516 217142
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 361860 41938 403028 41980
rect 361860 41702 361902 41938
rect 362138 41702 402750 41938
rect 402986 41702 403028 41938
rect 361860 41660 403028 41702
rect 403444 41660 412044 41980
rect 403444 41300 403764 41660
rect 365540 41258 403764 41300
rect 365540 41022 365582 41258
rect 365818 41022 403764 41258
rect 365540 40980 403764 41022
rect 411724 41300 412044 41660
rect 412460 41660 421796 41980
rect 422120 41938 451420 41980
rect 422120 41702 422162 41938
rect 422398 41702 451142 41938
rect 451378 41702 451420 41938
rect 422120 41660 451420 41702
rect 451836 41660 461080 41980
rect 412460 41300 412780 41660
rect 411724 40980 412780 41300
rect 421476 41300 421796 41660
rect 451836 41300 452156 41660
rect 421476 40980 452156 41300
rect 460760 41300 461080 41660
rect 461404 41938 463932 41980
rect 461404 41702 463654 41938
rect 463890 41702 463932 41938
rect 461404 41660 463932 41702
rect 461404 41300 461724 41660
rect 460760 40980 461724 41300
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravan_logo  caravan_logo
timestamp 1636751500
transform 1 0 255300 0 1 6032
box 2240 2560 37000 11520
use caravan_motto  caravan_motto
timestamp 1637698689
transform 1 0 -54560 0 1 -52
box 367960 10204 399802 14768
use caravan_power_routing  caravan_power_routing
timestamp 1666269678
transform 1 0 0 0 1 0
box 6022 30806 711814 997678
use caravan_signal_routing  caravan_signal_routing
timestamp 1666277172
transform 1 0 0 0 1 0
box 39764 415548 677806 997846
use caravel_clocking  clock_ctrl
timestamp 1666097791
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use copyright_block_a  copyright_block_a
timestamp 1665519472
transform 1 0 149582 0 1 16298
box -262 -10162 35048 2764
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1665682149
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666126335
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666126335
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666126335
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666126335
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666126335
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666126335
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666126335
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666126335
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666126335
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666126335
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666126335
transform -1 0 710203 0 1 884800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666126335
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666126335
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666126335
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666126335
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666126335
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666126335
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666126335
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666126335
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666126335
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666126335
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666126335
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666126335
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666126335
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666126335
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666126335
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666126335
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1638587925
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1638587925
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1638587925
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1638587925
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1638587925
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1638587925
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1638587925
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1638587925
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1638587925
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1638587925
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1638587925
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1638587925
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1638587925
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1638587925
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1638587925
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1638587925
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1638587925
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1638587925
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1638587925
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1638587925
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1638587925
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1638587925
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1638587925
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1638587925
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1638587925
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1638587925
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1638587925
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666084955
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use mgmt_protect  mgmt_buffers
timestamp 1666114774
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use user_analog_project_wrapper  mprj
timestamp 1632839657
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use open_source  open_source
timestamp 1666123577
transform 1 0 206074 0 1 2336
box 752 5164 29030 16242
use chip_io_alt  padframe
timestamp 1666377896
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use digital_pll  pll
timestamp 1666101174
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1650914729
transform 1 0 650146 0 -1 55282
box -52 -62 11344 8684
use xres_buf  rstb_level
timestamp 1649268499
transform -1 0 145710 0 -1 50488
box 374 -400 3540 3800
use gpio_signal_buffering_alt  sigbuf
timestamp 1666028682
transform 1 0 0 0 1 0
box 40023 41960 677583 728321
use mgmt_core_wrapper  soc
timestamp 1665963385
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use spare_logic_block  spare_logic\[0\]
timestamp 1638030917
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1638030917
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1638030917
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1638030917
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use user_id_textblock  user_id_textblock
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use user_id_programming  user_id_value
timestamp 1650371074
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698624 953022 710789 965190 0 FreeSans 16000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628410 1018624 640578 1030789 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526610 1018624 538778 1030789 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475210 1018624 487378 1030789 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386210 1018624 398378 1030789 0 FreeSans 16000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284410 1018624 296578 1030789 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 231810 1018624 243978 1030789 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181410 1018624 193578 1030789 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 130010 1018624 142178 1030789 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78610 1018624 90778 1030789 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6811 956610 18976 968778 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144150 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19620 80934 0 FreeSans 16000 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 697980 909666 711433 920546 0 FreeSans 16000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19620 924934 0 FreeSans 16000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18976 0 FreeSans 16000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710789 831990 0 FreeSans 16000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710789 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18976 496578 0 FreeSans 16000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18976 123778 0 FreeSans 16000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18976 883378 0 FreeSans 16000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18976 0 FreeSans 16000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030789 0 FreeSans 16000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710789 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18976 841178 0 FreeSans 16000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19620 0 FreeSans 16000 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 697980 461866 711433 472746 0 FreeSans 16000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19620 453734 0 FreeSans 16000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18976 0 FreeSans 16000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030789 0 FreeSans 16000 0 0 0 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
