magic
tech sky130A
magscale 1 2
timestamp 1677077417
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< metal1 >>
rect 41866 995682 675734 995734
rect 41866 42225 41918 995682
rect 411070 42466 411076 42518
rect 411128 42506 411134 42518
rect 419718 42506 419724 42518
rect 411128 42478 419724 42506
rect 411128 42466 411134 42478
rect 419718 42466 419724 42478
rect 419776 42466 419782 42518
rect 465810 42476 465816 42528
rect 465868 42516 465874 42528
rect 474458 42516 474464 42528
rect 465868 42488 474464 42516
rect 465868 42476 465874 42488
rect 474458 42476 474464 42488
rect 474516 42476 474522 42528
rect 409230 42340 409236 42392
rect 409288 42380 409294 42392
rect 412266 42380 412272 42392
rect 409288 42352 412272 42380
rect 409288 42340 409294 42352
rect 412266 42340 412272 42352
rect 412324 42380 412330 42392
rect 415394 42380 415400 42392
rect 412324 42352 415400 42380
rect 412324 42340 412330 42352
rect 415394 42340 415400 42352
rect 415452 42340 415458 42392
rect 464004 42328 464010 42380
rect 464062 42368 464068 42380
rect 467040 42368 467046 42380
rect 464062 42340 467046 42368
rect 464062 42328 464068 42340
rect 467040 42328 467046 42340
rect 467098 42368 467104 42380
rect 470167 42368 470173 42380
rect 467098 42340 470173 42368
rect 467098 42328 467104 42340
rect 470167 42328 470173 42340
rect 470225 42328 470231 42380
rect 518802 42340 518808 42392
rect 518860 42380 518866 42392
rect 524966 42380 524972 42392
rect 518860 42352 524972 42380
rect 518860 42340 518866 42352
rect 524966 42340 524972 42352
rect 525024 42340 525030 42392
rect 675682 42225 675734 995682
rect 41866 42173 145063 42225
rect 145115 42173 145127 42225
rect 145179 42173 195328 42225
rect 195380 42173 199653 42225
rect 199705 42173 303929 42225
rect 303981 42173 308066 42225
rect 308118 42173 358732 42225
rect 358784 42173 363053 42225
rect 363105 42173 413524 42225
rect 413576 42173 417858 42225
rect 417910 42173 468330 42225
rect 468382 42173 472656 42225
rect 472708 42173 523126 42225
rect 523178 42173 527457 42225
rect 527509 42173 675734 42225
rect 186548 42089 188522 42141
rect 188574 42089 192845 42141
rect 192897 42089 201494 42141
rect 201546 42089 202717 42141
rect 202769 42089 202775 42141
rect 295162 42089 297125 42141
rect 297177 42089 299607 42141
rect 299659 42089 305774 42141
rect 305826 42089 311317 42141
rect 311369 42089 311375 42141
rect 349962 42089 351925 42141
rect 351977 42089 354406 42141
rect 354458 42089 360570 42141
rect 360622 42089 366117 42141
rect 366169 42089 366175 42141
rect 404762 42089 406719 42141
rect 406771 42089 420917 42141
rect 420969 42089 420975 42141
rect 459562 42089 461524 42141
rect 461576 42089 475717 42141
rect 475769 42089 475775 42141
rect 514362 42089 516320 42141
rect 516372 42089 530517 42141
rect 530569 42089 530575 42141
rect 186548 42005 189163 42057
rect 189215 42005 191003 42057
rect 191055 42005 192202 42057
rect 192254 42005 193489 42057
rect 193541 42005 196528 42057
rect 196580 42005 197170 42057
rect 197222 42005 197813 42057
rect 197865 42005 198368 42057
rect 198420 42005 200206 42057
rect 200258 42005 200857 42057
rect 200909 42005 205928 42057
rect 205980 42005 205986 42057
rect 295162 42005 297768 42057
rect 297820 42005 300804 42057
rect 300856 42005 301451 42057
rect 301503 42005 302094 42057
rect 302146 42005 302643 42057
rect 302695 42005 305133 42057
rect 305185 42005 306418 42057
rect 306470 42005 308809 42057
rect 308861 42005 309452 42057
rect 309504 42005 315497 42057
rect 315549 42005 315555 42057
rect 349962 42005 352568 42057
rect 352620 42005 355600 42057
rect 355652 42005 356246 42057
rect 356298 42005 356889 42057
rect 356941 42005 357444 42057
rect 357496 42005 359928 42057
rect 359980 42005 361217 42057
rect 361269 42005 363607 42057
rect 363659 42005 364252 42057
rect 364304 42005 370302 42057
rect 370354 42005 370360 42057
rect 404762 42005 407367 42057
rect 407419 42005 410398 42057
rect 410450 42005 411691 42057
rect 411743 42005 414725 42057
rect 414777 42005 416013 42057
rect 416065 42005 418404 42057
rect 418456 42005 419045 42057
rect 419097 42005 425115 42057
rect 425167 42005 425173 42057
rect 459562 42005 462162 42057
rect 462214 42005 465201 42057
rect 465253 42005 466488 42057
rect 466540 42005 469522 42057
rect 469574 42005 470810 42057
rect 470862 42005 473201 42057
rect 473253 42005 473849 42057
rect 473901 42005 479915 42057
rect 479967 42005 479973 42057
rect 514362 42005 516969 42057
rect 517021 42005 520004 42057
rect 520056 42005 521293 42057
rect 521345 42005 524328 42057
rect 524380 42005 525615 42057
rect 525667 42005 528009 42057
rect 528061 42005 528652 42057
rect 528704 42005 534772 42057
rect 534824 42005 534830 42057
rect 186548 41921 187968 41973
rect 188020 41921 195973 41973
rect 196025 41921 202162 41973
rect 295162 41921 296576 41973
rect 296628 41921 304577 41973
rect 304629 41921 310827 41973
rect 349962 41921 351375 41973
rect 351427 41921 359374 41973
rect 359426 41921 365627 41973
rect 404762 41921 406170 41973
rect 406222 41921 414174 41973
rect 414226 41921 420427 41973
rect 459562 41921 460971 41973
rect 461023 41921 468967 41973
rect 469019 41921 475227 41973
rect 514362 41921 515772 41973
rect 515824 41921 523773 41973
rect 523825 41921 530027 41973
rect 186548 41837 186683 41889
rect 186735 41837 194688 41889
rect 194740 41837 199012 41889
rect 199064 41837 202162 41889
rect 295162 41837 295283 41889
rect 295335 41837 303290 41889
rect 303342 41837 307616 41889
rect 307668 41837 310827 41889
rect 349962 41837 350086 41889
rect 350138 41837 358090 41889
rect 358142 41837 362412 41889
rect 362464 41837 365627 41889
rect 404762 41837 404877 41889
rect 404929 41837 412888 41889
rect 412940 41837 417210 41889
rect 417262 41837 420427 41889
rect 459562 41837 459678 41889
rect 459730 41837 467684 41889
rect 467736 41837 472010 41889
rect 472062 41837 475227 41889
rect 514362 41837 514487 41889
rect 514539 41837 522486 41889
rect 522538 41837 526810 41889
rect 526862 41837 530027 41889
rect 140990 40073 140996 40125
rect 141048 40118 141054 40125
rect 141986 40118 141992 40125
rect 141048 40080 141992 40118
rect 141048 40073 141054 40080
rect 141986 40073 141992 40080
rect 142044 40118 142050 40125
rect 143062 40118 143068 40125
rect 142044 40080 143068 40118
rect 142044 40073 142050 40080
rect 142573 40000 142619 40080
rect 143062 40073 143068 40080
rect 143120 40118 143126 40125
rect 143401 40118 143437 40125
rect 143120 40080 143437 40118
rect 143120 40073 143126 40080
rect 143401 40073 143437 40080
rect 143489 40118 143525 40125
rect 144597 40118 144603 40125
rect 143489 40080 144603 40118
rect 143489 40073 143525 40080
rect 144597 40073 144603 40080
rect 144655 40073 144661 40125
<< via1 >>
rect 411076 42466 411128 42518
rect 419724 42466 419776 42518
rect 465816 42476 465868 42528
rect 474464 42476 474516 42528
rect 409236 42340 409288 42392
rect 412272 42340 412324 42392
rect 415400 42340 415452 42392
rect 464010 42328 464062 42380
rect 467046 42328 467098 42380
rect 470173 42328 470225 42380
rect 518808 42340 518860 42392
rect 524972 42340 525024 42392
rect 145063 42173 145115 42225
rect 145127 42173 145179 42225
rect 195328 42173 195380 42225
rect 199653 42173 199705 42225
rect 303929 42173 303981 42225
rect 308066 42173 308118 42225
rect 358732 42173 358784 42225
rect 363053 42173 363105 42225
rect 413524 42173 413576 42225
rect 417858 42173 417910 42225
rect 468330 42173 468382 42225
rect 472656 42173 472708 42225
rect 523126 42173 523178 42225
rect 527457 42173 527509 42225
rect 188522 42089 188574 42141
rect 192845 42089 192897 42141
rect 201494 42089 201546 42141
rect 202717 42089 202769 42141
rect 297125 42089 297177 42141
rect 299607 42089 299659 42141
rect 305774 42089 305826 42141
rect 311317 42089 311369 42141
rect 351925 42089 351977 42141
rect 354406 42089 354458 42141
rect 360570 42089 360622 42141
rect 366117 42089 366169 42141
rect 406719 42089 406771 42141
rect 420917 42089 420969 42141
rect 461524 42089 461576 42141
rect 475717 42089 475769 42141
rect 516320 42089 516372 42141
rect 530517 42089 530569 42141
rect 189163 42005 189215 42057
rect 191003 42005 191055 42057
rect 192202 42005 192254 42057
rect 193489 42005 193541 42057
rect 196528 42005 196580 42057
rect 197170 42005 197222 42057
rect 197813 42005 197865 42057
rect 198368 42005 198420 42057
rect 200206 42005 200258 42057
rect 200857 42005 200909 42057
rect 205928 42005 205980 42057
rect 297768 42005 297820 42057
rect 300804 42005 300856 42057
rect 301451 42005 301503 42057
rect 302094 42005 302146 42057
rect 302643 42005 302695 42057
rect 305133 42005 305185 42057
rect 306418 42005 306470 42057
rect 308809 42005 308861 42057
rect 309452 42005 309504 42057
rect 315497 42005 315549 42057
rect 352568 42005 352620 42057
rect 355600 42005 355652 42057
rect 356246 42005 356298 42057
rect 356889 42005 356941 42057
rect 357444 42005 357496 42057
rect 359928 42005 359980 42057
rect 361217 42005 361269 42057
rect 363607 42005 363659 42057
rect 364252 42005 364304 42057
rect 370302 42005 370354 42057
rect 407367 42005 407419 42057
rect 410398 42005 410450 42057
rect 411691 42005 411743 42057
rect 414725 42005 414777 42057
rect 416013 42005 416065 42057
rect 418404 42005 418456 42057
rect 419045 42005 419097 42057
rect 425115 42005 425167 42057
rect 462162 42005 462214 42057
rect 465201 42005 465253 42057
rect 466488 42005 466540 42057
rect 469522 42005 469574 42057
rect 470810 42005 470862 42057
rect 473201 42005 473253 42057
rect 473849 42005 473901 42057
rect 479915 42005 479967 42057
rect 516969 42005 517021 42057
rect 520004 42005 520056 42057
rect 521293 42005 521345 42057
rect 524328 42005 524380 42057
rect 525615 42005 525667 42057
rect 528009 42005 528061 42057
rect 528652 42005 528704 42057
rect 534772 42005 534824 42057
rect 187968 41921 188020 41973
rect 195973 41921 196025 41973
rect 296576 41921 296628 41973
rect 304577 41921 304629 41973
rect 351375 41921 351427 41973
rect 359374 41921 359426 41973
rect 406170 41921 406222 41973
rect 414174 41921 414226 41973
rect 460971 41921 461023 41973
rect 468967 41921 469019 41973
rect 515772 41921 515824 41973
rect 523773 41921 523825 41973
rect 186683 41837 186735 41889
rect 194688 41837 194740 41889
rect 199012 41837 199064 41889
rect 295283 41837 295335 41889
rect 303290 41837 303342 41889
rect 307616 41837 307668 41889
rect 350086 41837 350138 41889
rect 358090 41837 358142 41889
rect 362412 41837 362464 41889
rect 404877 41837 404929 41889
rect 412888 41837 412940 41889
rect 417210 41837 417262 41889
rect 459678 41837 459730 41889
rect 467684 41837 467736 41889
rect 472010 41837 472062 41889
rect 514487 41837 514539 41889
rect 522486 41837 522538 41889
rect 526810 41837 526862 41889
rect 140996 40073 141048 40125
rect 141992 40073 142044 40125
rect 143068 40073 143120 40125
rect 143437 40073 143489 40125
rect 144603 40073 144655 40125
<< metal2 >>
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 90021 995407 90077 995887
rect 91217 995407 91273 995887
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 141421 995407 141477 995887
rect 142617 995407 142673 995887
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 192821 995407 192877 995887
rect 194017 995407 194073 995887
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 244221 995407 244277 995887
rect 245417 995407 245473 995887
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 295821 995407 295877 995887
rect 297017 995407 297073 995887
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 397621 995407 397677 995887
rect 398817 995407 398873 995887
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 486621 995407 486677 995887
rect 487817 995407 487873 995887
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 538021 995407 538077 995887
rect 539217 995407 539273 995887
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 639821 995407 639877 995887
rect 641017 995407 641073 995887
rect 41863 969273 42193 969280
rect 41713 969217 41883 969273
rect 41939 969217 41963 969273
rect 42019 969217 42043 969273
rect 42099 969217 42123 969273
rect 42179 969217 42193 969273
rect 41863 969210 42193 969217
rect 41863 968077 42193 968084
rect 41713 968021 41883 968077
rect 41939 968021 41963 968077
rect 42019 968021 42043 968077
rect 42099 968021 42123 968077
rect 42179 968021 42193 968077
rect 41863 968014 42193 968021
rect 41863 967433 42193 967440
rect 41713 967377 41883 967433
rect 41939 967377 41963 967433
rect 42019 967377 42043 967433
rect 42099 967377 42123 967433
rect 42179 967377 42193 967433
rect 41863 967370 42193 967377
rect 41863 966789 42193 966796
rect 41713 966733 41883 966789
rect 41939 966733 41963 966789
rect 42019 966733 42043 966789
rect 42099 966733 42123 966789
rect 42179 966733 42193 966789
rect 41863 966726 42193 966733
rect 675407 966751 675737 966758
rect 675407 966695 675427 966751
rect 675483 966695 675507 966751
rect 675563 966695 675587 966751
rect 675643 966695 675667 966751
rect 675723 966695 675887 966751
rect 675407 966688 675737 966695
rect 675407 966107 675737 966114
rect 675407 966051 675427 966107
rect 675483 966051 675507 966107
rect 675563 966051 675587 966107
rect 675643 966051 675667 966107
rect 675723 966051 675887 966107
rect 675407 966044 675737 966051
rect 41863 965593 42193 965600
rect 41713 965537 41883 965593
rect 41939 965537 41963 965593
rect 42019 965537 42043 965593
rect 42099 965537 42123 965593
rect 42179 965537 42193 965593
rect 41863 965530 42193 965537
rect 675407 965463 675737 965470
rect 675407 965407 675427 965463
rect 675483 965407 675507 965463
rect 675563 965407 675587 965463
rect 675643 965407 675667 965463
rect 675723 965407 675887 965463
rect 675407 965400 675737 965407
rect 41863 964397 42193 964404
rect 41713 964341 41883 964397
rect 41939 964341 41963 964397
rect 42019 964341 42043 964397
rect 42099 964341 42123 964397
rect 42179 964341 42193 964397
rect 41863 964334 42193 964341
rect 41863 963753 42193 963760
rect 41713 963697 41883 963753
rect 41939 963697 41963 963753
rect 42019 963697 42043 963753
rect 42099 963697 42123 963753
rect 42179 963697 42193 963753
rect 41863 963690 42193 963697
rect 675407 963623 675737 963630
rect 675407 963567 675427 963623
rect 675483 963567 675507 963623
rect 675563 963567 675587 963623
rect 675643 963567 675667 963623
rect 675723 963567 675887 963623
rect 675407 963560 675737 963567
rect 41863 963109 42193 963116
rect 41713 963053 41883 963109
rect 41939 963053 41963 963109
rect 42019 963053 42043 963109
rect 42099 963053 42123 963109
rect 42179 963053 42193 963109
rect 41863 963046 42193 963053
rect 675407 963071 675737 963078
rect 675407 963015 675427 963071
rect 675483 963015 675507 963071
rect 675563 963015 675587 963071
rect 675643 963015 675667 963071
rect 675723 963015 675887 963071
rect 675407 963008 675737 963015
rect 41863 962557 42193 962564
rect 41713 962501 41883 962557
rect 41939 962501 41963 962557
rect 42019 962501 42043 962557
rect 42099 962501 42123 962557
rect 42179 962501 42193 962557
rect 41863 962494 42193 962501
rect 675407 962427 675737 962434
rect 675407 962371 675427 962427
rect 675483 962371 675507 962427
rect 675563 962371 675587 962427
rect 675643 962371 675667 962427
rect 675723 962371 675887 962427
rect 675407 962364 675737 962371
rect 675407 961783 675737 961790
rect 675407 961727 675427 961783
rect 675483 961727 675507 961783
rect 675563 961727 675587 961783
rect 675643 961727 675667 961783
rect 675723 961727 675887 961783
rect 675407 961720 675737 961727
rect 41863 960073 42193 960080
rect 41713 960017 41883 960073
rect 41939 960017 41963 960073
rect 42019 960017 42043 960073
rect 42099 960017 42123 960073
rect 42179 960017 42193 960073
rect 41863 960010 42193 960017
rect 41863 959429 42193 959436
rect 41713 959373 41883 959429
rect 41939 959373 41963 959429
rect 42019 959373 42043 959429
rect 42099 959373 42123 959429
rect 42179 959373 42193 959429
rect 41863 959366 42193 959373
rect 675407 959299 675737 959306
rect 675407 959243 675427 959299
rect 675483 959243 675507 959299
rect 675563 959243 675587 959299
rect 675643 959243 675667 959299
rect 675723 959243 675887 959299
rect 675407 959236 675737 959243
rect 41863 958785 42193 958792
rect 41713 958729 41883 958785
rect 41939 958729 41963 958785
rect 42019 958729 42043 958785
rect 42099 958729 42123 958785
rect 42179 958729 42193 958785
rect 41863 958722 42193 958729
rect 675407 958747 675737 958754
rect 675407 958691 675427 958747
rect 675483 958691 675507 958747
rect 675563 958691 675587 958747
rect 675643 958691 675667 958747
rect 675723 958691 675887 958747
rect 675407 958684 675737 958691
rect 41863 958233 42193 958240
rect 41713 958177 41883 958233
rect 41939 958177 41963 958233
rect 42019 958177 42043 958233
rect 42099 958177 42123 958233
rect 42179 958177 42193 958233
rect 41863 958170 42193 958177
rect 675407 958103 675737 958110
rect 675407 958047 675427 958103
rect 675483 958047 675507 958103
rect 675563 958047 675587 958103
rect 675643 958047 675667 958103
rect 675723 958047 675887 958103
rect 675407 958040 675737 958047
rect 675407 957459 675737 957466
rect 675407 957403 675427 957459
rect 675483 957403 675507 957459
rect 675563 957403 675587 957459
rect 675643 957403 675667 957459
rect 675723 957403 675887 957459
rect 675407 957396 675737 957403
rect 41863 956393 42193 956400
rect 41713 956337 41883 956393
rect 41939 956337 41963 956393
rect 42019 956337 42043 956393
rect 42099 956337 42123 956393
rect 42179 956337 42193 956393
rect 41863 956330 42193 956337
rect 675407 956263 675737 956270
rect 675407 956207 675427 956263
rect 675483 956207 675507 956263
rect 675563 956207 675587 956263
rect 675643 956207 675667 956263
rect 675723 956207 675887 956263
rect 675407 956200 675737 956207
rect 41863 955749 42193 955756
rect 41713 955693 41883 955749
rect 41939 955693 41963 955749
rect 42019 955693 42043 955749
rect 42099 955693 42123 955749
rect 42179 955693 42193 955749
rect 41863 955686 42193 955693
rect 41863 955105 42193 955112
rect 41713 955049 41883 955105
rect 41939 955049 41963 955105
rect 42019 955049 42043 955105
rect 42099 955049 42123 955105
rect 42179 955049 42193 955105
rect 41863 955042 42193 955049
rect 675407 955067 675737 955074
rect 675407 955011 675427 955067
rect 675483 955011 675507 955067
rect 675563 955011 675587 955067
rect 675643 955011 675667 955067
rect 675723 955011 675887 955067
rect 675407 955004 675737 955011
rect 675407 954423 675737 954430
rect 675407 954367 675427 954423
rect 675483 954367 675507 954423
rect 675563 954367 675587 954423
rect 675643 954367 675667 954423
rect 675723 954367 675887 954423
rect 675407 954360 675737 954367
rect 675407 953779 675737 953786
rect 675407 953723 675427 953779
rect 675483 953723 675507 953779
rect 675563 953723 675587 953779
rect 675643 953723 675667 953779
rect 675723 953723 675887 953779
rect 675407 953716 675737 953723
rect 675407 952583 675737 952590
rect 675407 952527 675427 952583
rect 675483 952527 675507 952583
rect 675563 952527 675587 952583
rect 675643 952527 675667 952583
rect 675723 952527 675887 952583
rect 675407 952520 675737 952527
rect 675407 877551 675737 877558
rect 675407 877495 675427 877551
rect 675483 877495 675507 877551
rect 675563 877495 675587 877551
rect 675643 877495 675667 877551
rect 675723 877495 675887 877551
rect 675407 877488 675737 877495
rect 675407 876907 675737 876914
rect 675407 876851 675427 876907
rect 675483 876851 675507 876907
rect 675563 876851 675587 876907
rect 675643 876851 675667 876907
rect 675723 876851 675887 876907
rect 675407 876844 675737 876851
rect 675407 876263 675737 876270
rect 675407 876207 675427 876263
rect 675483 876207 675507 876263
rect 675563 876207 675587 876263
rect 675643 876207 675667 876263
rect 675723 876207 675887 876263
rect 675407 876200 675737 876207
rect 675407 874423 675737 874430
rect 675407 874367 675427 874423
rect 675483 874367 675507 874423
rect 675563 874367 675587 874423
rect 675643 874367 675667 874423
rect 675723 874367 675887 874423
rect 675407 874360 675737 874367
rect 675407 873871 675737 873878
rect 675407 873815 675427 873871
rect 675483 873815 675507 873871
rect 675563 873815 675587 873871
rect 675643 873815 675667 873871
rect 675723 873815 675887 873871
rect 675407 873808 675737 873815
rect 675407 873227 675737 873234
rect 675407 873171 675427 873227
rect 675483 873171 675507 873227
rect 675563 873171 675587 873227
rect 675643 873171 675667 873227
rect 675723 873171 675887 873227
rect 675407 873164 675737 873171
rect 675407 872583 675737 872590
rect 675407 872527 675427 872583
rect 675483 872527 675507 872583
rect 675563 872527 675587 872583
rect 675643 872527 675667 872583
rect 675723 872527 675887 872583
rect 675407 872520 675737 872527
rect 675407 870099 675737 870106
rect 675407 870043 675427 870099
rect 675483 870043 675507 870099
rect 675563 870043 675587 870099
rect 675643 870043 675667 870099
rect 675723 870043 675887 870099
rect 675407 870036 675737 870043
rect 675407 869547 675737 869554
rect 675407 869491 675427 869547
rect 675483 869491 675507 869547
rect 675563 869491 675587 869547
rect 675643 869491 675667 869547
rect 675723 869491 675887 869547
rect 675407 869484 675737 869491
rect 675407 868903 675737 868910
rect 675407 868847 675427 868903
rect 675483 868847 675507 868903
rect 675563 868847 675587 868903
rect 675643 868847 675667 868903
rect 675723 868847 675887 868903
rect 675407 868840 675737 868847
rect 675407 868259 675737 868266
rect 675407 868203 675427 868259
rect 675483 868203 675507 868259
rect 675563 868203 675587 868259
rect 675643 868203 675667 868259
rect 675723 868203 675887 868259
rect 675407 868196 675737 868203
rect 675407 867063 675737 867070
rect 675407 867007 675427 867063
rect 675483 867007 675507 867063
rect 675563 867007 675587 867063
rect 675643 867007 675667 867063
rect 675723 867007 675887 867063
rect 675407 867000 675737 867007
rect 675407 865867 675737 865874
rect 675407 865811 675427 865867
rect 675483 865811 675507 865867
rect 675563 865811 675587 865867
rect 675643 865811 675667 865867
rect 675723 865811 675887 865867
rect 675407 865804 675737 865811
rect 675407 865223 675737 865230
rect 675407 865167 675427 865223
rect 675483 865167 675507 865223
rect 675563 865167 675587 865223
rect 675643 865167 675667 865223
rect 675723 865167 675887 865223
rect 675407 865160 675737 865167
rect 675407 864579 675737 864586
rect 675407 864523 675427 864579
rect 675483 864523 675507 864579
rect 675563 864523 675587 864579
rect 675643 864523 675667 864579
rect 675723 864523 675887 864579
rect 675407 864516 675737 864523
rect 675407 863383 675737 863390
rect 675407 863327 675427 863383
rect 675483 863327 675507 863383
rect 675563 863327 675587 863383
rect 675643 863327 675667 863383
rect 675723 863327 675887 863383
rect 675407 863320 675737 863327
rect 41863 799473 42193 799480
rect 41713 799417 41883 799473
rect 41939 799417 41963 799473
rect 42019 799417 42043 799473
rect 42099 799417 42123 799473
rect 42179 799417 42193 799473
rect 41863 799410 42193 799417
rect 41863 798277 42193 798284
rect 41713 798221 41883 798277
rect 41939 798221 41963 798277
rect 42019 798221 42043 798277
rect 42099 798221 42123 798277
rect 42179 798221 42193 798277
rect 41863 798214 42193 798221
rect 41863 797633 42193 797640
rect 41713 797577 41883 797633
rect 41939 797577 41963 797633
rect 42019 797577 42043 797633
rect 42099 797577 42123 797633
rect 42179 797577 42193 797633
rect 41863 797570 42193 797577
rect 41863 796989 42193 796996
rect 41713 796933 41883 796989
rect 41939 796933 41963 796989
rect 42019 796933 42043 796989
rect 42099 796933 42123 796989
rect 42179 796933 42193 796989
rect 41863 796926 42193 796933
rect 41863 795793 42193 795800
rect 41713 795737 41883 795793
rect 41939 795737 41963 795793
rect 42019 795737 42043 795793
rect 42099 795737 42123 795793
rect 42179 795737 42193 795793
rect 41863 795730 42193 795737
rect 41863 794597 42193 794604
rect 41713 794541 41883 794597
rect 41939 794541 41963 794597
rect 42019 794541 42043 794597
rect 42099 794541 42123 794597
rect 42179 794541 42193 794597
rect 41863 794534 42193 794541
rect 41863 793953 42193 793960
rect 41713 793897 41883 793953
rect 41939 793897 41963 793953
rect 42019 793897 42043 793953
rect 42099 793897 42123 793953
rect 42179 793897 42193 793953
rect 41863 793890 42193 793897
rect 41863 793309 42193 793316
rect 41713 793253 41883 793309
rect 41939 793253 41963 793309
rect 42019 793253 42043 793309
rect 42099 793253 42123 793309
rect 42179 793253 42193 793309
rect 41863 793246 42193 793253
rect 41863 792757 42193 792764
rect 41713 792701 41883 792757
rect 41939 792701 41963 792757
rect 42019 792701 42043 792757
rect 42099 792701 42123 792757
rect 42179 792701 42193 792757
rect 41863 792694 42193 792701
rect 41863 790273 42193 790280
rect 41713 790217 41883 790273
rect 41939 790217 41963 790273
rect 42019 790217 42043 790273
rect 42099 790217 42123 790273
rect 42179 790217 42193 790273
rect 41863 790210 42193 790217
rect 41863 789629 42193 789636
rect 41713 789573 41883 789629
rect 41939 789573 41963 789629
rect 42019 789573 42043 789629
rect 42099 789573 42123 789629
rect 42179 789573 42193 789629
rect 41863 789566 42193 789573
rect 41863 788985 42193 788992
rect 41713 788929 41883 788985
rect 41939 788929 41963 788985
rect 42019 788929 42043 788985
rect 42099 788929 42123 788985
rect 42179 788929 42193 788985
rect 41863 788922 42193 788929
rect 41863 788433 42193 788440
rect 41713 788377 41883 788433
rect 41939 788377 41963 788433
rect 42019 788377 42043 788433
rect 42099 788377 42123 788433
rect 42179 788377 42193 788433
rect 41863 788370 42193 788377
rect 675407 788351 675737 788358
rect 675407 788295 675427 788351
rect 675483 788295 675507 788351
rect 675563 788295 675587 788351
rect 675643 788295 675667 788351
rect 675723 788295 675887 788351
rect 675407 788288 675737 788295
rect 675407 787707 675737 787714
rect 675407 787651 675427 787707
rect 675483 787651 675507 787707
rect 675563 787651 675587 787707
rect 675643 787651 675667 787707
rect 675723 787651 675887 787707
rect 675407 787644 675737 787651
rect 675407 787063 675737 787070
rect 675407 787007 675427 787063
rect 675483 787007 675507 787063
rect 675563 787007 675587 787063
rect 675643 787007 675667 787063
rect 675723 787007 675887 787063
rect 675407 787000 675737 787007
rect 41863 786593 42193 786600
rect 41713 786537 41883 786593
rect 41939 786537 41963 786593
rect 42019 786537 42043 786593
rect 42099 786537 42123 786593
rect 42179 786537 42193 786593
rect 41863 786530 42193 786537
rect 41863 785949 42193 785956
rect 41713 785893 41883 785949
rect 41939 785893 41963 785949
rect 42019 785893 42043 785949
rect 42099 785893 42123 785949
rect 42179 785893 42193 785949
rect 41863 785886 42193 785893
rect 41863 785305 42193 785312
rect 41713 785249 41883 785305
rect 41939 785249 41963 785305
rect 42019 785249 42043 785305
rect 42099 785249 42123 785305
rect 42179 785249 42193 785305
rect 41863 785242 42193 785249
rect 675407 785223 675737 785230
rect 675407 785167 675427 785223
rect 675483 785167 675507 785223
rect 675563 785167 675587 785223
rect 675643 785167 675667 785223
rect 675723 785167 675887 785223
rect 675407 785160 675737 785167
rect 675407 784671 675737 784678
rect 675407 784615 675427 784671
rect 675483 784615 675507 784671
rect 675563 784615 675587 784671
rect 675643 784615 675667 784671
rect 675723 784615 675887 784671
rect 675407 784608 675737 784615
rect 675407 784027 675737 784034
rect 675407 783971 675427 784027
rect 675483 783971 675507 784027
rect 675563 783971 675587 784027
rect 675643 783971 675667 784027
rect 675723 783971 675887 784027
rect 675407 783964 675737 783971
rect 675407 783383 675737 783390
rect 675407 783327 675427 783383
rect 675483 783327 675507 783383
rect 675563 783327 675587 783383
rect 675643 783327 675667 783383
rect 675723 783327 675887 783383
rect 675407 783320 675737 783327
rect 675407 780899 675737 780906
rect 675407 780843 675427 780899
rect 675483 780843 675507 780899
rect 675563 780843 675587 780899
rect 675643 780843 675667 780899
rect 675723 780843 675887 780899
rect 675407 780836 675737 780843
rect 675407 780347 675737 780354
rect 675407 780291 675427 780347
rect 675483 780291 675507 780347
rect 675563 780291 675587 780347
rect 675643 780291 675667 780347
rect 675723 780291 675887 780347
rect 675407 780284 675737 780291
rect 675407 779703 675737 779710
rect 675407 779647 675427 779703
rect 675483 779647 675507 779703
rect 675563 779647 675587 779703
rect 675643 779647 675667 779703
rect 675723 779647 675887 779703
rect 675407 779640 675737 779647
rect 675407 779059 675737 779066
rect 675407 779003 675427 779059
rect 675483 779003 675507 779059
rect 675563 779003 675587 779059
rect 675643 779003 675667 779059
rect 675723 779003 675887 779059
rect 675407 778996 675737 779003
rect 675407 777863 675737 777870
rect 675407 777807 675427 777863
rect 675483 777807 675507 777863
rect 675563 777807 675587 777863
rect 675643 777807 675667 777863
rect 675723 777807 675887 777863
rect 675407 777800 675737 777807
rect 675407 776667 675737 776674
rect 675407 776611 675427 776667
rect 675483 776611 675507 776667
rect 675563 776611 675587 776667
rect 675643 776611 675667 776667
rect 675723 776611 675887 776667
rect 675407 776604 675737 776611
rect 675407 776023 675737 776030
rect 675407 775967 675427 776023
rect 675483 775967 675507 776023
rect 675563 775967 675587 776023
rect 675643 775967 675667 776023
rect 675723 775967 675887 776023
rect 675407 775960 675737 775967
rect 675407 775379 675737 775386
rect 675407 775323 675427 775379
rect 675483 775323 675507 775379
rect 675563 775323 675587 775379
rect 675643 775323 675667 775379
rect 675723 775323 675887 775379
rect 675407 775316 675737 775323
rect 675407 774183 675737 774190
rect 675407 774127 675427 774183
rect 675483 774127 675507 774183
rect 675563 774127 675587 774183
rect 675643 774127 675667 774183
rect 675723 774127 675887 774183
rect 675407 774120 675737 774127
rect 41863 756273 42193 756280
rect 41713 756217 41883 756273
rect 41939 756217 41963 756273
rect 42019 756217 42043 756273
rect 42099 756217 42123 756273
rect 42179 756217 42193 756273
rect 41863 756210 42193 756217
rect 41863 755077 42193 755084
rect 41713 755021 41883 755077
rect 41939 755021 41963 755077
rect 42019 755021 42043 755077
rect 42099 755021 42123 755077
rect 42179 755021 42193 755077
rect 41863 755014 42193 755021
rect 41863 754433 42193 754440
rect 41713 754377 41883 754433
rect 41939 754377 41963 754433
rect 42019 754377 42043 754433
rect 42099 754377 42123 754433
rect 42179 754377 42193 754433
rect 41863 754370 42193 754377
rect 41863 753789 42193 753796
rect 41713 753733 41883 753789
rect 41939 753733 41963 753789
rect 42019 753733 42043 753789
rect 42099 753733 42123 753789
rect 42179 753733 42193 753789
rect 41863 753726 42193 753733
rect 41863 752593 42193 752600
rect 41713 752537 41883 752593
rect 41939 752537 41963 752593
rect 42019 752537 42043 752593
rect 42099 752537 42123 752593
rect 42179 752537 42193 752593
rect 41863 752530 42193 752537
rect 41863 751397 42193 751404
rect 41713 751341 41883 751397
rect 41939 751341 41963 751397
rect 42019 751341 42043 751397
rect 42099 751341 42123 751397
rect 42179 751341 42193 751397
rect 41863 751334 42193 751341
rect 41863 750753 42193 750760
rect 41713 750697 41883 750753
rect 41939 750697 41963 750753
rect 42019 750697 42043 750753
rect 42099 750697 42123 750753
rect 42179 750697 42193 750753
rect 41863 750690 42193 750697
rect 41863 750109 42193 750116
rect 41713 750053 41883 750109
rect 41939 750053 41963 750109
rect 42019 750053 42043 750109
rect 42099 750053 42123 750109
rect 42179 750053 42193 750109
rect 41863 750046 42193 750053
rect 41863 749557 42193 749564
rect 41713 749501 41883 749557
rect 41939 749501 41963 749557
rect 42019 749501 42043 749557
rect 42099 749501 42123 749557
rect 42179 749501 42193 749557
rect 41863 749494 42193 749501
rect 41863 747073 42193 747080
rect 41713 747017 41883 747073
rect 41939 747017 41963 747073
rect 42019 747017 42043 747073
rect 42099 747017 42123 747073
rect 42179 747017 42193 747073
rect 41863 747010 42193 747017
rect 41863 746429 42193 746436
rect 41713 746373 41883 746429
rect 41939 746373 41963 746429
rect 42019 746373 42043 746429
rect 42099 746373 42123 746429
rect 42179 746373 42193 746429
rect 41863 746366 42193 746373
rect 41863 745785 42193 745792
rect 41713 745729 41883 745785
rect 41939 745729 41963 745785
rect 42019 745729 42043 745785
rect 42099 745729 42123 745785
rect 42179 745729 42193 745785
rect 41863 745722 42193 745729
rect 41863 745233 42193 745240
rect 41713 745177 41883 745233
rect 41939 745177 41963 745233
rect 42019 745177 42043 745233
rect 42099 745177 42123 745233
rect 42179 745177 42193 745233
rect 41863 745170 42193 745177
rect 41863 743393 42193 743400
rect 41713 743337 41883 743393
rect 41939 743337 41963 743393
rect 42019 743337 42043 743393
rect 42099 743337 42123 743393
rect 42179 743337 42193 743393
rect 41863 743330 42193 743337
rect 675407 743351 675737 743358
rect 675407 743295 675427 743351
rect 675483 743295 675507 743351
rect 675563 743295 675587 743351
rect 675643 743295 675667 743351
rect 675723 743295 675887 743351
rect 675407 743288 675737 743295
rect 41863 742749 42193 742756
rect 41713 742693 41883 742749
rect 41939 742693 41963 742749
rect 42019 742693 42043 742749
rect 42099 742693 42123 742749
rect 42179 742693 42193 742749
rect 41863 742686 42193 742693
rect 675407 742707 675737 742714
rect 675407 742651 675427 742707
rect 675483 742651 675507 742707
rect 675563 742651 675587 742707
rect 675643 742651 675667 742707
rect 675723 742651 675887 742707
rect 675407 742644 675737 742651
rect 41863 742105 42193 742112
rect 41713 742049 41883 742105
rect 41939 742049 41963 742105
rect 42019 742049 42043 742105
rect 42099 742049 42123 742105
rect 42179 742049 42193 742105
rect 41863 742042 42193 742049
rect 675407 742063 675737 742070
rect 675407 742007 675427 742063
rect 675483 742007 675507 742063
rect 675563 742007 675587 742063
rect 675643 742007 675667 742063
rect 675723 742007 675887 742063
rect 675407 742000 675737 742007
rect 675407 740223 675737 740230
rect 675407 740167 675427 740223
rect 675483 740167 675507 740223
rect 675563 740167 675587 740223
rect 675643 740167 675667 740223
rect 675723 740167 675887 740223
rect 675407 740160 675737 740167
rect 675407 739671 675737 739678
rect 675407 739615 675427 739671
rect 675483 739615 675507 739671
rect 675563 739615 675587 739671
rect 675643 739615 675667 739671
rect 675723 739615 675887 739671
rect 675407 739608 675737 739615
rect 675407 739027 675737 739034
rect 675407 738971 675427 739027
rect 675483 738971 675507 739027
rect 675563 738971 675587 739027
rect 675643 738971 675667 739027
rect 675723 738971 675887 739027
rect 675407 738964 675737 738971
rect 675407 738383 675737 738390
rect 675407 738327 675427 738383
rect 675483 738327 675507 738383
rect 675563 738327 675587 738383
rect 675643 738327 675667 738383
rect 675723 738327 675887 738383
rect 675407 738320 675737 738327
rect 675407 735899 675737 735906
rect 675407 735843 675427 735899
rect 675483 735843 675507 735899
rect 675563 735843 675587 735899
rect 675643 735843 675667 735899
rect 675723 735843 675887 735899
rect 675407 735836 675737 735843
rect 675407 735347 675737 735354
rect 675407 735291 675427 735347
rect 675483 735291 675507 735347
rect 675563 735291 675587 735347
rect 675643 735291 675667 735347
rect 675723 735291 675887 735347
rect 675407 735284 675737 735291
rect 675407 734703 675737 734710
rect 675407 734647 675427 734703
rect 675483 734647 675507 734703
rect 675563 734647 675587 734703
rect 675643 734647 675667 734703
rect 675723 734647 675887 734703
rect 675407 734640 675737 734647
rect 675407 734059 675737 734066
rect 675407 734003 675427 734059
rect 675483 734003 675507 734059
rect 675563 734003 675587 734059
rect 675643 734003 675667 734059
rect 675723 734003 675887 734059
rect 675407 733996 675737 734003
rect 675407 732863 675737 732870
rect 675407 732807 675427 732863
rect 675483 732807 675507 732863
rect 675563 732807 675587 732863
rect 675643 732807 675667 732863
rect 675723 732807 675887 732863
rect 675407 732800 675737 732807
rect 675407 731667 675737 731674
rect 675407 731611 675427 731667
rect 675483 731611 675507 731667
rect 675563 731611 675587 731667
rect 675643 731611 675667 731667
rect 675723 731611 675887 731667
rect 675407 731604 675737 731611
rect 675407 731023 675737 731030
rect 675407 730967 675427 731023
rect 675483 730967 675507 731023
rect 675563 730967 675587 731023
rect 675643 730967 675667 731023
rect 675723 730967 675887 731023
rect 675407 730960 675737 730967
rect 675407 730379 675737 730386
rect 675407 730323 675427 730379
rect 675483 730323 675507 730379
rect 675563 730323 675587 730379
rect 675643 730323 675667 730379
rect 675723 730323 675887 730379
rect 675407 730316 675737 730323
rect 675407 729183 675737 729190
rect 675407 729127 675427 729183
rect 675483 729127 675507 729183
rect 675563 729127 675587 729183
rect 675643 729127 675667 729183
rect 675723 729127 675887 729183
rect 675407 729120 675737 729127
rect 41863 713073 42193 713080
rect 41713 713017 41883 713073
rect 41939 713017 41963 713073
rect 42019 713017 42043 713073
rect 42099 713017 42123 713073
rect 42179 713017 42193 713073
rect 41863 713010 42193 713017
rect 41863 711877 42193 711884
rect 41713 711821 41883 711877
rect 41939 711821 41963 711877
rect 42019 711821 42043 711877
rect 42099 711821 42123 711877
rect 42179 711821 42193 711877
rect 41863 711814 42193 711821
rect 41863 711233 42193 711240
rect 41713 711177 41883 711233
rect 41939 711177 41963 711233
rect 42019 711177 42043 711233
rect 42099 711177 42123 711233
rect 42179 711177 42193 711233
rect 41863 711170 42193 711177
rect 41863 710589 42193 710596
rect 41713 710533 41883 710589
rect 41939 710533 41963 710589
rect 42019 710533 42043 710589
rect 42099 710533 42123 710589
rect 42179 710533 42193 710589
rect 41863 710526 42193 710533
rect 41863 709393 42193 709400
rect 41713 709337 41883 709393
rect 41939 709337 41963 709393
rect 42019 709337 42043 709393
rect 42099 709337 42123 709393
rect 42179 709337 42193 709393
rect 41863 709330 42193 709337
rect 41863 708197 42193 708204
rect 41713 708141 41883 708197
rect 41939 708141 41963 708197
rect 42019 708141 42043 708197
rect 42099 708141 42123 708197
rect 42179 708141 42193 708197
rect 41863 708134 42193 708141
rect 41863 707553 42193 707560
rect 41713 707497 41883 707553
rect 41939 707497 41963 707553
rect 42019 707497 42043 707553
rect 42099 707497 42123 707553
rect 42179 707497 42193 707553
rect 41863 707490 42193 707497
rect 41863 706909 42193 706916
rect 41713 706853 41883 706909
rect 41939 706853 41963 706909
rect 42019 706853 42043 706909
rect 42099 706853 42123 706909
rect 42179 706853 42193 706909
rect 41863 706846 42193 706853
rect 41863 706357 42193 706364
rect 41713 706301 41883 706357
rect 41939 706301 41963 706357
rect 42019 706301 42043 706357
rect 42099 706301 42123 706357
rect 42179 706301 42193 706357
rect 41863 706294 42193 706301
rect 41863 703873 42193 703880
rect 41713 703817 41883 703873
rect 41939 703817 41963 703873
rect 42019 703817 42043 703873
rect 42099 703817 42123 703873
rect 42179 703817 42193 703873
rect 41863 703810 42193 703817
rect 41863 703229 42193 703236
rect 41713 703173 41883 703229
rect 41939 703173 41963 703229
rect 42019 703173 42043 703229
rect 42099 703173 42123 703229
rect 42179 703173 42193 703229
rect 41863 703166 42193 703173
rect 41863 702585 42193 702592
rect 41713 702529 41883 702585
rect 41939 702529 41963 702585
rect 42019 702529 42043 702585
rect 42099 702529 42123 702585
rect 42179 702529 42193 702585
rect 41863 702522 42193 702529
rect 41863 702033 42193 702040
rect 41713 701977 41883 702033
rect 41939 701977 41963 702033
rect 42019 701977 42043 702033
rect 42099 701977 42123 702033
rect 42179 701977 42193 702033
rect 41863 701970 42193 701977
rect 41863 700193 42193 700200
rect 41713 700137 41883 700193
rect 41939 700137 41963 700193
rect 42019 700137 42043 700193
rect 42099 700137 42123 700193
rect 42179 700137 42193 700193
rect 41863 700130 42193 700137
rect 41863 699549 42193 699556
rect 41713 699493 41883 699549
rect 41939 699493 41963 699549
rect 42019 699493 42043 699549
rect 42099 699493 42123 699549
rect 42179 699493 42193 699549
rect 41863 699486 42193 699493
rect 41863 698905 42193 698912
rect 41713 698849 41883 698905
rect 41939 698849 41963 698905
rect 42019 698849 42043 698905
rect 42099 698849 42123 698905
rect 42179 698849 42193 698905
rect 41863 698842 42193 698849
rect 675407 698351 675737 698358
rect 675407 698295 675427 698351
rect 675483 698295 675507 698351
rect 675563 698295 675587 698351
rect 675643 698295 675667 698351
rect 675723 698295 675887 698351
rect 675407 698288 675737 698295
rect 675407 697707 675737 697714
rect 675407 697651 675427 697707
rect 675483 697651 675507 697707
rect 675563 697651 675587 697707
rect 675643 697651 675667 697707
rect 675723 697651 675887 697707
rect 675407 697644 675737 697651
rect 675407 697063 675737 697070
rect 675407 697007 675427 697063
rect 675483 697007 675507 697063
rect 675563 697007 675587 697063
rect 675643 697007 675667 697063
rect 675723 697007 675887 697063
rect 675407 697000 675737 697007
rect 675407 695223 675737 695230
rect 675407 695167 675427 695223
rect 675483 695167 675507 695223
rect 675563 695167 675587 695223
rect 675643 695167 675667 695223
rect 675723 695167 675887 695223
rect 675407 695160 675737 695167
rect 675407 694671 675737 694678
rect 675407 694615 675427 694671
rect 675483 694615 675507 694671
rect 675563 694615 675587 694671
rect 675643 694615 675667 694671
rect 675723 694615 675887 694671
rect 675407 694608 675737 694615
rect 675407 694027 675737 694034
rect 675407 693971 675427 694027
rect 675483 693971 675507 694027
rect 675563 693971 675587 694027
rect 675643 693971 675667 694027
rect 675723 693971 675887 694027
rect 675407 693964 675737 693971
rect 675407 693383 675737 693390
rect 675407 693327 675427 693383
rect 675483 693327 675507 693383
rect 675563 693327 675587 693383
rect 675643 693327 675667 693383
rect 675723 693327 675887 693383
rect 675407 693320 675737 693327
rect 675407 690899 675737 690906
rect 675407 690843 675427 690899
rect 675483 690843 675507 690899
rect 675563 690843 675587 690899
rect 675643 690843 675667 690899
rect 675723 690843 675887 690899
rect 675407 690836 675737 690843
rect 675407 690347 675737 690354
rect 675407 690291 675427 690347
rect 675483 690291 675507 690347
rect 675563 690291 675587 690347
rect 675643 690291 675667 690347
rect 675723 690291 675887 690347
rect 675407 690284 675737 690291
rect 675407 689703 675737 689710
rect 675407 689647 675427 689703
rect 675483 689647 675507 689703
rect 675563 689647 675587 689703
rect 675643 689647 675667 689703
rect 675723 689647 675887 689703
rect 675407 689640 675737 689647
rect 675407 689059 675737 689066
rect 675407 689003 675427 689059
rect 675483 689003 675507 689059
rect 675563 689003 675587 689059
rect 675643 689003 675667 689059
rect 675723 689003 675887 689059
rect 675407 688996 675737 689003
rect 675407 687863 675737 687870
rect 675407 687807 675427 687863
rect 675483 687807 675507 687863
rect 675563 687807 675587 687863
rect 675643 687807 675667 687863
rect 675723 687807 675887 687863
rect 675407 687800 675737 687807
rect 675407 686667 675737 686674
rect 675407 686611 675427 686667
rect 675483 686611 675507 686667
rect 675563 686611 675587 686667
rect 675643 686611 675667 686667
rect 675723 686611 675887 686667
rect 675407 686604 675737 686611
rect 675407 686023 675737 686030
rect 675407 685967 675427 686023
rect 675483 685967 675507 686023
rect 675563 685967 675587 686023
rect 675643 685967 675667 686023
rect 675723 685967 675887 686023
rect 675407 685960 675737 685967
rect 675407 685379 675737 685386
rect 675407 685323 675427 685379
rect 675483 685323 675507 685379
rect 675563 685323 675587 685379
rect 675643 685323 675667 685379
rect 675723 685323 675887 685379
rect 675407 685316 675737 685323
rect 675407 684183 675737 684190
rect 675407 684127 675427 684183
rect 675483 684127 675507 684183
rect 675563 684127 675587 684183
rect 675643 684127 675667 684183
rect 675723 684127 675887 684183
rect 675407 684120 675737 684127
rect 41863 669873 42193 669880
rect 41713 669817 41883 669873
rect 41939 669817 41963 669873
rect 42019 669817 42043 669873
rect 42099 669817 42123 669873
rect 42179 669817 42193 669873
rect 41863 669810 42193 669817
rect 41863 668677 42193 668684
rect 41713 668621 41883 668677
rect 41939 668621 41963 668677
rect 42019 668621 42043 668677
rect 42099 668621 42123 668677
rect 42179 668621 42193 668677
rect 41863 668614 42193 668621
rect 41863 668033 42193 668040
rect 41713 667977 41883 668033
rect 41939 667977 41963 668033
rect 42019 667977 42043 668033
rect 42099 667977 42123 668033
rect 42179 667977 42193 668033
rect 41863 667970 42193 667977
rect 41863 667389 42193 667396
rect 41713 667333 41883 667389
rect 41939 667333 41963 667389
rect 42019 667333 42043 667389
rect 42099 667333 42123 667389
rect 42179 667333 42193 667389
rect 41863 667326 42193 667333
rect 41863 666193 42193 666200
rect 41713 666137 41883 666193
rect 41939 666137 41963 666193
rect 42019 666137 42043 666193
rect 42099 666137 42123 666193
rect 42179 666137 42193 666193
rect 41863 666130 42193 666137
rect 41863 664997 42193 665004
rect 41713 664941 41883 664997
rect 41939 664941 41963 664997
rect 42019 664941 42043 664997
rect 42099 664941 42123 664997
rect 42179 664941 42193 664997
rect 41863 664934 42193 664941
rect 41863 664353 42193 664360
rect 41713 664297 41883 664353
rect 41939 664297 41963 664353
rect 42019 664297 42043 664353
rect 42099 664297 42123 664353
rect 42179 664297 42193 664353
rect 41863 664290 42193 664297
rect 41863 663709 42193 663716
rect 41713 663653 41883 663709
rect 41939 663653 41963 663709
rect 42019 663653 42043 663709
rect 42099 663653 42123 663709
rect 42179 663653 42193 663709
rect 41863 663646 42193 663653
rect 41863 663157 42193 663164
rect 41713 663101 41883 663157
rect 41939 663101 41963 663157
rect 42019 663101 42043 663157
rect 42099 663101 42123 663157
rect 42179 663101 42193 663157
rect 41863 663094 42193 663101
rect 41863 660673 42193 660680
rect 41713 660617 41883 660673
rect 41939 660617 41963 660673
rect 42019 660617 42043 660673
rect 42099 660617 42123 660673
rect 42179 660617 42193 660673
rect 41863 660610 42193 660617
rect 41863 660029 42193 660036
rect 41713 659973 41883 660029
rect 41939 659973 41963 660029
rect 42019 659973 42043 660029
rect 42099 659973 42123 660029
rect 42179 659973 42193 660029
rect 41863 659966 42193 659973
rect 41863 659385 42193 659392
rect 41713 659329 41883 659385
rect 41939 659329 41963 659385
rect 42019 659329 42043 659385
rect 42099 659329 42123 659385
rect 42179 659329 42193 659385
rect 41863 659322 42193 659329
rect 41863 658833 42193 658840
rect 41713 658777 41883 658833
rect 41939 658777 41963 658833
rect 42019 658777 42043 658833
rect 42099 658777 42123 658833
rect 42179 658777 42193 658833
rect 41863 658770 42193 658777
rect 41863 656993 42193 657000
rect 41713 656937 41883 656993
rect 41939 656937 41963 656993
rect 42019 656937 42043 656993
rect 42099 656937 42123 656993
rect 42179 656937 42193 656993
rect 41863 656930 42193 656937
rect 41863 656349 42193 656356
rect 41713 656293 41883 656349
rect 41939 656293 41963 656349
rect 42019 656293 42043 656349
rect 42099 656293 42123 656349
rect 42179 656293 42193 656349
rect 41863 656286 42193 656293
rect 41863 655705 42193 655712
rect 41713 655649 41883 655705
rect 41939 655649 41963 655705
rect 42019 655649 42043 655705
rect 42099 655649 42123 655705
rect 42179 655649 42193 655705
rect 41863 655642 42193 655649
rect 675407 653151 675737 653158
rect 675407 653095 675427 653151
rect 675483 653095 675507 653151
rect 675563 653095 675587 653151
rect 675643 653095 675667 653151
rect 675723 653095 675887 653151
rect 675407 653088 675737 653095
rect 675407 652507 675737 652514
rect 675407 652451 675427 652507
rect 675483 652451 675507 652507
rect 675563 652451 675587 652507
rect 675643 652451 675667 652507
rect 675723 652451 675887 652507
rect 675407 652444 675737 652451
rect 675407 651863 675737 651870
rect 675407 651807 675427 651863
rect 675483 651807 675507 651863
rect 675563 651807 675587 651863
rect 675643 651807 675667 651863
rect 675723 651807 675887 651863
rect 675407 651800 675737 651807
rect 675407 650023 675737 650030
rect 675407 649967 675427 650023
rect 675483 649967 675507 650023
rect 675563 649967 675587 650023
rect 675643 649967 675667 650023
rect 675723 649967 675887 650023
rect 675407 649960 675737 649967
rect 675407 649471 675737 649478
rect 675407 649415 675427 649471
rect 675483 649415 675507 649471
rect 675563 649415 675587 649471
rect 675643 649415 675667 649471
rect 675723 649415 675887 649471
rect 675407 649408 675737 649415
rect 675407 648827 675737 648834
rect 675407 648771 675427 648827
rect 675483 648771 675507 648827
rect 675563 648771 675587 648827
rect 675643 648771 675667 648827
rect 675723 648771 675887 648827
rect 675407 648764 675737 648771
rect 675407 648183 675737 648190
rect 675407 648127 675427 648183
rect 675483 648127 675507 648183
rect 675563 648127 675587 648183
rect 675643 648127 675667 648183
rect 675723 648127 675887 648183
rect 675407 648120 675737 648127
rect 675407 645699 675737 645706
rect 675407 645643 675427 645699
rect 675483 645643 675507 645699
rect 675563 645643 675587 645699
rect 675643 645643 675667 645699
rect 675723 645643 675887 645699
rect 675407 645636 675737 645643
rect 675407 645147 675737 645154
rect 675407 645091 675427 645147
rect 675483 645091 675507 645147
rect 675563 645091 675587 645147
rect 675643 645091 675667 645147
rect 675723 645091 675887 645147
rect 675407 645084 675737 645091
rect 675407 644503 675737 644510
rect 675407 644447 675427 644503
rect 675483 644447 675507 644503
rect 675563 644447 675587 644503
rect 675643 644447 675667 644503
rect 675723 644447 675887 644503
rect 675407 644440 675737 644447
rect 675407 643859 675737 643866
rect 675407 643803 675427 643859
rect 675483 643803 675507 643859
rect 675563 643803 675587 643859
rect 675643 643803 675667 643859
rect 675723 643803 675887 643859
rect 675407 643796 675737 643803
rect 675407 642663 675737 642670
rect 675407 642607 675427 642663
rect 675483 642607 675507 642663
rect 675563 642607 675587 642663
rect 675643 642607 675667 642663
rect 675723 642607 675887 642663
rect 675407 642600 675737 642607
rect 675407 641467 675737 641474
rect 675407 641411 675427 641467
rect 675483 641411 675507 641467
rect 675563 641411 675587 641467
rect 675643 641411 675667 641467
rect 675723 641411 675887 641467
rect 675407 641404 675737 641411
rect 675407 640823 675737 640830
rect 675407 640767 675427 640823
rect 675483 640767 675507 640823
rect 675563 640767 675587 640823
rect 675643 640767 675667 640823
rect 675723 640767 675887 640823
rect 675407 640760 675737 640767
rect 675407 640179 675737 640186
rect 675407 640123 675427 640179
rect 675483 640123 675507 640179
rect 675563 640123 675587 640179
rect 675643 640123 675667 640179
rect 675723 640123 675887 640179
rect 675407 640116 675737 640123
rect 675407 638983 675737 638990
rect 675407 638927 675427 638983
rect 675483 638927 675507 638983
rect 675563 638927 675587 638983
rect 675643 638927 675667 638983
rect 675723 638927 675887 638983
rect 675407 638920 675737 638927
rect 41863 626673 42193 626680
rect 41713 626617 41883 626673
rect 41939 626617 41963 626673
rect 42019 626617 42043 626673
rect 42099 626617 42123 626673
rect 42179 626617 42193 626673
rect 41863 626610 42193 626617
rect 41863 625477 42193 625484
rect 41713 625421 41883 625477
rect 41939 625421 41963 625477
rect 42019 625421 42043 625477
rect 42099 625421 42123 625477
rect 42179 625421 42193 625477
rect 41863 625414 42193 625421
rect 41863 624833 42193 624840
rect 41713 624777 41883 624833
rect 41939 624777 41963 624833
rect 42019 624777 42043 624833
rect 42099 624777 42123 624833
rect 42179 624777 42193 624833
rect 41863 624770 42193 624777
rect 41863 624189 42193 624196
rect 41713 624133 41883 624189
rect 41939 624133 41963 624189
rect 42019 624133 42043 624189
rect 42099 624133 42123 624189
rect 42179 624133 42193 624189
rect 41863 624126 42193 624133
rect 41863 622993 42193 623000
rect 41713 622937 41883 622993
rect 41939 622937 41963 622993
rect 42019 622937 42043 622993
rect 42099 622937 42123 622993
rect 42179 622937 42193 622993
rect 41863 622930 42193 622937
rect 41863 621797 42193 621804
rect 41713 621741 41883 621797
rect 41939 621741 41963 621797
rect 42019 621741 42043 621797
rect 42099 621741 42123 621797
rect 42179 621741 42193 621797
rect 41863 621734 42193 621741
rect 41863 621153 42193 621160
rect 41713 621097 41883 621153
rect 41939 621097 41963 621153
rect 42019 621097 42043 621153
rect 42099 621097 42123 621153
rect 42179 621097 42193 621153
rect 41863 621090 42193 621097
rect 41863 620509 42193 620516
rect 41713 620453 41883 620509
rect 41939 620453 41963 620509
rect 42019 620453 42043 620509
rect 42099 620453 42123 620509
rect 42179 620453 42193 620509
rect 41863 620446 42193 620453
rect 41863 619957 42193 619964
rect 41713 619901 41883 619957
rect 41939 619901 41963 619957
rect 42019 619901 42043 619957
rect 42099 619901 42123 619957
rect 42179 619901 42193 619957
rect 41863 619894 42193 619901
rect 41863 617473 42193 617480
rect 41713 617417 41883 617473
rect 41939 617417 41963 617473
rect 42019 617417 42043 617473
rect 42099 617417 42123 617473
rect 42179 617417 42193 617473
rect 41863 617410 42193 617417
rect 41863 616829 42193 616836
rect 41713 616773 41883 616829
rect 41939 616773 41963 616829
rect 42019 616773 42043 616829
rect 42099 616773 42123 616829
rect 42179 616773 42193 616829
rect 41863 616766 42193 616773
rect 41863 616185 42193 616192
rect 41713 616129 41883 616185
rect 41939 616129 41963 616185
rect 42019 616129 42043 616185
rect 42099 616129 42123 616185
rect 42179 616129 42193 616185
rect 41863 616122 42193 616129
rect 41863 615633 42193 615640
rect 41713 615577 41883 615633
rect 41939 615577 41963 615633
rect 42019 615577 42043 615633
rect 42099 615577 42123 615633
rect 42179 615577 42193 615633
rect 41863 615570 42193 615577
rect 41863 613793 42193 613800
rect 41713 613737 41883 613793
rect 41939 613737 41963 613793
rect 42019 613737 42043 613793
rect 42099 613737 42123 613793
rect 42179 613737 42193 613793
rect 41863 613730 42193 613737
rect 41863 613149 42193 613156
rect 41713 613093 41883 613149
rect 41939 613093 41963 613149
rect 42019 613093 42043 613149
rect 42099 613093 42123 613149
rect 42179 613093 42193 613149
rect 41863 613086 42193 613093
rect 41863 612505 42193 612512
rect 41713 612449 41883 612505
rect 41939 612449 41963 612505
rect 42019 612449 42043 612505
rect 42099 612449 42123 612505
rect 42179 612449 42193 612505
rect 41863 612442 42193 612449
rect 675407 608151 675737 608158
rect 675407 608095 675427 608151
rect 675483 608095 675507 608151
rect 675563 608095 675587 608151
rect 675643 608095 675667 608151
rect 675723 608095 675887 608151
rect 675407 608088 675737 608095
rect 675407 607507 675737 607514
rect 675407 607451 675427 607507
rect 675483 607451 675507 607507
rect 675563 607451 675587 607507
rect 675643 607451 675667 607507
rect 675723 607451 675887 607507
rect 675407 607444 675737 607451
rect 675407 606863 675737 606870
rect 675407 606807 675427 606863
rect 675483 606807 675507 606863
rect 675563 606807 675587 606863
rect 675643 606807 675667 606863
rect 675723 606807 675887 606863
rect 675407 606800 675737 606807
rect 675407 605023 675737 605030
rect 675407 604967 675427 605023
rect 675483 604967 675507 605023
rect 675563 604967 675587 605023
rect 675643 604967 675667 605023
rect 675723 604967 675887 605023
rect 675407 604960 675737 604967
rect 675407 604471 675737 604478
rect 675407 604415 675427 604471
rect 675483 604415 675507 604471
rect 675563 604415 675587 604471
rect 675643 604415 675667 604471
rect 675723 604415 675887 604471
rect 675407 604408 675737 604415
rect 675407 603827 675737 603834
rect 675407 603771 675427 603827
rect 675483 603771 675507 603827
rect 675563 603771 675587 603827
rect 675643 603771 675667 603827
rect 675723 603771 675887 603827
rect 675407 603764 675737 603771
rect 675407 603183 675737 603190
rect 675407 603127 675427 603183
rect 675483 603127 675507 603183
rect 675563 603127 675587 603183
rect 675643 603127 675667 603183
rect 675723 603127 675887 603183
rect 675407 603120 675737 603127
rect 675407 600699 675737 600706
rect 675407 600643 675427 600699
rect 675483 600643 675507 600699
rect 675563 600643 675587 600699
rect 675643 600643 675667 600699
rect 675723 600643 675887 600699
rect 675407 600636 675737 600643
rect 675407 600147 675737 600154
rect 675407 600091 675427 600147
rect 675483 600091 675507 600147
rect 675563 600091 675587 600147
rect 675643 600091 675667 600147
rect 675723 600091 675887 600147
rect 675407 600084 675737 600091
rect 675407 599503 675737 599510
rect 675407 599447 675427 599503
rect 675483 599447 675507 599503
rect 675563 599447 675587 599503
rect 675643 599447 675667 599503
rect 675723 599447 675887 599503
rect 675407 599440 675737 599447
rect 675407 598859 675737 598866
rect 675407 598803 675427 598859
rect 675483 598803 675507 598859
rect 675563 598803 675587 598859
rect 675643 598803 675667 598859
rect 675723 598803 675887 598859
rect 675407 598796 675737 598803
rect 675407 597663 675737 597670
rect 675407 597607 675427 597663
rect 675483 597607 675507 597663
rect 675563 597607 675587 597663
rect 675643 597607 675667 597663
rect 675723 597607 675887 597663
rect 675407 597600 675737 597607
rect 675407 596467 675737 596474
rect 675407 596411 675427 596467
rect 675483 596411 675507 596467
rect 675563 596411 675587 596467
rect 675643 596411 675667 596467
rect 675723 596411 675887 596467
rect 675407 596404 675737 596411
rect 675407 595823 675737 595830
rect 675407 595767 675427 595823
rect 675483 595767 675507 595823
rect 675563 595767 675587 595823
rect 675643 595767 675667 595823
rect 675723 595767 675887 595823
rect 675407 595760 675737 595767
rect 675407 595179 675737 595186
rect 675407 595123 675427 595179
rect 675483 595123 675507 595179
rect 675563 595123 675587 595179
rect 675643 595123 675667 595179
rect 675723 595123 675887 595179
rect 675407 595116 675737 595123
rect 675407 593983 675737 593990
rect 675407 593927 675427 593983
rect 675483 593927 675507 593983
rect 675563 593927 675587 593983
rect 675643 593927 675667 593983
rect 675723 593927 675887 593983
rect 675407 593920 675737 593927
rect 41863 583473 42193 583480
rect 41713 583417 41883 583473
rect 41939 583417 41963 583473
rect 42019 583417 42043 583473
rect 42099 583417 42123 583473
rect 42179 583417 42193 583473
rect 41863 583410 42193 583417
rect 41863 582277 42193 582284
rect 41713 582221 41883 582277
rect 41939 582221 41963 582277
rect 42019 582221 42043 582277
rect 42099 582221 42123 582277
rect 42179 582221 42193 582277
rect 41863 582214 42193 582221
rect 41863 581633 42193 581640
rect 41713 581577 41883 581633
rect 41939 581577 41963 581633
rect 42019 581577 42043 581633
rect 42099 581577 42123 581633
rect 42179 581577 42193 581633
rect 41863 581570 42193 581577
rect 41863 580989 42193 580996
rect 41713 580933 41883 580989
rect 41939 580933 41963 580989
rect 42019 580933 42043 580989
rect 42099 580933 42123 580989
rect 42179 580933 42193 580989
rect 41863 580926 42193 580933
rect 41863 579793 42193 579800
rect 41713 579737 41883 579793
rect 41939 579737 41963 579793
rect 42019 579737 42043 579793
rect 42099 579737 42123 579793
rect 42179 579737 42193 579793
rect 41863 579730 42193 579737
rect 41863 578597 42193 578604
rect 41713 578541 41883 578597
rect 41939 578541 41963 578597
rect 42019 578541 42043 578597
rect 42099 578541 42123 578597
rect 42179 578541 42193 578597
rect 41863 578534 42193 578541
rect 41863 577953 42193 577960
rect 41713 577897 41883 577953
rect 41939 577897 41963 577953
rect 42019 577897 42043 577953
rect 42099 577897 42123 577953
rect 42179 577897 42193 577953
rect 41863 577890 42193 577897
rect 41863 577309 42193 577316
rect 41713 577253 41883 577309
rect 41939 577253 41963 577309
rect 42019 577253 42043 577309
rect 42099 577253 42123 577309
rect 42179 577253 42193 577309
rect 41863 577246 42193 577253
rect 41863 576757 42193 576764
rect 41713 576701 41883 576757
rect 41939 576701 41963 576757
rect 42019 576701 42043 576757
rect 42099 576701 42123 576757
rect 42179 576701 42193 576757
rect 41863 576694 42193 576701
rect 41863 574273 42193 574280
rect 41713 574217 41883 574273
rect 41939 574217 41963 574273
rect 42019 574217 42043 574273
rect 42099 574217 42123 574273
rect 42179 574217 42193 574273
rect 41863 574210 42193 574217
rect 41863 573629 42193 573636
rect 41713 573573 41883 573629
rect 41939 573573 41963 573629
rect 42019 573573 42043 573629
rect 42099 573573 42123 573629
rect 42179 573573 42193 573629
rect 41863 573566 42193 573573
rect 41863 572985 42193 572992
rect 41713 572929 41883 572985
rect 41939 572929 41963 572985
rect 42019 572929 42043 572985
rect 42099 572929 42123 572985
rect 42179 572929 42193 572985
rect 41863 572922 42193 572929
rect 41863 572433 42193 572440
rect 41713 572377 41883 572433
rect 41939 572377 41963 572433
rect 42019 572377 42043 572433
rect 42099 572377 42123 572433
rect 42179 572377 42193 572433
rect 41863 572370 42193 572377
rect 41863 570593 42193 570600
rect 41713 570537 41883 570593
rect 41939 570537 41963 570593
rect 42019 570537 42043 570593
rect 42099 570537 42123 570593
rect 42179 570537 42193 570593
rect 41863 570530 42193 570537
rect 41863 569949 42193 569956
rect 41713 569893 41883 569949
rect 41939 569893 41963 569949
rect 42019 569893 42043 569949
rect 42099 569893 42123 569949
rect 42179 569893 42193 569949
rect 41863 569886 42193 569893
rect 41863 569305 42193 569312
rect 41713 569249 41883 569305
rect 41939 569249 41963 569305
rect 42019 569249 42043 569305
rect 42099 569249 42123 569305
rect 42179 569249 42193 569305
rect 41863 569242 42193 569249
rect 675407 562951 675737 562958
rect 675407 562895 675427 562951
rect 675483 562895 675507 562951
rect 675563 562895 675587 562951
rect 675643 562895 675667 562951
rect 675723 562895 675887 562951
rect 675407 562888 675737 562895
rect 675407 562307 675737 562314
rect 675407 562251 675427 562307
rect 675483 562251 675507 562307
rect 675563 562251 675587 562307
rect 675643 562251 675667 562307
rect 675723 562251 675887 562307
rect 675407 562244 675737 562251
rect 675407 561663 675737 561670
rect 675407 561607 675427 561663
rect 675483 561607 675507 561663
rect 675563 561607 675587 561663
rect 675643 561607 675667 561663
rect 675723 561607 675887 561663
rect 675407 561600 675737 561607
rect 675407 559823 675737 559830
rect 675407 559767 675427 559823
rect 675483 559767 675507 559823
rect 675563 559767 675587 559823
rect 675643 559767 675667 559823
rect 675723 559767 675887 559823
rect 675407 559760 675737 559767
rect 675407 559271 675737 559278
rect 675407 559215 675427 559271
rect 675483 559215 675507 559271
rect 675563 559215 675587 559271
rect 675643 559215 675667 559271
rect 675723 559215 675887 559271
rect 675407 559208 675737 559215
rect 675407 558627 675737 558634
rect 675407 558571 675427 558627
rect 675483 558571 675507 558627
rect 675563 558571 675587 558627
rect 675643 558571 675667 558627
rect 675723 558571 675887 558627
rect 675407 558564 675737 558571
rect 675407 557983 675737 557990
rect 675407 557927 675427 557983
rect 675483 557927 675507 557983
rect 675563 557927 675587 557983
rect 675643 557927 675667 557983
rect 675723 557927 675887 557983
rect 675407 557920 675737 557927
rect 675407 555499 675737 555506
rect 675407 555443 675427 555499
rect 675483 555443 675507 555499
rect 675563 555443 675587 555499
rect 675643 555443 675667 555499
rect 675723 555443 675887 555499
rect 675407 555436 675737 555443
rect 675407 554947 675737 554954
rect 675407 554891 675427 554947
rect 675483 554891 675507 554947
rect 675563 554891 675587 554947
rect 675643 554891 675667 554947
rect 675723 554891 675887 554947
rect 675407 554884 675737 554891
rect 675407 554303 675737 554310
rect 675407 554247 675427 554303
rect 675483 554247 675507 554303
rect 675563 554247 675587 554303
rect 675643 554247 675667 554303
rect 675723 554247 675887 554303
rect 675407 554240 675737 554247
rect 675407 553659 675737 553666
rect 675407 553603 675427 553659
rect 675483 553603 675507 553659
rect 675563 553603 675587 553659
rect 675643 553603 675667 553659
rect 675723 553603 675887 553659
rect 675407 553596 675737 553603
rect 675407 552463 675737 552470
rect 675407 552407 675427 552463
rect 675483 552407 675507 552463
rect 675563 552407 675587 552463
rect 675643 552407 675667 552463
rect 675723 552407 675887 552463
rect 675407 552400 675737 552407
rect 675407 551267 675737 551274
rect 675407 551211 675427 551267
rect 675483 551211 675507 551267
rect 675563 551211 675587 551267
rect 675643 551211 675667 551267
rect 675723 551211 675887 551267
rect 675407 551204 675737 551211
rect 675407 550623 675737 550630
rect 675407 550567 675427 550623
rect 675483 550567 675507 550623
rect 675563 550567 675587 550623
rect 675643 550567 675667 550623
rect 675723 550567 675887 550623
rect 675407 550560 675737 550567
rect 675407 549979 675737 549986
rect 675407 549923 675427 549979
rect 675483 549923 675507 549979
rect 675563 549923 675587 549979
rect 675643 549923 675667 549979
rect 675723 549923 675887 549979
rect 675407 549916 675737 549923
rect 675407 548783 675737 548790
rect 675407 548727 675427 548783
rect 675483 548727 675507 548783
rect 675563 548727 675587 548783
rect 675643 548727 675667 548783
rect 675723 548727 675887 548783
rect 675407 548720 675737 548727
rect 41863 540273 42193 540280
rect 41713 540217 41883 540273
rect 41939 540217 41963 540273
rect 42019 540217 42043 540273
rect 42099 540217 42123 540273
rect 42179 540217 42193 540273
rect 41863 540210 42193 540217
rect 41863 539077 42193 539084
rect 41713 539021 41883 539077
rect 41939 539021 41963 539077
rect 42019 539021 42043 539077
rect 42099 539021 42123 539077
rect 42179 539021 42193 539077
rect 41863 539014 42193 539021
rect 41863 538433 42193 538440
rect 41713 538377 41883 538433
rect 41939 538377 41963 538433
rect 42019 538377 42043 538433
rect 42099 538377 42123 538433
rect 42179 538377 42193 538433
rect 41863 538370 42193 538377
rect 41863 537789 42193 537796
rect 41713 537733 41883 537789
rect 41939 537733 41963 537789
rect 42019 537733 42043 537789
rect 42099 537733 42123 537789
rect 42179 537733 42193 537789
rect 41863 537726 42193 537733
rect 41863 536593 42193 536600
rect 41713 536537 41883 536593
rect 41939 536537 41963 536593
rect 42019 536537 42043 536593
rect 42099 536537 42123 536593
rect 42179 536537 42193 536593
rect 41863 536530 42193 536537
rect 41863 535397 42193 535404
rect 41713 535341 41883 535397
rect 41939 535341 41963 535397
rect 42019 535341 42043 535397
rect 42099 535341 42123 535397
rect 42179 535341 42193 535397
rect 41863 535334 42193 535341
rect 41863 534753 42193 534760
rect 41713 534697 41883 534753
rect 41939 534697 41963 534753
rect 42019 534697 42043 534753
rect 42099 534697 42123 534753
rect 42179 534697 42193 534753
rect 41863 534690 42193 534697
rect 41863 534109 42193 534116
rect 41713 534053 41883 534109
rect 41939 534053 41963 534109
rect 42019 534053 42043 534109
rect 42099 534053 42123 534109
rect 42179 534053 42193 534109
rect 41863 534046 42193 534053
rect 41863 533557 42193 533564
rect 41713 533501 41883 533557
rect 41939 533501 41963 533557
rect 42019 533501 42043 533557
rect 42099 533501 42123 533557
rect 42179 533501 42193 533557
rect 41863 533494 42193 533501
rect 41863 531073 42193 531080
rect 41713 531017 41883 531073
rect 41939 531017 41963 531073
rect 42019 531017 42043 531073
rect 42099 531017 42123 531073
rect 42179 531017 42193 531073
rect 41863 531010 42193 531017
rect 41863 530429 42193 530436
rect 41713 530373 41883 530429
rect 41939 530373 41963 530429
rect 42019 530373 42043 530429
rect 42099 530373 42123 530429
rect 42179 530373 42193 530429
rect 41863 530366 42193 530373
rect 41863 529785 42193 529792
rect 41713 529729 41883 529785
rect 41939 529729 41963 529785
rect 42019 529729 42043 529785
rect 42099 529729 42123 529785
rect 42179 529729 42193 529785
rect 41863 529722 42193 529729
rect 41863 529233 42193 529240
rect 41713 529177 41883 529233
rect 41939 529177 41963 529233
rect 42019 529177 42043 529233
rect 42099 529177 42123 529233
rect 42179 529177 42193 529233
rect 41863 529170 42193 529177
rect 41863 527393 42193 527400
rect 41713 527337 41883 527393
rect 41939 527337 41963 527393
rect 42019 527337 42043 527393
rect 42099 527337 42123 527393
rect 42179 527337 42193 527393
rect 41863 527330 42193 527337
rect 41863 526749 42193 526756
rect 41713 526693 41883 526749
rect 41939 526693 41963 526749
rect 42019 526693 42043 526749
rect 42099 526693 42123 526749
rect 42179 526693 42193 526749
rect 41863 526686 42193 526693
rect 41863 526105 42193 526112
rect 41713 526049 41883 526105
rect 41939 526049 41963 526105
rect 42019 526049 42043 526105
rect 42099 526049 42123 526105
rect 42179 526049 42193 526105
rect 41863 526042 42193 526049
rect 41863 412673 42193 412680
rect 41713 412617 41883 412673
rect 41939 412617 41963 412673
rect 42019 412617 42043 412673
rect 42099 412617 42123 412673
rect 42179 412617 42193 412673
rect 41863 412610 42193 412617
rect 41863 411477 42193 411484
rect 41713 411421 41883 411477
rect 41939 411421 41963 411477
rect 42019 411421 42043 411477
rect 42099 411421 42123 411477
rect 42179 411421 42193 411477
rect 41863 411414 42193 411421
rect 41863 410833 42193 410840
rect 41713 410777 41883 410833
rect 41939 410777 41963 410833
rect 42019 410777 42043 410833
rect 42099 410777 42123 410833
rect 42179 410777 42193 410833
rect 41863 410770 42193 410777
rect 41863 410189 42193 410196
rect 41713 410133 41883 410189
rect 41939 410133 41963 410189
rect 42019 410133 42043 410189
rect 42099 410133 42123 410189
rect 42179 410133 42193 410189
rect 41863 410126 42193 410133
rect 41863 408993 42193 409000
rect 41713 408937 41883 408993
rect 41939 408937 41963 408993
rect 42019 408937 42043 408993
rect 42099 408937 42123 408993
rect 42179 408937 42193 408993
rect 41863 408930 42193 408937
rect 41863 407797 42193 407804
rect 41713 407741 41883 407797
rect 41939 407741 41963 407797
rect 42019 407741 42043 407797
rect 42099 407741 42123 407797
rect 42179 407741 42193 407797
rect 41863 407734 42193 407741
rect 41863 407153 42193 407160
rect 41713 407097 41883 407153
rect 41939 407097 41963 407153
rect 42019 407097 42043 407153
rect 42099 407097 42123 407153
rect 42179 407097 42193 407153
rect 41863 407090 42193 407097
rect 41863 406509 42193 406516
rect 41713 406453 41883 406509
rect 41939 406453 41963 406509
rect 42019 406453 42043 406509
rect 42099 406453 42123 406509
rect 42179 406453 42193 406509
rect 41863 406446 42193 406453
rect 41863 405957 42193 405964
rect 41713 405901 41883 405957
rect 41939 405901 41963 405957
rect 42019 405901 42043 405957
rect 42099 405901 42123 405957
rect 42179 405901 42193 405957
rect 41863 405894 42193 405901
rect 41863 403473 42193 403480
rect 41713 403417 41883 403473
rect 41939 403417 41963 403473
rect 42019 403417 42043 403473
rect 42099 403417 42123 403473
rect 42179 403417 42193 403473
rect 41863 403410 42193 403417
rect 41863 402829 42193 402836
rect 41713 402773 41883 402829
rect 41939 402773 41963 402829
rect 42019 402773 42043 402829
rect 42099 402773 42123 402829
rect 42179 402773 42193 402829
rect 41863 402766 42193 402773
rect 41863 402185 42193 402192
rect 41713 402129 41883 402185
rect 41939 402129 41963 402185
rect 42019 402129 42043 402185
rect 42099 402129 42123 402185
rect 42179 402129 42193 402185
rect 41863 402122 42193 402129
rect 41863 401633 42193 401640
rect 41713 401577 41883 401633
rect 41939 401577 41963 401633
rect 42019 401577 42043 401633
rect 42099 401577 42123 401633
rect 42179 401577 42193 401633
rect 41863 401570 42193 401577
rect 41863 399793 42193 399800
rect 41713 399737 41883 399793
rect 41939 399737 41963 399793
rect 42019 399737 42043 399793
rect 42099 399737 42123 399793
rect 42179 399737 42193 399793
rect 41863 399730 42193 399737
rect 41863 399149 42193 399156
rect 41713 399093 41883 399149
rect 41939 399093 41963 399149
rect 42019 399093 42043 399149
rect 42099 399093 42123 399149
rect 42179 399093 42193 399149
rect 41863 399086 42193 399093
rect 41863 398505 42193 398512
rect 41713 398449 41883 398505
rect 41939 398449 41963 398505
rect 42019 398449 42043 398505
rect 42099 398449 42123 398505
rect 42179 398449 42193 398505
rect 41863 398442 42193 398449
rect 675407 385751 675737 385758
rect 675407 385695 675427 385751
rect 675483 385695 675507 385751
rect 675563 385695 675587 385751
rect 675643 385695 675667 385751
rect 675723 385695 675887 385751
rect 675407 385688 675737 385695
rect 675407 385107 675737 385114
rect 675407 385051 675427 385107
rect 675483 385051 675507 385107
rect 675563 385051 675587 385107
rect 675643 385051 675667 385107
rect 675723 385051 675887 385107
rect 675407 385044 675737 385051
rect 675407 384463 675737 384470
rect 675407 384407 675427 384463
rect 675483 384407 675507 384463
rect 675563 384407 675587 384463
rect 675643 384407 675667 384463
rect 675723 384407 675887 384463
rect 675407 384400 675737 384407
rect 675407 382623 675737 382630
rect 675407 382567 675427 382623
rect 675483 382567 675507 382623
rect 675563 382567 675587 382623
rect 675643 382567 675667 382623
rect 675723 382567 675887 382623
rect 675407 382560 675737 382567
rect 675407 382071 675737 382078
rect 675407 382015 675427 382071
rect 675483 382015 675507 382071
rect 675563 382015 675587 382071
rect 675643 382015 675667 382071
rect 675723 382015 675887 382071
rect 675407 382008 675737 382015
rect 675407 381427 675737 381434
rect 675407 381371 675427 381427
rect 675483 381371 675507 381427
rect 675563 381371 675587 381427
rect 675643 381371 675667 381427
rect 675723 381371 675887 381427
rect 675407 381364 675737 381371
rect 675407 380783 675737 380790
rect 675407 380727 675427 380783
rect 675483 380727 675507 380783
rect 675563 380727 675587 380783
rect 675643 380727 675667 380783
rect 675723 380727 675887 380783
rect 675407 380720 675737 380727
rect 675407 378299 675737 378306
rect 675407 378243 675427 378299
rect 675483 378243 675507 378299
rect 675563 378243 675587 378299
rect 675643 378243 675667 378299
rect 675723 378243 675887 378299
rect 675407 378236 675737 378243
rect 675407 377747 675737 377754
rect 675407 377691 675427 377747
rect 675483 377691 675507 377747
rect 675563 377691 675587 377747
rect 675643 377691 675667 377747
rect 675723 377691 675887 377747
rect 675407 377684 675737 377691
rect 675407 377103 675737 377110
rect 675407 377047 675427 377103
rect 675483 377047 675507 377103
rect 675563 377047 675587 377103
rect 675643 377047 675667 377103
rect 675723 377047 675887 377103
rect 675407 377040 675737 377047
rect 675407 376459 675737 376466
rect 675407 376403 675427 376459
rect 675483 376403 675507 376459
rect 675563 376403 675587 376459
rect 675643 376403 675667 376459
rect 675723 376403 675887 376459
rect 675407 376396 675737 376403
rect 675407 375263 675737 375270
rect 675407 375207 675427 375263
rect 675483 375207 675507 375263
rect 675563 375207 675587 375263
rect 675643 375207 675667 375263
rect 675723 375207 675887 375263
rect 675407 375200 675737 375207
rect 675407 373423 675737 373430
rect 675407 373367 675427 373423
rect 675483 373367 675507 373423
rect 675563 373367 675587 373423
rect 675643 373367 675667 373423
rect 675723 373367 675887 373423
rect 675407 373360 675737 373367
rect 675407 372779 675737 372786
rect 675407 372723 675427 372779
rect 675483 372723 675507 372779
rect 675563 372723 675587 372779
rect 675643 372723 675667 372779
rect 675723 372723 675887 372779
rect 675407 372716 675737 372723
rect 675407 371583 675737 371590
rect 675407 371527 675427 371583
rect 675483 371527 675507 371583
rect 675563 371527 675587 371583
rect 675643 371527 675667 371583
rect 675723 371527 675887 371583
rect 675407 371520 675737 371527
rect 41863 369473 42193 369480
rect 41713 369417 41883 369473
rect 41939 369417 41963 369473
rect 42019 369417 42043 369473
rect 42099 369417 42123 369473
rect 42179 369417 42193 369473
rect 41863 369410 42193 369417
rect 41863 368277 42193 368284
rect 41713 368221 41883 368277
rect 41939 368221 41963 368277
rect 42019 368221 42043 368277
rect 42099 368221 42123 368277
rect 42179 368221 42193 368277
rect 41863 368214 42193 368221
rect 41863 367633 42193 367640
rect 41713 367577 41883 367633
rect 41939 367577 41963 367633
rect 42019 367577 42043 367633
rect 42099 367577 42123 367633
rect 42179 367577 42193 367633
rect 41863 367570 42193 367577
rect 41863 366989 42193 366996
rect 41713 366933 41883 366989
rect 41939 366933 41963 366989
rect 42019 366933 42043 366989
rect 42099 366933 42123 366989
rect 42179 366933 42193 366989
rect 41863 366926 42193 366933
rect 41863 365793 42193 365800
rect 41713 365737 41883 365793
rect 41939 365737 41963 365793
rect 42019 365737 42043 365793
rect 42099 365737 42123 365793
rect 42179 365737 42193 365793
rect 41863 365730 42193 365737
rect 41863 364597 42193 364604
rect 41713 364541 41883 364597
rect 41939 364541 41963 364597
rect 42019 364541 42043 364597
rect 42099 364541 42123 364597
rect 42179 364541 42193 364597
rect 41863 364534 42193 364541
rect 41863 363953 42193 363960
rect 41713 363897 41883 363953
rect 41939 363897 41963 363953
rect 42019 363897 42043 363953
rect 42099 363897 42123 363953
rect 42179 363897 42193 363953
rect 41863 363890 42193 363897
rect 41863 363309 42193 363316
rect 41713 363253 41883 363309
rect 41939 363253 41963 363309
rect 42019 363253 42043 363309
rect 42099 363253 42123 363309
rect 42179 363253 42193 363309
rect 41863 363246 42193 363253
rect 41863 362757 42193 362764
rect 41713 362701 41883 362757
rect 41939 362701 41963 362757
rect 42019 362701 42043 362757
rect 42099 362701 42123 362757
rect 42179 362701 42193 362757
rect 41863 362694 42193 362701
rect 41863 360273 42193 360280
rect 41713 360217 41883 360273
rect 41939 360217 41963 360273
rect 42019 360217 42043 360273
rect 42099 360217 42123 360273
rect 42179 360217 42193 360273
rect 41863 360210 42193 360217
rect 41863 359629 42193 359636
rect 41713 359573 41883 359629
rect 41939 359573 41963 359629
rect 42019 359573 42043 359629
rect 42099 359573 42123 359629
rect 42179 359573 42193 359629
rect 41863 359566 42193 359573
rect 41863 358985 42193 358992
rect 41713 358929 41883 358985
rect 41939 358929 41963 358985
rect 42019 358929 42043 358985
rect 42099 358929 42123 358985
rect 42179 358929 42193 358985
rect 41863 358922 42193 358929
rect 41863 358433 42193 358440
rect 41713 358377 41883 358433
rect 41939 358377 41963 358433
rect 42019 358377 42043 358433
rect 42099 358377 42123 358433
rect 42179 358377 42193 358433
rect 41863 358370 42193 358377
rect 41863 356593 42193 356600
rect 41713 356537 41883 356593
rect 41939 356537 41963 356593
rect 42019 356537 42043 356593
rect 42099 356537 42123 356593
rect 42179 356537 42193 356593
rect 41863 356530 42193 356537
rect 41863 355949 42193 355956
rect 41713 355893 41883 355949
rect 41939 355893 41963 355949
rect 42019 355893 42043 355949
rect 42099 355893 42123 355949
rect 42179 355893 42193 355949
rect 41863 355886 42193 355893
rect 41863 355305 42193 355312
rect 41713 355249 41883 355305
rect 41939 355249 41963 355305
rect 42019 355249 42043 355305
rect 42099 355249 42123 355305
rect 42179 355249 42193 355305
rect 41863 355242 42193 355249
rect 675407 340551 675737 340558
rect 675407 340495 675427 340551
rect 675483 340495 675507 340551
rect 675563 340495 675587 340551
rect 675643 340495 675667 340551
rect 675723 340495 675887 340551
rect 675407 340488 675737 340495
rect 675407 339907 675737 339914
rect 675407 339851 675427 339907
rect 675483 339851 675507 339907
rect 675563 339851 675587 339907
rect 675643 339851 675667 339907
rect 675723 339851 675887 339907
rect 675407 339844 675737 339851
rect 675407 339263 675737 339270
rect 675407 339207 675427 339263
rect 675483 339207 675507 339263
rect 675563 339207 675587 339263
rect 675643 339207 675667 339263
rect 675723 339207 675887 339263
rect 675407 339200 675737 339207
rect 675407 337423 675737 337430
rect 675407 337367 675427 337423
rect 675483 337367 675507 337423
rect 675563 337367 675587 337423
rect 675643 337367 675667 337423
rect 675723 337367 675887 337423
rect 675407 337360 675737 337367
rect 675407 336871 675737 336878
rect 675407 336815 675427 336871
rect 675483 336815 675507 336871
rect 675563 336815 675587 336871
rect 675643 336815 675667 336871
rect 675723 336815 675887 336871
rect 675407 336808 675737 336815
rect 675407 336227 675737 336234
rect 675407 336171 675427 336227
rect 675483 336171 675507 336227
rect 675563 336171 675587 336227
rect 675643 336171 675667 336227
rect 675723 336171 675887 336227
rect 675407 336164 675737 336171
rect 675407 335583 675737 335590
rect 675407 335527 675427 335583
rect 675483 335527 675507 335583
rect 675563 335527 675587 335583
rect 675643 335527 675667 335583
rect 675723 335527 675887 335583
rect 675407 335520 675737 335527
rect 675407 333099 675737 333106
rect 675407 333043 675427 333099
rect 675483 333043 675507 333099
rect 675563 333043 675587 333099
rect 675643 333043 675667 333099
rect 675723 333043 675887 333099
rect 675407 333036 675737 333043
rect 675407 332547 675737 332554
rect 675407 332491 675427 332547
rect 675483 332491 675507 332547
rect 675563 332491 675587 332547
rect 675643 332491 675667 332547
rect 675723 332491 675887 332547
rect 675407 332484 675737 332491
rect 675407 331903 675737 331910
rect 675407 331847 675427 331903
rect 675483 331847 675507 331903
rect 675563 331847 675587 331903
rect 675643 331847 675667 331903
rect 675723 331847 675887 331903
rect 675407 331840 675737 331847
rect 675407 331259 675737 331266
rect 675407 331203 675427 331259
rect 675483 331203 675507 331259
rect 675563 331203 675587 331259
rect 675643 331203 675667 331259
rect 675723 331203 675887 331259
rect 675407 331196 675737 331203
rect 675407 330063 675737 330070
rect 675407 330007 675427 330063
rect 675483 330007 675507 330063
rect 675563 330007 675587 330063
rect 675643 330007 675667 330063
rect 675723 330007 675887 330063
rect 675407 330000 675737 330007
rect 675407 328223 675737 328230
rect 675407 328167 675427 328223
rect 675483 328167 675507 328223
rect 675563 328167 675587 328223
rect 675643 328167 675667 328223
rect 675723 328167 675887 328223
rect 675407 328160 675737 328167
rect 675407 327579 675737 327586
rect 675407 327523 675427 327579
rect 675483 327523 675507 327579
rect 675563 327523 675587 327579
rect 675643 327523 675667 327579
rect 675723 327523 675887 327579
rect 675407 327516 675737 327523
rect 675407 326383 675737 326390
rect 675407 326327 675427 326383
rect 675483 326327 675507 326383
rect 675563 326327 675587 326383
rect 675643 326327 675667 326383
rect 675723 326327 675887 326383
rect 675407 326320 675737 326327
rect 41863 326273 42193 326280
rect 41713 326217 41883 326273
rect 41939 326217 41963 326273
rect 42019 326217 42043 326273
rect 42099 326217 42123 326273
rect 42179 326217 42193 326273
rect 41863 326210 42193 326217
rect 41863 325077 42193 325084
rect 41713 325021 41883 325077
rect 41939 325021 41963 325077
rect 42019 325021 42043 325077
rect 42099 325021 42123 325077
rect 42179 325021 42193 325077
rect 41863 325014 42193 325021
rect 41863 324433 42193 324440
rect 41713 324377 41883 324433
rect 41939 324377 41963 324433
rect 42019 324377 42043 324433
rect 42099 324377 42123 324433
rect 42179 324377 42193 324433
rect 41863 324370 42193 324377
rect 41863 323789 42193 323796
rect 41713 323733 41883 323789
rect 41939 323733 41963 323789
rect 42019 323733 42043 323789
rect 42099 323733 42123 323789
rect 42179 323733 42193 323789
rect 41863 323726 42193 323733
rect 41863 322593 42193 322600
rect 41713 322537 41883 322593
rect 41939 322537 41963 322593
rect 42019 322537 42043 322593
rect 42099 322537 42123 322593
rect 42179 322537 42193 322593
rect 41863 322530 42193 322537
rect 41863 321397 42193 321404
rect 41713 321341 41883 321397
rect 41939 321341 41963 321397
rect 42019 321341 42043 321397
rect 42099 321341 42123 321397
rect 42179 321341 42193 321397
rect 41863 321334 42193 321341
rect 41863 320753 42193 320760
rect 41713 320697 41883 320753
rect 41939 320697 41963 320753
rect 42019 320697 42043 320753
rect 42099 320697 42123 320753
rect 42179 320697 42193 320753
rect 41863 320690 42193 320697
rect 41863 320109 42193 320116
rect 41713 320053 41883 320109
rect 41939 320053 41963 320109
rect 42019 320053 42043 320109
rect 42099 320053 42123 320109
rect 42179 320053 42193 320109
rect 41863 320046 42193 320053
rect 41863 319557 42193 319564
rect 41713 319501 41883 319557
rect 41939 319501 41963 319557
rect 42019 319501 42043 319557
rect 42099 319501 42123 319557
rect 42179 319501 42193 319557
rect 41863 319494 42193 319501
rect 41863 317073 42193 317080
rect 41713 317017 41883 317073
rect 41939 317017 41963 317073
rect 42019 317017 42043 317073
rect 42099 317017 42123 317073
rect 42179 317017 42193 317073
rect 41863 317010 42193 317017
rect 41863 316429 42193 316436
rect 41713 316373 41883 316429
rect 41939 316373 41963 316429
rect 42019 316373 42043 316429
rect 42099 316373 42123 316429
rect 42179 316373 42193 316429
rect 41863 316366 42193 316373
rect 41863 315785 42193 315792
rect 41713 315729 41883 315785
rect 41939 315729 41963 315785
rect 42019 315729 42043 315785
rect 42099 315729 42123 315785
rect 42179 315729 42193 315785
rect 41863 315722 42193 315729
rect 41863 315233 42193 315240
rect 41713 315177 41883 315233
rect 41939 315177 41963 315233
rect 42019 315177 42043 315233
rect 42099 315177 42123 315233
rect 42179 315177 42193 315233
rect 41863 315170 42193 315177
rect 41863 313393 42193 313400
rect 41713 313337 41883 313393
rect 41939 313337 41963 313393
rect 42019 313337 42043 313393
rect 42099 313337 42123 313393
rect 42179 313337 42193 313393
rect 41863 313330 42193 313337
rect 41863 312749 42193 312756
rect 41713 312693 41883 312749
rect 41939 312693 41963 312749
rect 42019 312693 42043 312749
rect 42099 312693 42123 312749
rect 42179 312693 42193 312749
rect 41863 312686 42193 312693
rect 41863 312105 42193 312112
rect 41713 312049 41883 312105
rect 41939 312049 41963 312105
rect 42019 312049 42043 312105
rect 42099 312049 42123 312105
rect 42179 312049 42193 312105
rect 41863 312042 42193 312049
rect 675407 295551 675737 295558
rect 675407 295495 675427 295551
rect 675483 295495 675507 295551
rect 675563 295495 675587 295551
rect 675643 295495 675667 295551
rect 675723 295495 675887 295551
rect 675407 295488 675737 295495
rect 675407 294907 675737 294914
rect 675407 294851 675427 294907
rect 675483 294851 675507 294907
rect 675563 294851 675587 294907
rect 675643 294851 675667 294907
rect 675723 294851 675887 294907
rect 675407 294844 675737 294851
rect 675407 294263 675737 294270
rect 675407 294207 675427 294263
rect 675483 294207 675507 294263
rect 675563 294207 675587 294263
rect 675643 294207 675667 294263
rect 675723 294207 675887 294263
rect 675407 294200 675737 294207
rect 675407 292423 675737 292430
rect 675407 292367 675427 292423
rect 675483 292367 675507 292423
rect 675563 292367 675587 292423
rect 675643 292367 675667 292423
rect 675723 292367 675887 292423
rect 675407 292360 675737 292367
rect 675407 291871 675737 291878
rect 675407 291815 675427 291871
rect 675483 291815 675507 291871
rect 675563 291815 675587 291871
rect 675643 291815 675667 291871
rect 675723 291815 675887 291871
rect 675407 291808 675737 291815
rect 675407 291227 675737 291234
rect 675407 291171 675427 291227
rect 675483 291171 675507 291227
rect 675563 291171 675587 291227
rect 675643 291171 675667 291227
rect 675723 291171 675887 291227
rect 675407 291164 675737 291171
rect 675407 290583 675737 290590
rect 675407 290527 675427 290583
rect 675483 290527 675507 290583
rect 675563 290527 675587 290583
rect 675643 290527 675667 290583
rect 675723 290527 675887 290583
rect 675407 290520 675737 290527
rect 675407 288099 675737 288106
rect 675407 288043 675427 288099
rect 675483 288043 675507 288099
rect 675563 288043 675587 288099
rect 675643 288043 675667 288099
rect 675723 288043 675887 288099
rect 675407 288036 675737 288043
rect 675407 287547 675737 287554
rect 675407 287491 675427 287547
rect 675483 287491 675507 287547
rect 675563 287491 675587 287547
rect 675643 287491 675667 287547
rect 675723 287491 675887 287547
rect 675407 287484 675737 287491
rect 675407 286903 675737 286910
rect 675407 286847 675427 286903
rect 675483 286847 675507 286903
rect 675563 286847 675587 286903
rect 675643 286847 675667 286903
rect 675723 286847 675887 286903
rect 675407 286840 675737 286847
rect 675407 286259 675737 286266
rect 675407 286203 675427 286259
rect 675483 286203 675507 286259
rect 675563 286203 675587 286259
rect 675643 286203 675667 286259
rect 675723 286203 675887 286259
rect 675407 286196 675737 286203
rect 675407 285063 675737 285070
rect 675407 285007 675427 285063
rect 675483 285007 675507 285063
rect 675563 285007 675587 285063
rect 675643 285007 675667 285063
rect 675723 285007 675887 285063
rect 675407 285000 675737 285007
rect 675407 283223 675737 283230
rect 675407 283167 675427 283223
rect 675483 283167 675507 283223
rect 675563 283167 675587 283223
rect 675643 283167 675667 283223
rect 675723 283167 675887 283223
rect 675407 283160 675737 283167
rect 41863 283073 42193 283080
rect 41713 283017 41883 283073
rect 41939 283017 41963 283073
rect 42019 283017 42043 283073
rect 42099 283017 42123 283073
rect 42179 283017 42193 283073
rect 41863 283010 42193 283017
rect 675407 282579 675737 282586
rect 675407 282523 675427 282579
rect 675483 282523 675507 282579
rect 675563 282523 675587 282579
rect 675643 282523 675667 282579
rect 675723 282523 675887 282579
rect 675407 282516 675737 282523
rect 41863 281877 42193 281884
rect 41713 281821 41883 281877
rect 41939 281821 41963 281877
rect 42019 281821 42043 281877
rect 42099 281821 42123 281877
rect 42179 281821 42193 281877
rect 41863 281814 42193 281821
rect 675407 281383 675737 281390
rect 675407 281327 675427 281383
rect 675483 281327 675507 281383
rect 675563 281327 675587 281383
rect 675643 281327 675667 281383
rect 675723 281327 675887 281383
rect 675407 281320 675737 281327
rect 41863 281233 42193 281240
rect 41713 281177 41883 281233
rect 41939 281177 41963 281233
rect 42019 281177 42043 281233
rect 42099 281177 42123 281233
rect 42179 281177 42193 281233
rect 41863 281170 42193 281177
rect 41863 280589 42193 280596
rect 41713 280533 41883 280589
rect 41939 280533 41963 280589
rect 42019 280533 42043 280589
rect 42099 280533 42123 280589
rect 42179 280533 42193 280589
rect 41863 280526 42193 280533
rect 41863 279393 42193 279400
rect 41713 279337 41883 279393
rect 41939 279337 41963 279393
rect 42019 279337 42043 279393
rect 42099 279337 42123 279393
rect 42179 279337 42193 279393
rect 41863 279330 42193 279337
rect 41863 278197 42193 278204
rect 41713 278141 41883 278197
rect 41939 278141 41963 278197
rect 42019 278141 42043 278197
rect 42099 278141 42123 278197
rect 42179 278141 42193 278197
rect 41863 278134 42193 278141
rect 41863 277553 42193 277560
rect 41713 277497 41883 277553
rect 41939 277497 41963 277553
rect 42019 277497 42043 277553
rect 42099 277497 42123 277553
rect 42179 277497 42193 277553
rect 41863 277490 42193 277497
rect 41863 276909 42193 276916
rect 41713 276853 41883 276909
rect 41939 276853 41963 276909
rect 42019 276853 42043 276909
rect 42099 276853 42123 276909
rect 42179 276853 42193 276909
rect 41863 276846 42193 276853
rect 41863 276357 42193 276364
rect 41713 276301 41883 276357
rect 41939 276301 41963 276357
rect 42019 276301 42043 276357
rect 42099 276301 42123 276357
rect 42179 276301 42193 276357
rect 41863 276294 42193 276301
rect 41863 273873 42193 273880
rect 41713 273817 41883 273873
rect 41939 273817 41963 273873
rect 42019 273817 42043 273873
rect 42099 273817 42123 273873
rect 42179 273817 42193 273873
rect 41863 273810 42193 273817
rect 41863 273229 42193 273236
rect 41713 273173 41883 273229
rect 41939 273173 41963 273229
rect 42019 273173 42043 273229
rect 42099 273173 42123 273229
rect 42179 273173 42193 273229
rect 41863 273166 42193 273173
rect 41863 272585 42193 272592
rect 41713 272529 41883 272585
rect 41939 272529 41963 272585
rect 42019 272529 42043 272585
rect 42099 272529 42123 272585
rect 42179 272529 42193 272585
rect 41863 272522 42193 272529
rect 41863 272033 42193 272040
rect 41713 271977 41883 272033
rect 41939 271977 41963 272033
rect 42019 271977 42043 272033
rect 42099 271977 42123 272033
rect 42179 271977 42193 272033
rect 41863 271970 42193 271977
rect 41863 270193 42193 270200
rect 41713 270137 41883 270193
rect 41939 270137 41963 270193
rect 42019 270137 42043 270193
rect 42099 270137 42123 270193
rect 42179 270137 42193 270193
rect 41863 270130 42193 270137
rect 41863 269549 42193 269556
rect 41713 269493 41883 269549
rect 41939 269493 41963 269549
rect 42019 269493 42043 269549
rect 42099 269493 42123 269549
rect 42179 269493 42193 269549
rect 41863 269486 42193 269493
rect 41863 268905 42193 268912
rect 41713 268849 41883 268905
rect 41939 268849 41963 268905
rect 42019 268849 42043 268905
rect 42099 268849 42123 268905
rect 42179 268849 42193 268905
rect 41863 268842 42193 268849
rect 675407 250551 675737 250558
rect 675407 250495 675427 250551
rect 675483 250495 675507 250551
rect 675563 250495 675587 250551
rect 675643 250495 675667 250551
rect 675723 250495 675887 250551
rect 675407 250488 675737 250495
rect 675407 249907 675737 249914
rect 675407 249851 675427 249907
rect 675483 249851 675507 249907
rect 675563 249851 675587 249907
rect 675643 249851 675667 249907
rect 675723 249851 675887 249907
rect 675407 249844 675737 249851
rect 675407 249263 675737 249270
rect 675407 249207 675427 249263
rect 675483 249207 675507 249263
rect 675563 249207 675587 249263
rect 675643 249207 675667 249263
rect 675723 249207 675887 249263
rect 675407 249200 675737 249207
rect 675407 247423 675737 247430
rect 675407 247367 675427 247423
rect 675483 247367 675507 247423
rect 675563 247367 675587 247423
rect 675643 247367 675667 247423
rect 675723 247367 675887 247423
rect 675407 247360 675737 247367
rect 675407 246871 675737 246878
rect 675407 246815 675427 246871
rect 675483 246815 675507 246871
rect 675563 246815 675587 246871
rect 675643 246815 675667 246871
rect 675723 246815 675887 246871
rect 675407 246808 675737 246815
rect 675407 246227 675737 246234
rect 675407 246171 675427 246227
rect 675483 246171 675507 246227
rect 675563 246171 675587 246227
rect 675643 246171 675667 246227
rect 675723 246171 675887 246227
rect 675407 246164 675737 246171
rect 675407 245583 675737 245590
rect 675407 245527 675427 245583
rect 675483 245527 675507 245583
rect 675563 245527 675587 245583
rect 675643 245527 675667 245583
rect 675723 245527 675887 245583
rect 675407 245520 675737 245527
rect 675407 243099 675737 243106
rect 675407 243043 675427 243099
rect 675483 243043 675507 243099
rect 675563 243043 675587 243099
rect 675643 243043 675667 243099
rect 675723 243043 675887 243099
rect 675407 243036 675737 243043
rect 675407 242547 675737 242554
rect 675407 242491 675427 242547
rect 675483 242491 675507 242547
rect 675563 242491 675587 242547
rect 675643 242491 675667 242547
rect 675723 242491 675887 242547
rect 675407 242484 675737 242491
rect 675407 241903 675737 241910
rect 675407 241847 675427 241903
rect 675483 241847 675507 241903
rect 675563 241847 675587 241903
rect 675643 241847 675667 241903
rect 675723 241847 675887 241903
rect 675407 241840 675737 241847
rect 675407 241259 675737 241266
rect 675407 241203 675427 241259
rect 675483 241203 675507 241259
rect 675563 241203 675587 241259
rect 675643 241203 675667 241259
rect 675723 241203 675887 241259
rect 675407 241196 675737 241203
rect 675407 240063 675737 240070
rect 675407 240007 675427 240063
rect 675483 240007 675507 240063
rect 675563 240007 675587 240063
rect 675643 240007 675667 240063
rect 675723 240007 675887 240063
rect 675407 240000 675737 240007
rect 41863 239873 42193 239880
rect 41713 239817 41883 239873
rect 41939 239817 41963 239873
rect 42019 239817 42043 239873
rect 42099 239817 42123 239873
rect 42179 239817 42193 239873
rect 41863 239810 42193 239817
rect 41863 238677 42193 238684
rect 41713 238621 41883 238677
rect 41939 238621 41963 238677
rect 42019 238621 42043 238677
rect 42099 238621 42123 238677
rect 42179 238621 42193 238677
rect 41863 238614 42193 238621
rect 675407 238223 675737 238230
rect 675407 238167 675427 238223
rect 675483 238167 675507 238223
rect 675563 238167 675587 238223
rect 675643 238167 675667 238223
rect 675723 238167 675887 238223
rect 675407 238160 675737 238167
rect 41863 238033 42193 238040
rect 41713 237977 41883 238033
rect 41939 237977 41963 238033
rect 42019 237977 42043 238033
rect 42099 237977 42123 238033
rect 42179 237977 42193 238033
rect 41863 237970 42193 237977
rect 675407 237579 675737 237586
rect 675407 237523 675427 237579
rect 675483 237523 675507 237579
rect 675563 237523 675587 237579
rect 675643 237523 675667 237579
rect 675723 237523 675887 237579
rect 675407 237516 675737 237523
rect 675407 236383 675737 236390
rect 675407 236327 675427 236383
rect 675483 236327 675507 236383
rect 675563 236327 675587 236383
rect 675643 236327 675667 236383
rect 675723 236327 675887 236383
rect 675407 236320 675737 236327
rect 41863 236193 42193 236200
rect 41713 236137 41883 236193
rect 41939 236137 41963 236193
rect 42019 236137 42043 236193
rect 42099 236137 42123 236193
rect 42179 236137 42193 236193
rect 41863 236130 42193 236137
rect 41863 234997 42193 235004
rect 41713 234941 41883 234997
rect 41939 234941 41963 234997
rect 42019 234941 42043 234997
rect 42099 234941 42123 234997
rect 42179 234941 42193 234997
rect 41863 234934 42193 234941
rect 41863 234353 42193 234360
rect 41713 234297 41883 234353
rect 41939 234297 41963 234353
rect 42019 234297 42043 234353
rect 42099 234297 42123 234353
rect 42179 234297 42193 234353
rect 41863 234290 42193 234297
rect 41863 233709 42193 233716
rect 41713 233653 41883 233709
rect 41939 233653 41963 233709
rect 42019 233653 42043 233709
rect 42099 233653 42123 233709
rect 42179 233653 42193 233709
rect 41863 233646 42193 233653
rect 41863 233157 42193 233164
rect 41713 233101 41883 233157
rect 41939 233101 41963 233157
rect 42019 233101 42043 233157
rect 42099 233101 42123 233157
rect 42179 233101 42193 233157
rect 41863 233094 42193 233101
rect 41863 230673 42193 230680
rect 41713 230617 41883 230673
rect 41939 230617 41963 230673
rect 42019 230617 42043 230673
rect 42099 230617 42123 230673
rect 42179 230617 42193 230673
rect 41863 230610 42193 230617
rect 41863 230029 42193 230036
rect 41713 229973 41883 230029
rect 41939 229973 41963 230029
rect 42019 229973 42043 230029
rect 42099 229973 42123 230029
rect 42179 229973 42193 230029
rect 41863 229966 42193 229973
rect 41863 229385 42193 229392
rect 41713 229329 41883 229385
rect 41939 229329 41963 229385
rect 42019 229329 42043 229385
rect 42099 229329 42123 229385
rect 42179 229329 42193 229385
rect 41863 229322 42193 229329
rect 41863 228833 42193 228840
rect 41713 228777 41883 228833
rect 41939 228777 41963 228833
rect 42019 228777 42043 228833
rect 42099 228777 42123 228833
rect 42179 228777 42193 228833
rect 41863 228770 42193 228777
rect 41863 226993 42193 227000
rect 41713 226937 41883 226993
rect 41939 226937 41963 226993
rect 42019 226937 42043 226993
rect 42099 226937 42123 226993
rect 42179 226937 42193 226993
rect 41863 226930 42193 226937
rect 41863 226349 42193 226356
rect 41713 226293 41883 226349
rect 41939 226293 41963 226349
rect 42019 226293 42043 226349
rect 42099 226293 42123 226349
rect 42179 226293 42193 226349
rect 41863 226286 42193 226293
rect 41863 225705 42193 225712
rect 41713 225649 41883 225705
rect 41939 225649 41963 225705
rect 42019 225649 42043 225705
rect 42099 225649 42123 225705
rect 42179 225649 42193 225705
rect 41863 225642 42193 225649
rect 675407 205351 675737 205358
rect 675407 205295 675427 205351
rect 675483 205295 675507 205351
rect 675563 205295 675587 205351
rect 675643 205295 675667 205351
rect 675723 205295 675887 205351
rect 675407 205288 675737 205295
rect 675407 204707 675737 204714
rect 675407 204651 675427 204707
rect 675483 204651 675507 204707
rect 675563 204651 675587 204707
rect 675643 204651 675667 204707
rect 675723 204651 675887 204707
rect 675407 204644 675737 204651
rect 675407 204063 675737 204070
rect 675407 204007 675427 204063
rect 675483 204007 675507 204063
rect 675563 204007 675587 204063
rect 675643 204007 675667 204063
rect 675723 204007 675887 204063
rect 675407 204000 675737 204007
rect 675407 202223 675737 202230
rect 675407 202167 675427 202223
rect 675483 202167 675507 202223
rect 675563 202167 675587 202223
rect 675643 202167 675667 202223
rect 675723 202167 675887 202223
rect 675407 202160 675737 202167
rect 675407 201671 675737 201678
rect 675407 201615 675427 201671
rect 675483 201615 675507 201671
rect 675563 201615 675587 201671
rect 675643 201615 675667 201671
rect 675723 201615 675887 201671
rect 675407 201608 675737 201615
rect 675407 201027 675737 201034
rect 675407 200971 675427 201027
rect 675483 200971 675507 201027
rect 675563 200971 675587 201027
rect 675643 200971 675667 201027
rect 675723 200971 675887 201027
rect 675407 200964 675737 200971
rect 675407 200383 675737 200390
rect 675407 200327 675427 200383
rect 675483 200327 675507 200383
rect 675563 200327 675587 200383
rect 675643 200327 675667 200383
rect 675723 200327 675887 200383
rect 675407 200320 675737 200327
rect 675407 197899 675737 197906
rect 675407 197843 675427 197899
rect 675483 197843 675507 197899
rect 675563 197843 675587 197899
rect 675643 197843 675667 197899
rect 675723 197843 675887 197899
rect 675407 197836 675737 197843
rect 675407 197347 675737 197354
rect 675407 197291 675427 197347
rect 675483 197291 675507 197347
rect 675563 197291 675587 197347
rect 675643 197291 675667 197347
rect 675723 197291 675887 197347
rect 675407 197284 675737 197291
rect 675407 196703 675737 196710
rect 41863 196673 42193 196680
rect 41713 196617 41883 196673
rect 41939 196617 41963 196673
rect 42019 196617 42043 196673
rect 42099 196617 42123 196673
rect 42179 196617 42193 196673
rect 675407 196647 675427 196703
rect 675483 196647 675507 196703
rect 675563 196647 675587 196703
rect 675643 196647 675667 196703
rect 675723 196647 675887 196703
rect 675407 196640 675737 196647
rect 41863 196610 42193 196617
rect 675407 196059 675737 196066
rect 675407 196003 675427 196059
rect 675483 196003 675507 196059
rect 675563 196003 675587 196059
rect 675643 196003 675667 196059
rect 675723 196003 675887 196059
rect 675407 195996 675737 196003
rect 41863 195477 42193 195484
rect 41713 195421 41883 195477
rect 41939 195421 41963 195477
rect 42019 195421 42043 195477
rect 42099 195421 42123 195477
rect 42179 195421 42193 195477
rect 41863 195414 42193 195421
rect 675407 194863 675737 194870
rect 41863 194833 42193 194840
rect 41713 194777 41883 194833
rect 41939 194777 41963 194833
rect 42019 194777 42043 194833
rect 42099 194777 42123 194833
rect 42179 194777 42193 194833
rect 675407 194807 675427 194863
rect 675483 194807 675507 194863
rect 675563 194807 675587 194863
rect 675643 194807 675667 194863
rect 675723 194807 675887 194863
rect 675407 194800 675737 194807
rect 41863 194770 42193 194777
rect 675407 193023 675737 193030
rect 41863 192993 42193 193000
rect 41713 192937 41883 192993
rect 41939 192937 41963 192993
rect 42019 192937 42043 192993
rect 42099 192937 42123 192993
rect 42179 192937 42193 192993
rect 675407 192967 675427 193023
rect 675483 192967 675507 193023
rect 675563 192967 675587 193023
rect 675643 192967 675667 193023
rect 675723 192967 675887 193023
rect 675407 192960 675737 192967
rect 41863 192930 42193 192937
rect 675407 192379 675737 192386
rect 675407 192323 675427 192379
rect 675483 192323 675507 192379
rect 675563 192323 675587 192379
rect 675643 192323 675667 192379
rect 675723 192323 675887 192379
rect 675407 192316 675737 192323
rect 41863 191797 42193 191804
rect 41713 191741 41883 191797
rect 41939 191741 41963 191797
rect 42019 191741 42043 191797
rect 42099 191741 42123 191797
rect 42179 191741 42193 191797
rect 41863 191734 42193 191741
rect 675407 191183 675737 191190
rect 41863 191153 42193 191160
rect 41713 191097 41883 191153
rect 41939 191097 41963 191153
rect 42019 191097 42043 191153
rect 42099 191097 42123 191153
rect 42179 191097 42193 191153
rect 675407 191127 675427 191183
rect 675483 191127 675507 191183
rect 675563 191127 675587 191183
rect 675643 191127 675667 191183
rect 675723 191127 675887 191183
rect 675407 191120 675737 191127
rect 41863 191090 42193 191097
rect 41863 190509 42193 190516
rect 41713 190453 41883 190509
rect 41939 190453 41963 190509
rect 42019 190453 42043 190509
rect 42099 190453 42123 190509
rect 42179 190453 42193 190509
rect 41863 190446 42193 190453
rect 41863 189957 42193 189964
rect 41713 189901 41883 189957
rect 41939 189901 41963 189957
rect 42019 189901 42043 189957
rect 42099 189901 42123 189957
rect 42179 189901 42193 189957
rect 41863 189894 42193 189901
rect 41863 187473 42193 187480
rect 41713 187417 41883 187473
rect 41939 187417 41963 187473
rect 42019 187417 42043 187473
rect 42099 187417 42123 187473
rect 42179 187417 42193 187473
rect 41863 187410 42193 187417
rect 41863 186829 42193 186836
rect 41713 186773 41883 186829
rect 41939 186773 41963 186829
rect 42019 186773 42043 186829
rect 42099 186773 42123 186829
rect 42179 186773 42193 186829
rect 41863 186766 42193 186773
rect 41863 186185 42193 186192
rect 41713 186129 41883 186185
rect 41939 186129 41963 186185
rect 42019 186129 42043 186185
rect 42099 186129 42123 186185
rect 42179 186129 42193 186185
rect 41863 186122 42193 186129
rect 41863 185633 42193 185640
rect 41713 185577 41883 185633
rect 41939 185577 41963 185633
rect 42019 185577 42043 185633
rect 42099 185577 42123 185633
rect 42179 185577 42193 185633
rect 41863 185570 42193 185577
rect 41863 183793 42193 183800
rect 41713 183737 41883 183793
rect 41939 183737 41963 183793
rect 42019 183737 42043 183793
rect 42099 183737 42123 183793
rect 42179 183737 42193 183793
rect 41863 183730 42193 183737
rect 41863 183149 42193 183156
rect 41713 183093 41883 183149
rect 41939 183093 41963 183149
rect 42019 183093 42043 183149
rect 42099 183093 42123 183149
rect 42179 183093 42193 183149
rect 41863 183086 42193 183093
rect 41863 182505 42193 182512
rect 41713 182449 41883 182505
rect 41939 182449 41963 182505
rect 42019 182449 42043 182505
rect 42099 182449 42123 182505
rect 42179 182449 42193 182505
rect 41863 182442 42193 182449
rect 675407 160351 675737 160358
rect 675407 160295 675427 160351
rect 675483 160295 675507 160351
rect 675563 160295 675587 160351
rect 675643 160295 675667 160351
rect 675723 160295 675887 160351
rect 675407 160288 675737 160295
rect 675407 159707 675737 159714
rect 675407 159651 675427 159707
rect 675483 159651 675507 159707
rect 675563 159651 675587 159707
rect 675643 159651 675667 159707
rect 675723 159651 675887 159707
rect 675407 159644 675737 159651
rect 675407 159063 675737 159070
rect 675407 159007 675427 159063
rect 675483 159007 675507 159063
rect 675563 159007 675587 159063
rect 675643 159007 675667 159063
rect 675723 159007 675887 159063
rect 675407 159000 675737 159007
rect 675407 157223 675737 157230
rect 675407 157167 675427 157223
rect 675483 157167 675507 157223
rect 675563 157167 675587 157223
rect 675643 157167 675667 157223
rect 675723 157167 675887 157223
rect 675407 157160 675737 157167
rect 675407 156671 675737 156678
rect 675407 156615 675427 156671
rect 675483 156615 675507 156671
rect 675563 156615 675587 156671
rect 675643 156615 675667 156671
rect 675723 156615 675887 156671
rect 675407 156608 675737 156615
rect 675407 156027 675737 156034
rect 675407 155971 675427 156027
rect 675483 155971 675507 156027
rect 675563 155971 675587 156027
rect 675643 155971 675667 156027
rect 675723 155971 675887 156027
rect 675407 155964 675737 155971
rect 675407 155383 675737 155390
rect 675407 155327 675427 155383
rect 675483 155327 675507 155383
rect 675563 155327 675587 155383
rect 675643 155327 675667 155383
rect 675723 155327 675887 155383
rect 675407 155320 675737 155327
rect 675407 152899 675737 152906
rect 675407 152843 675427 152899
rect 675483 152843 675507 152899
rect 675563 152843 675587 152899
rect 675643 152843 675667 152899
rect 675723 152843 675887 152899
rect 675407 152836 675737 152843
rect 675407 152347 675737 152354
rect 675407 152291 675427 152347
rect 675483 152291 675507 152347
rect 675563 152291 675587 152347
rect 675643 152291 675667 152347
rect 675723 152291 675887 152347
rect 675407 152284 675737 152291
rect 675407 151703 675737 151710
rect 675407 151647 675427 151703
rect 675483 151647 675507 151703
rect 675563 151647 675587 151703
rect 675643 151647 675667 151703
rect 675723 151647 675887 151703
rect 675407 151640 675737 151647
rect 675407 151059 675737 151066
rect 675407 151003 675427 151059
rect 675483 151003 675507 151059
rect 675563 151003 675587 151059
rect 675643 151003 675667 151059
rect 675723 151003 675887 151059
rect 675407 150996 675737 151003
rect 675407 149863 675737 149870
rect 675407 149807 675427 149863
rect 675483 149807 675507 149863
rect 675563 149807 675587 149863
rect 675643 149807 675667 149863
rect 675723 149807 675887 149863
rect 675407 149800 675737 149807
rect 675407 148023 675737 148030
rect 675407 147967 675427 148023
rect 675483 147967 675507 148023
rect 675563 147967 675587 148023
rect 675643 147967 675667 148023
rect 675723 147967 675887 148023
rect 675407 147960 675737 147967
rect 675407 147379 675737 147386
rect 675407 147323 675427 147379
rect 675483 147323 675507 147379
rect 675563 147323 675587 147379
rect 675643 147323 675667 147379
rect 675723 147323 675887 147379
rect 675407 147316 675737 147323
rect 675407 146183 675737 146190
rect 675407 146127 675427 146183
rect 675483 146127 675507 146183
rect 675563 146127 675587 146183
rect 675643 146127 675667 146183
rect 675723 146127 675887 146183
rect 675407 146120 675737 146127
rect 675407 115151 675737 115158
rect 675407 115095 675427 115151
rect 675483 115095 675507 115151
rect 675563 115095 675587 115151
rect 675643 115095 675667 115151
rect 675723 115095 675887 115151
rect 675407 115088 675737 115095
rect 675407 114507 675737 114514
rect 675407 114451 675427 114507
rect 675483 114451 675507 114507
rect 675563 114451 675587 114507
rect 675643 114451 675667 114507
rect 675723 114451 675887 114507
rect 675407 114444 675737 114451
rect 675407 113863 675737 113870
rect 675407 113807 675427 113863
rect 675483 113807 675507 113863
rect 675563 113807 675587 113863
rect 675643 113807 675667 113863
rect 675723 113807 675887 113863
rect 675407 113800 675737 113807
rect 675407 112023 675737 112030
rect 675407 111967 675427 112023
rect 675483 111967 675507 112023
rect 675563 111967 675587 112023
rect 675643 111967 675667 112023
rect 675723 111967 675887 112023
rect 675407 111960 675737 111967
rect 675407 111471 675737 111478
rect 675407 111415 675427 111471
rect 675483 111415 675507 111471
rect 675563 111415 675587 111471
rect 675643 111415 675667 111471
rect 675723 111415 675887 111471
rect 675407 111408 675737 111415
rect 675407 110827 675737 110834
rect 675407 110771 675427 110827
rect 675483 110771 675507 110827
rect 675563 110771 675587 110827
rect 675643 110771 675667 110827
rect 675723 110771 675887 110827
rect 675407 110764 675737 110771
rect 675407 110183 675737 110190
rect 675407 110127 675427 110183
rect 675483 110127 675507 110183
rect 675563 110127 675587 110183
rect 675643 110127 675667 110183
rect 675723 110127 675887 110183
rect 675407 110120 675737 110127
rect 675407 107699 675737 107706
rect 675407 107643 675427 107699
rect 675483 107643 675507 107699
rect 675563 107643 675587 107699
rect 675643 107643 675667 107699
rect 675723 107643 675887 107699
rect 675407 107636 675737 107643
rect 675407 107147 675737 107154
rect 675407 107091 675427 107147
rect 675483 107091 675507 107147
rect 675563 107091 675587 107147
rect 675643 107091 675667 107147
rect 675723 107091 675887 107147
rect 675407 107084 675737 107091
rect 675407 106503 675737 106510
rect 675407 106447 675427 106503
rect 675483 106447 675507 106503
rect 675563 106447 675587 106503
rect 675643 106447 675667 106503
rect 675723 106447 675887 106503
rect 675407 106440 675737 106447
rect 675407 105859 675737 105866
rect 675407 105803 675427 105859
rect 675483 105803 675507 105859
rect 675563 105803 675587 105859
rect 675643 105803 675667 105859
rect 675723 105803 675887 105859
rect 675407 105796 675737 105803
rect 675407 104663 675737 104670
rect 675407 104607 675427 104663
rect 675483 104607 675507 104663
rect 675563 104607 675587 104663
rect 675643 104607 675667 104663
rect 675723 104607 675887 104663
rect 675407 104600 675737 104607
rect 675407 102823 675737 102830
rect 675407 102767 675427 102823
rect 675483 102767 675507 102823
rect 675563 102767 675587 102823
rect 675643 102767 675667 102823
rect 675723 102767 675887 102823
rect 675407 102760 675737 102767
rect 675407 102179 675737 102186
rect 675407 102123 675427 102179
rect 675483 102123 675507 102179
rect 675563 102123 675587 102179
rect 675643 102123 675667 102179
rect 675723 102123 675887 102179
rect 675407 102116 675737 102123
rect 675407 100983 675737 100990
rect 675407 100927 675427 100983
rect 675483 100927 675507 100983
rect 675563 100927 675587 100983
rect 675643 100927 675667 100983
rect 675723 100927 675887 100983
rect 675407 100920 675737 100927
rect 465816 42528 465868 42534
rect 411076 42518 411128 42524
rect 411076 42460 411128 42466
rect 419724 42518 419776 42524
rect 465816 42470 465868 42476
rect 474464 42528 474516 42534
rect 474464 42470 474516 42476
rect 419724 42460 419776 42466
rect 409236 42392 409288 42398
rect 409236 42334 409288 42340
rect 195331 42231 195387 42242
rect 199655 42231 199711 42243
rect 303931 42231 303987 42240
rect 145035 42225 145207 42231
rect 145035 42173 145063 42225
rect 145115 42173 145127 42225
rect 145179 42173 145207 42225
rect 195328 42225 195387 42231
rect 145035 42167 145207 42173
rect 140996 40125 141048 40131
rect 141992 40125 142044 40131
rect 140996 40067 141048 40073
rect 141986 40073 141992 40120
rect 143068 40125 143120 40131
rect 142044 40073 142050 40120
rect 141004 39990 141042 40067
rect 141667 39934 141813 40000
rect 141986 39998 142050 40073
rect 143407 40125 143519 40131
rect 143407 40090 143437 40125
rect 143489 40090 143519 40125
rect 144603 40125 144655 40131
rect 143068 40067 143120 40073
rect 143078 39996 143110 40067
rect 143398 40034 143435 40090
rect 143491 40034 143528 40090
rect 144603 40067 144655 40073
rect 144610 39990 144652 40067
rect 145106 39990 145136 42167
rect 186683 41889 186735 41895
rect 186683 41831 186735 41837
rect 187327 41713 187383 42193
rect 188522 42141 188574 42147
rect 188522 42083 188574 42089
rect 192845 42141 192897 42147
rect 192845 42083 192897 42089
rect 189163 42057 189215 42063
rect 189163 41999 189215 42005
rect 191003 42057 191055 42063
rect 191003 41999 191055 42005
rect 192202 42057 192254 42063
rect 192202 41999 192254 42005
rect 193489 42057 193541 42063
rect 193489 41999 193541 42005
rect 187968 41973 188020 41979
rect 187968 41915 188020 41921
rect 194043 41713 194099 42193
rect 195380 42173 195387 42225
rect 195328 42167 195387 42173
rect 199653 42225 199711 42231
rect 199705 42173 199711 42225
rect 199653 42167 199711 42173
rect 303929 42225 303987 42231
rect 303981 42173 303987 42225
rect 308065 42225 308121 42248
rect 303929 42167 303987 42173
rect 195331 42137 195387 42167
rect 199655 42137 199711 42167
rect 201494 42141 201546 42147
rect 201494 42083 201546 42089
rect 202717 42141 202769 42147
rect 196528 42057 196580 42063
rect 196528 41999 196580 42005
rect 197170 42057 197222 42063
rect 197170 41999 197222 42005
rect 197813 42057 197865 42063
rect 197813 41999 197865 42005
rect 198368 42057 198420 42063
rect 198368 41999 198420 42005
rect 200206 42057 200258 42063
rect 200206 41999 200258 42005
rect 200857 42057 200909 42063
rect 200857 41999 200909 42005
rect 195973 41973 196025 41979
rect 195973 41915 196025 41921
rect 194688 41889 194740 41895
rect 194688 41831 194740 41837
rect 199012 41889 199064 41895
rect 199012 41831 199064 41837
rect 202717 40982 202769 42089
rect 297125 42141 297177 42147
rect 297125 42083 297177 42089
rect 299607 42141 299659 42147
rect 303931 42137 303987 42167
rect 305774 42141 305826 42147
rect 299607 42083 299659 42089
rect 305774 42083 305826 42089
rect 205928 42057 205980 42063
rect 145830 40974 145888 40981
rect 145828 40972 145888 40974
rect 145828 40916 145830 40972
rect 145886 40916 145888 40972
rect 145828 40903 145888 40916
rect 202713 40971 202773 40982
rect 205928 40981 205980 42005
rect 297768 42057 297820 42063
rect 297768 41999 297820 42005
rect 300804 42057 300856 42063
rect 300804 41999 300856 42005
rect 301451 42057 301503 42063
rect 301451 41999 301503 42005
rect 302094 42057 302146 42063
rect 302094 41999 302146 42005
rect 302643 42057 302695 42063
rect 302643 41999 302695 42005
rect 305133 42057 305185 42063
rect 305133 41999 305185 42005
rect 306418 42057 306470 42063
rect 306418 41999 306470 42005
rect 296576 41973 296628 41979
rect 296576 41915 296628 41921
rect 304577 41973 304629 41979
rect 304577 41915 304629 41921
rect 295283 41889 295335 41895
rect 295283 41831 295335 41837
rect 303290 41889 303342 41895
rect 303290 41831 303342 41837
rect 306967 41713 307023 42193
rect 308065 42173 308066 42225
rect 308118 42173 308121 42225
rect 358731 42225 358787 42240
rect 363055 42231 363111 42240
rect 308065 42129 308121 42173
rect 308255 42129 308311 42193
rect 308065 42073 308311 42129
rect 307616 41889 307668 41895
rect 307616 41831 307668 41837
rect 308255 41713 308311 42073
rect 308809 42057 308861 42063
rect 308809 41999 308861 42005
rect 309452 42057 309504 42063
rect 309452 41999 309504 42005
rect 310095 41713 310151 42193
rect 358731 42173 358732 42225
rect 358784 42173 358787 42225
rect 363053 42225 363111 42231
rect 311317 42141 311369 42147
rect 311317 40982 311369 42089
rect 351925 42141 351977 42147
rect 351925 42083 351977 42089
rect 354406 42141 354458 42147
rect 358731 42137 358787 42173
rect 360570 42141 360622 42147
rect 354406 42083 354458 42089
rect 360570 42083 360622 42089
rect 315497 42057 315549 42063
rect 202713 40915 202715 40971
rect 202771 40915 202773 40971
rect 202713 40904 202773 40915
rect 205924 40970 205984 40981
rect 205924 40914 205926 40970
rect 205982 40914 205984 40970
rect 205924 40903 205984 40914
rect 311313 40971 311373 40982
rect 315497 40976 315549 42005
rect 352568 42057 352620 42063
rect 352568 41999 352620 42005
rect 355600 42057 355652 42063
rect 355600 41999 355652 42005
rect 356246 42057 356298 42063
rect 356246 41999 356298 42005
rect 356889 42057 356941 42063
rect 356889 41999 356941 42005
rect 357444 42057 357496 42063
rect 357444 41999 357496 42005
rect 359928 42057 359980 42063
rect 359928 41999 359980 42005
rect 361217 42057 361269 42063
rect 361217 41999 361269 42005
rect 351375 41973 351427 41979
rect 351375 41915 351427 41921
rect 359374 41973 359426 41979
rect 359374 41915 359426 41921
rect 350086 41889 350138 41895
rect 350086 41831 350138 41837
rect 358090 41889 358142 41895
rect 358090 41831 358142 41837
rect 361767 41713 361823 42193
rect 363105 42173 363111 42225
rect 363053 42167 363111 42173
rect 363055 42137 363111 42167
rect 363607 42057 363659 42063
rect 363607 41999 363659 42005
rect 364252 42057 364304 42063
rect 364252 41999 364304 42005
rect 362412 41889 362464 41895
rect 362412 41831 362464 41837
rect 364895 41713 364951 42193
rect 366117 42141 366169 42147
rect 366117 40982 366169 42089
rect 370302 42057 370354 42063
rect 311313 40915 311315 40971
rect 311371 40915 311373 40971
rect 315484 40974 315562 40976
rect 315484 40918 315495 40974
rect 315551 40918 315562 40974
rect 315484 40916 315562 40918
rect 366113 40971 366173 40982
rect 370302 40981 370354 42005
rect 404877 41889 404929 41895
rect 404877 41831 404929 41837
rect 405527 41713 405583 42193
rect 406719 42141 406771 42147
rect 406719 42083 406771 42089
rect 407367 42057 407419 42063
rect 407367 41999 407419 42005
rect 406170 41973 406222 41979
rect 406170 41915 406222 41921
rect 409248 41820 409276 42334
rect 410398 42057 410450 42063
rect 410398 41999 410450 42005
rect 411088 41820 411116 42460
rect 412272 42392 412324 42398
rect 412272 42334 412324 42340
rect 415400 42392 415452 42398
rect 415400 42334 415452 42340
rect 412284 42193 412312 42334
rect 413531 42231 413587 42240
rect 411691 42057 411743 42063
rect 411691 41999 411743 42005
rect 412243 41820 412312 42193
rect 413524 42225 413587 42231
rect 413576 42173 413587 42225
rect 413524 42167 413587 42173
rect 413531 42135 413587 42167
rect 414725 42057 414777 42063
rect 414725 41999 414777 42005
rect 414174 41973 414226 41979
rect 414174 41915 414226 41921
rect 412888 41889 412940 41895
rect 412888 41831 412940 41837
rect 415412 41820 415440 42334
rect 417855 42225 417911 42236
rect 416013 42057 416065 42063
rect 416013 41999 416065 42005
rect 412243 41713 412299 41820
rect 416567 41713 416623 42193
rect 417855 42173 417858 42225
rect 417910 42173 417911 42225
rect 419736 42193 419764 42460
rect 464010 42380 464062 42386
rect 417855 42137 417911 42173
rect 418404 42057 418456 42063
rect 418404 41999 418456 42005
rect 419045 42057 419097 42063
rect 419045 41999 419097 42005
rect 417210 41889 417262 41895
rect 417210 41831 417262 41837
rect 419695 41820 419764 42193
rect 420917 42141 420969 42147
rect 419695 41713 419751 41820
rect 420917 40982 420969 42089
rect 425115 42057 425167 42063
rect 311313 40904 311373 40915
rect 366113 40915 366115 40971
rect 366171 40915 366173 40971
rect 366113 40904 366173 40915
rect 370298 40970 370358 40981
rect 370298 40914 370300 40970
rect 370356 40914 370358 40970
rect 370298 40903 370358 40914
rect 420913 40971 420973 40982
rect 420913 40915 420915 40971
rect 420971 40915 420973 40971
rect 425115 40969 425167 42005
rect 459678 41889 459730 41895
rect 459678 41831 459730 41837
rect 460327 41713 460383 42193
rect 464010 42180 464062 42328
rect 461524 42141 461576 42147
rect 461524 42083 461576 42089
rect 462162 42057 462214 42063
rect 462162 41999 462214 42005
rect 465201 42057 465253 42063
rect 465201 41999 465253 42005
rect 460971 41973 461023 41979
rect 460971 41915 461023 41921
rect 465828 41834 465856 42470
rect 467046 42380 467098 42386
rect 467046 42193 467098 42328
rect 470173 42380 470225 42386
rect 468331 42231 468387 42245
rect 468330 42225 468387 42231
rect 466488 42057 466540 42063
rect 466488 41999 466540 42005
rect 465828 41806 465875 41834
rect 467043 41713 467099 42193
rect 468382 42173 468387 42225
rect 470173 42181 470225 42328
rect 472655 42225 472711 42235
rect 468330 42167 468387 42173
rect 468331 42135 468387 42167
rect 469522 42057 469574 42063
rect 469522 41999 469574 42005
rect 470810 42057 470862 42063
rect 470810 41999 470862 42005
rect 468967 41973 469019 41979
rect 468967 41915 469019 41921
rect 467684 41889 467736 41895
rect 467684 41831 467736 41837
rect 471367 41713 471423 42193
rect 472655 42173 472656 42225
rect 472708 42173 472711 42225
rect 472655 42132 472711 42173
rect 474476 42193 474504 42470
rect 518808 42392 518860 42398
rect 518808 42334 518860 42340
rect 524972 42392 525024 42398
rect 524972 42334 525024 42340
rect 473201 42057 473253 42063
rect 473201 41999 473253 42005
rect 473849 42057 473901 42063
rect 473849 41999 473901 42005
rect 472010 41889 472062 41895
rect 472010 41831 472062 41837
rect 474476 41806 474551 42193
rect 474495 41713 474551 41806
rect 475717 42141 475769 42147
rect 475717 40982 475769 42089
rect 479915 42057 479967 42063
rect 479915 40983 479967 42005
rect 514487 41889 514539 41895
rect 514487 41831 514539 41837
rect 515127 41713 515183 42193
rect 516320 42141 516372 42147
rect 516320 42083 516372 42089
rect 516969 42057 517021 42063
rect 516969 41999 517021 42005
rect 515772 41973 515824 41979
rect 515772 41915 515824 41921
rect 518820 41820 518848 42334
rect 523131 42231 523187 42251
rect 523126 42225 523187 42231
rect 520004 42057 520056 42063
rect 520004 41999 520056 42005
rect 520647 41713 520703 42193
rect 521293 42057 521345 42063
rect 521293 41999 521345 42005
rect 521843 41713 521899 42193
rect 523178 42173 523187 42225
rect 524984 42193 525012 42334
rect 527455 42225 527511 42249
rect 523126 42167 523187 42173
rect 523131 42128 523187 42167
rect 524328 42057 524380 42063
rect 524328 41999 524380 42005
rect 523773 41973 523825 41979
rect 523773 41915 523825 41921
rect 522486 41889 522538 41895
rect 522486 41831 522538 41837
rect 524971 41713 525027 42193
rect 525615 42057 525667 42063
rect 525615 41999 525667 42005
rect 526167 41713 526223 42193
rect 527455 42173 527457 42225
rect 527509 42173 527511 42225
rect 527455 42120 527511 42173
rect 528009 42057 528061 42063
rect 528009 41999 528061 42005
rect 528652 42057 528704 42063
rect 528652 41999 528704 42005
rect 526810 41889 526862 41895
rect 526810 41831 526862 41837
rect 529295 41713 529351 42193
rect 530517 42141 530569 42147
rect 475713 40971 475773 40982
rect 420913 40904 420973 40915
rect 425111 40958 425171 40969
rect 145852 40134 145888 40903
rect 425111 40902 425113 40958
rect 425169 40902 425171 40958
rect 475713 40915 475715 40971
rect 475771 40915 475773 40971
rect 475713 40904 475773 40915
rect 479911 40972 479971 40983
rect 530517 40982 530569 42089
rect 534772 42057 534824 42063
rect 479911 40916 479913 40972
rect 479969 40916 479971 40972
rect 479911 40905 479971 40916
rect 530513 40971 530573 40982
rect 534772 40971 534824 42005
rect 530513 40915 530515 40971
rect 530571 40915 530573 40971
rect 530513 40904 530573 40915
rect 534768 40960 534828 40971
rect 534768 40904 534770 40960
rect 534826 40904 534828 40960
rect 425111 40891 425171 40902
rect 534768 40893 534828 40904
rect 145828 40132 145906 40134
rect 145828 40076 145839 40132
rect 145895 40076 145906 40132
rect 145828 40074 145906 40076
<< via2 >>
rect 41883 969217 41939 969273
rect 41963 969217 42019 969273
rect 42043 969217 42099 969273
rect 42123 969217 42179 969273
rect 41883 968021 41939 968077
rect 41963 968021 42019 968077
rect 42043 968021 42099 968077
rect 42123 968021 42179 968077
rect 41883 967377 41939 967433
rect 41963 967377 42019 967433
rect 42043 967377 42099 967433
rect 42123 967377 42179 967433
rect 41883 966733 41939 966789
rect 41963 966733 42019 966789
rect 42043 966733 42099 966789
rect 42123 966733 42179 966789
rect 675427 966695 675483 966751
rect 675507 966695 675563 966751
rect 675587 966695 675643 966751
rect 675667 966695 675723 966751
rect 675427 966051 675483 966107
rect 675507 966051 675563 966107
rect 675587 966051 675643 966107
rect 675667 966051 675723 966107
rect 41883 965537 41939 965593
rect 41963 965537 42019 965593
rect 42043 965537 42099 965593
rect 42123 965537 42179 965593
rect 675427 965407 675483 965463
rect 675507 965407 675563 965463
rect 675587 965407 675643 965463
rect 675667 965407 675723 965463
rect 41883 964341 41939 964397
rect 41963 964341 42019 964397
rect 42043 964341 42099 964397
rect 42123 964341 42179 964397
rect 41883 963697 41939 963753
rect 41963 963697 42019 963753
rect 42043 963697 42099 963753
rect 42123 963697 42179 963753
rect 675427 963567 675483 963623
rect 675507 963567 675563 963623
rect 675587 963567 675643 963623
rect 675667 963567 675723 963623
rect 41883 963053 41939 963109
rect 41963 963053 42019 963109
rect 42043 963053 42099 963109
rect 42123 963053 42179 963109
rect 675427 963015 675483 963071
rect 675507 963015 675563 963071
rect 675587 963015 675643 963071
rect 675667 963015 675723 963071
rect 41883 962501 41939 962557
rect 41963 962501 42019 962557
rect 42043 962501 42099 962557
rect 42123 962501 42179 962557
rect 675427 962371 675483 962427
rect 675507 962371 675563 962427
rect 675587 962371 675643 962427
rect 675667 962371 675723 962427
rect 675427 961727 675483 961783
rect 675507 961727 675563 961783
rect 675587 961727 675643 961783
rect 675667 961727 675723 961783
rect 41883 960017 41939 960073
rect 41963 960017 42019 960073
rect 42043 960017 42099 960073
rect 42123 960017 42179 960073
rect 41883 959373 41939 959429
rect 41963 959373 42019 959429
rect 42043 959373 42099 959429
rect 42123 959373 42179 959429
rect 675427 959243 675483 959299
rect 675507 959243 675563 959299
rect 675587 959243 675643 959299
rect 675667 959243 675723 959299
rect 41883 958729 41939 958785
rect 41963 958729 42019 958785
rect 42043 958729 42099 958785
rect 42123 958729 42179 958785
rect 675427 958691 675483 958747
rect 675507 958691 675563 958747
rect 675587 958691 675643 958747
rect 675667 958691 675723 958747
rect 41883 958177 41939 958233
rect 41963 958177 42019 958233
rect 42043 958177 42099 958233
rect 42123 958177 42179 958233
rect 675427 958047 675483 958103
rect 675507 958047 675563 958103
rect 675587 958047 675643 958103
rect 675667 958047 675723 958103
rect 675427 957403 675483 957459
rect 675507 957403 675563 957459
rect 675587 957403 675643 957459
rect 675667 957403 675723 957459
rect 41883 956337 41939 956393
rect 41963 956337 42019 956393
rect 42043 956337 42099 956393
rect 42123 956337 42179 956393
rect 675427 956207 675483 956263
rect 675507 956207 675563 956263
rect 675587 956207 675643 956263
rect 675667 956207 675723 956263
rect 41883 955693 41939 955749
rect 41963 955693 42019 955749
rect 42043 955693 42099 955749
rect 42123 955693 42179 955749
rect 41883 955049 41939 955105
rect 41963 955049 42019 955105
rect 42043 955049 42099 955105
rect 42123 955049 42179 955105
rect 675427 955011 675483 955067
rect 675507 955011 675563 955067
rect 675587 955011 675643 955067
rect 675667 955011 675723 955067
rect 675427 954367 675483 954423
rect 675507 954367 675563 954423
rect 675587 954367 675643 954423
rect 675667 954367 675723 954423
rect 675427 953723 675483 953779
rect 675507 953723 675563 953779
rect 675587 953723 675643 953779
rect 675667 953723 675723 953779
rect 675427 952527 675483 952583
rect 675507 952527 675563 952583
rect 675587 952527 675643 952583
rect 675667 952527 675723 952583
rect 675427 877495 675483 877551
rect 675507 877495 675563 877551
rect 675587 877495 675643 877551
rect 675667 877495 675723 877551
rect 675427 876851 675483 876907
rect 675507 876851 675563 876907
rect 675587 876851 675643 876907
rect 675667 876851 675723 876907
rect 675427 876207 675483 876263
rect 675507 876207 675563 876263
rect 675587 876207 675643 876263
rect 675667 876207 675723 876263
rect 675427 874367 675483 874423
rect 675507 874367 675563 874423
rect 675587 874367 675643 874423
rect 675667 874367 675723 874423
rect 675427 873815 675483 873871
rect 675507 873815 675563 873871
rect 675587 873815 675643 873871
rect 675667 873815 675723 873871
rect 675427 873171 675483 873227
rect 675507 873171 675563 873227
rect 675587 873171 675643 873227
rect 675667 873171 675723 873227
rect 675427 872527 675483 872583
rect 675507 872527 675563 872583
rect 675587 872527 675643 872583
rect 675667 872527 675723 872583
rect 675427 870043 675483 870099
rect 675507 870043 675563 870099
rect 675587 870043 675643 870099
rect 675667 870043 675723 870099
rect 675427 869491 675483 869547
rect 675507 869491 675563 869547
rect 675587 869491 675643 869547
rect 675667 869491 675723 869547
rect 675427 868847 675483 868903
rect 675507 868847 675563 868903
rect 675587 868847 675643 868903
rect 675667 868847 675723 868903
rect 675427 868203 675483 868259
rect 675507 868203 675563 868259
rect 675587 868203 675643 868259
rect 675667 868203 675723 868259
rect 675427 867007 675483 867063
rect 675507 867007 675563 867063
rect 675587 867007 675643 867063
rect 675667 867007 675723 867063
rect 675427 865811 675483 865867
rect 675507 865811 675563 865867
rect 675587 865811 675643 865867
rect 675667 865811 675723 865867
rect 675427 865167 675483 865223
rect 675507 865167 675563 865223
rect 675587 865167 675643 865223
rect 675667 865167 675723 865223
rect 675427 864523 675483 864579
rect 675507 864523 675563 864579
rect 675587 864523 675643 864579
rect 675667 864523 675723 864579
rect 675427 863327 675483 863383
rect 675507 863327 675563 863383
rect 675587 863327 675643 863383
rect 675667 863327 675723 863383
rect 41883 799417 41939 799473
rect 41963 799417 42019 799473
rect 42043 799417 42099 799473
rect 42123 799417 42179 799473
rect 41883 798221 41939 798277
rect 41963 798221 42019 798277
rect 42043 798221 42099 798277
rect 42123 798221 42179 798277
rect 41883 797577 41939 797633
rect 41963 797577 42019 797633
rect 42043 797577 42099 797633
rect 42123 797577 42179 797633
rect 41883 796933 41939 796989
rect 41963 796933 42019 796989
rect 42043 796933 42099 796989
rect 42123 796933 42179 796989
rect 41883 795737 41939 795793
rect 41963 795737 42019 795793
rect 42043 795737 42099 795793
rect 42123 795737 42179 795793
rect 41883 794541 41939 794597
rect 41963 794541 42019 794597
rect 42043 794541 42099 794597
rect 42123 794541 42179 794597
rect 41883 793897 41939 793953
rect 41963 793897 42019 793953
rect 42043 793897 42099 793953
rect 42123 793897 42179 793953
rect 41883 793253 41939 793309
rect 41963 793253 42019 793309
rect 42043 793253 42099 793309
rect 42123 793253 42179 793309
rect 41883 792701 41939 792757
rect 41963 792701 42019 792757
rect 42043 792701 42099 792757
rect 42123 792701 42179 792757
rect 41883 790217 41939 790273
rect 41963 790217 42019 790273
rect 42043 790217 42099 790273
rect 42123 790217 42179 790273
rect 41883 789573 41939 789629
rect 41963 789573 42019 789629
rect 42043 789573 42099 789629
rect 42123 789573 42179 789629
rect 41883 788929 41939 788985
rect 41963 788929 42019 788985
rect 42043 788929 42099 788985
rect 42123 788929 42179 788985
rect 41883 788377 41939 788433
rect 41963 788377 42019 788433
rect 42043 788377 42099 788433
rect 42123 788377 42179 788433
rect 675427 788295 675483 788351
rect 675507 788295 675563 788351
rect 675587 788295 675643 788351
rect 675667 788295 675723 788351
rect 675427 787651 675483 787707
rect 675507 787651 675563 787707
rect 675587 787651 675643 787707
rect 675667 787651 675723 787707
rect 675427 787007 675483 787063
rect 675507 787007 675563 787063
rect 675587 787007 675643 787063
rect 675667 787007 675723 787063
rect 41883 786537 41939 786593
rect 41963 786537 42019 786593
rect 42043 786537 42099 786593
rect 42123 786537 42179 786593
rect 41883 785893 41939 785949
rect 41963 785893 42019 785949
rect 42043 785893 42099 785949
rect 42123 785893 42179 785949
rect 41883 785249 41939 785305
rect 41963 785249 42019 785305
rect 42043 785249 42099 785305
rect 42123 785249 42179 785305
rect 675427 785167 675483 785223
rect 675507 785167 675563 785223
rect 675587 785167 675643 785223
rect 675667 785167 675723 785223
rect 675427 784615 675483 784671
rect 675507 784615 675563 784671
rect 675587 784615 675643 784671
rect 675667 784615 675723 784671
rect 675427 783971 675483 784027
rect 675507 783971 675563 784027
rect 675587 783971 675643 784027
rect 675667 783971 675723 784027
rect 675427 783327 675483 783383
rect 675507 783327 675563 783383
rect 675587 783327 675643 783383
rect 675667 783327 675723 783383
rect 675427 780843 675483 780899
rect 675507 780843 675563 780899
rect 675587 780843 675643 780899
rect 675667 780843 675723 780899
rect 675427 780291 675483 780347
rect 675507 780291 675563 780347
rect 675587 780291 675643 780347
rect 675667 780291 675723 780347
rect 675427 779647 675483 779703
rect 675507 779647 675563 779703
rect 675587 779647 675643 779703
rect 675667 779647 675723 779703
rect 675427 779003 675483 779059
rect 675507 779003 675563 779059
rect 675587 779003 675643 779059
rect 675667 779003 675723 779059
rect 675427 777807 675483 777863
rect 675507 777807 675563 777863
rect 675587 777807 675643 777863
rect 675667 777807 675723 777863
rect 675427 776611 675483 776667
rect 675507 776611 675563 776667
rect 675587 776611 675643 776667
rect 675667 776611 675723 776667
rect 675427 775967 675483 776023
rect 675507 775967 675563 776023
rect 675587 775967 675643 776023
rect 675667 775967 675723 776023
rect 675427 775323 675483 775379
rect 675507 775323 675563 775379
rect 675587 775323 675643 775379
rect 675667 775323 675723 775379
rect 675427 774127 675483 774183
rect 675507 774127 675563 774183
rect 675587 774127 675643 774183
rect 675667 774127 675723 774183
rect 41883 756217 41939 756273
rect 41963 756217 42019 756273
rect 42043 756217 42099 756273
rect 42123 756217 42179 756273
rect 41883 755021 41939 755077
rect 41963 755021 42019 755077
rect 42043 755021 42099 755077
rect 42123 755021 42179 755077
rect 41883 754377 41939 754433
rect 41963 754377 42019 754433
rect 42043 754377 42099 754433
rect 42123 754377 42179 754433
rect 41883 753733 41939 753789
rect 41963 753733 42019 753789
rect 42043 753733 42099 753789
rect 42123 753733 42179 753789
rect 41883 752537 41939 752593
rect 41963 752537 42019 752593
rect 42043 752537 42099 752593
rect 42123 752537 42179 752593
rect 41883 751341 41939 751397
rect 41963 751341 42019 751397
rect 42043 751341 42099 751397
rect 42123 751341 42179 751397
rect 41883 750697 41939 750753
rect 41963 750697 42019 750753
rect 42043 750697 42099 750753
rect 42123 750697 42179 750753
rect 41883 750053 41939 750109
rect 41963 750053 42019 750109
rect 42043 750053 42099 750109
rect 42123 750053 42179 750109
rect 41883 749501 41939 749557
rect 41963 749501 42019 749557
rect 42043 749501 42099 749557
rect 42123 749501 42179 749557
rect 41883 747017 41939 747073
rect 41963 747017 42019 747073
rect 42043 747017 42099 747073
rect 42123 747017 42179 747073
rect 41883 746373 41939 746429
rect 41963 746373 42019 746429
rect 42043 746373 42099 746429
rect 42123 746373 42179 746429
rect 41883 745729 41939 745785
rect 41963 745729 42019 745785
rect 42043 745729 42099 745785
rect 42123 745729 42179 745785
rect 41883 745177 41939 745233
rect 41963 745177 42019 745233
rect 42043 745177 42099 745233
rect 42123 745177 42179 745233
rect 41883 743337 41939 743393
rect 41963 743337 42019 743393
rect 42043 743337 42099 743393
rect 42123 743337 42179 743393
rect 675427 743295 675483 743351
rect 675507 743295 675563 743351
rect 675587 743295 675643 743351
rect 675667 743295 675723 743351
rect 41883 742693 41939 742749
rect 41963 742693 42019 742749
rect 42043 742693 42099 742749
rect 42123 742693 42179 742749
rect 675427 742651 675483 742707
rect 675507 742651 675563 742707
rect 675587 742651 675643 742707
rect 675667 742651 675723 742707
rect 41883 742049 41939 742105
rect 41963 742049 42019 742105
rect 42043 742049 42099 742105
rect 42123 742049 42179 742105
rect 675427 742007 675483 742063
rect 675507 742007 675563 742063
rect 675587 742007 675643 742063
rect 675667 742007 675723 742063
rect 675427 740167 675483 740223
rect 675507 740167 675563 740223
rect 675587 740167 675643 740223
rect 675667 740167 675723 740223
rect 675427 739615 675483 739671
rect 675507 739615 675563 739671
rect 675587 739615 675643 739671
rect 675667 739615 675723 739671
rect 675427 738971 675483 739027
rect 675507 738971 675563 739027
rect 675587 738971 675643 739027
rect 675667 738971 675723 739027
rect 675427 738327 675483 738383
rect 675507 738327 675563 738383
rect 675587 738327 675643 738383
rect 675667 738327 675723 738383
rect 675427 735843 675483 735899
rect 675507 735843 675563 735899
rect 675587 735843 675643 735899
rect 675667 735843 675723 735899
rect 675427 735291 675483 735347
rect 675507 735291 675563 735347
rect 675587 735291 675643 735347
rect 675667 735291 675723 735347
rect 675427 734647 675483 734703
rect 675507 734647 675563 734703
rect 675587 734647 675643 734703
rect 675667 734647 675723 734703
rect 675427 734003 675483 734059
rect 675507 734003 675563 734059
rect 675587 734003 675643 734059
rect 675667 734003 675723 734059
rect 675427 732807 675483 732863
rect 675507 732807 675563 732863
rect 675587 732807 675643 732863
rect 675667 732807 675723 732863
rect 675427 731611 675483 731667
rect 675507 731611 675563 731667
rect 675587 731611 675643 731667
rect 675667 731611 675723 731667
rect 675427 730967 675483 731023
rect 675507 730967 675563 731023
rect 675587 730967 675643 731023
rect 675667 730967 675723 731023
rect 675427 730323 675483 730379
rect 675507 730323 675563 730379
rect 675587 730323 675643 730379
rect 675667 730323 675723 730379
rect 675427 729127 675483 729183
rect 675507 729127 675563 729183
rect 675587 729127 675643 729183
rect 675667 729127 675723 729183
rect 41883 713017 41939 713073
rect 41963 713017 42019 713073
rect 42043 713017 42099 713073
rect 42123 713017 42179 713073
rect 41883 711821 41939 711877
rect 41963 711821 42019 711877
rect 42043 711821 42099 711877
rect 42123 711821 42179 711877
rect 41883 711177 41939 711233
rect 41963 711177 42019 711233
rect 42043 711177 42099 711233
rect 42123 711177 42179 711233
rect 41883 710533 41939 710589
rect 41963 710533 42019 710589
rect 42043 710533 42099 710589
rect 42123 710533 42179 710589
rect 41883 709337 41939 709393
rect 41963 709337 42019 709393
rect 42043 709337 42099 709393
rect 42123 709337 42179 709393
rect 41883 708141 41939 708197
rect 41963 708141 42019 708197
rect 42043 708141 42099 708197
rect 42123 708141 42179 708197
rect 41883 707497 41939 707553
rect 41963 707497 42019 707553
rect 42043 707497 42099 707553
rect 42123 707497 42179 707553
rect 41883 706853 41939 706909
rect 41963 706853 42019 706909
rect 42043 706853 42099 706909
rect 42123 706853 42179 706909
rect 41883 706301 41939 706357
rect 41963 706301 42019 706357
rect 42043 706301 42099 706357
rect 42123 706301 42179 706357
rect 41883 703817 41939 703873
rect 41963 703817 42019 703873
rect 42043 703817 42099 703873
rect 42123 703817 42179 703873
rect 41883 703173 41939 703229
rect 41963 703173 42019 703229
rect 42043 703173 42099 703229
rect 42123 703173 42179 703229
rect 41883 702529 41939 702585
rect 41963 702529 42019 702585
rect 42043 702529 42099 702585
rect 42123 702529 42179 702585
rect 41883 701977 41939 702033
rect 41963 701977 42019 702033
rect 42043 701977 42099 702033
rect 42123 701977 42179 702033
rect 41883 700137 41939 700193
rect 41963 700137 42019 700193
rect 42043 700137 42099 700193
rect 42123 700137 42179 700193
rect 41883 699493 41939 699549
rect 41963 699493 42019 699549
rect 42043 699493 42099 699549
rect 42123 699493 42179 699549
rect 41883 698849 41939 698905
rect 41963 698849 42019 698905
rect 42043 698849 42099 698905
rect 42123 698849 42179 698905
rect 675427 698295 675483 698351
rect 675507 698295 675563 698351
rect 675587 698295 675643 698351
rect 675667 698295 675723 698351
rect 675427 697651 675483 697707
rect 675507 697651 675563 697707
rect 675587 697651 675643 697707
rect 675667 697651 675723 697707
rect 675427 697007 675483 697063
rect 675507 697007 675563 697063
rect 675587 697007 675643 697063
rect 675667 697007 675723 697063
rect 675427 695167 675483 695223
rect 675507 695167 675563 695223
rect 675587 695167 675643 695223
rect 675667 695167 675723 695223
rect 675427 694615 675483 694671
rect 675507 694615 675563 694671
rect 675587 694615 675643 694671
rect 675667 694615 675723 694671
rect 675427 693971 675483 694027
rect 675507 693971 675563 694027
rect 675587 693971 675643 694027
rect 675667 693971 675723 694027
rect 675427 693327 675483 693383
rect 675507 693327 675563 693383
rect 675587 693327 675643 693383
rect 675667 693327 675723 693383
rect 675427 690843 675483 690899
rect 675507 690843 675563 690899
rect 675587 690843 675643 690899
rect 675667 690843 675723 690899
rect 675427 690291 675483 690347
rect 675507 690291 675563 690347
rect 675587 690291 675643 690347
rect 675667 690291 675723 690347
rect 675427 689647 675483 689703
rect 675507 689647 675563 689703
rect 675587 689647 675643 689703
rect 675667 689647 675723 689703
rect 675427 689003 675483 689059
rect 675507 689003 675563 689059
rect 675587 689003 675643 689059
rect 675667 689003 675723 689059
rect 675427 687807 675483 687863
rect 675507 687807 675563 687863
rect 675587 687807 675643 687863
rect 675667 687807 675723 687863
rect 675427 686611 675483 686667
rect 675507 686611 675563 686667
rect 675587 686611 675643 686667
rect 675667 686611 675723 686667
rect 675427 685967 675483 686023
rect 675507 685967 675563 686023
rect 675587 685967 675643 686023
rect 675667 685967 675723 686023
rect 675427 685323 675483 685379
rect 675507 685323 675563 685379
rect 675587 685323 675643 685379
rect 675667 685323 675723 685379
rect 675427 684127 675483 684183
rect 675507 684127 675563 684183
rect 675587 684127 675643 684183
rect 675667 684127 675723 684183
rect 41883 669817 41939 669873
rect 41963 669817 42019 669873
rect 42043 669817 42099 669873
rect 42123 669817 42179 669873
rect 41883 668621 41939 668677
rect 41963 668621 42019 668677
rect 42043 668621 42099 668677
rect 42123 668621 42179 668677
rect 41883 667977 41939 668033
rect 41963 667977 42019 668033
rect 42043 667977 42099 668033
rect 42123 667977 42179 668033
rect 41883 667333 41939 667389
rect 41963 667333 42019 667389
rect 42043 667333 42099 667389
rect 42123 667333 42179 667389
rect 41883 666137 41939 666193
rect 41963 666137 42019 666193
rect 42043 666137 42099 666193
rect 42123 666137 42179 666193
rect 41883 664941 41939 664997
rect 41963 664941 42019 664997
rect 42043 664941 42099 664997
rect 42123 664941 42179 664997
rect 41883 664297 41939 664353
rect 41963 664297 42019 664353
rect 42043 664297 42099 664353
rect 42123 664297 42179 664353
rect 41883 663653 41939 663709
rect 41963 663653 42019 663709
rect 42043 663653 42099 663709
rect 42123 663653 42179 663709
rect 41883 663101 41939 663157
rect 41963 663101 42019 663157
rect 42043 663101 42099 663157
rect 42123 663101 42179 663157
rect 41883 660617 41939 660673
rect 41963 660617 42019 660673
rect 42043 660617 42099 660673
rect 42123 660617 42179 660673
rect 41883 659973 41939 660029
rect 41963 659973 42019 660029
rect 42043 659973 42099 660029
rect 42123 659973 42179 660029
rect 41883 659329 41939 659385
rect 41963 659329 42019 659385
rect 42043 659329 42099 659385
rect 42123 659329 42179 659385
rect 41883 658777 41939 658833
rect 41963 658777 42019 658833
rect 42043 658777 42099 658833
rect 42123 658777 42179 658833
rect 41883 656937 41939 656993
rect 41963 656937 42019 656993
rect 42043 656937 42099 656993
rect 42123 656937 42179 656993
rect 41883 656293 41939 656349
rect 41963 656293 42019 656349
rect 42043 656293 42099 656349
rect 42123 656293 42179 656349
rect 41883 655649 41939 655705
rect 41963 655649 42019 655705
rect 42043 655649 42099 655705
rect 42123 655649 42179 655705
rect 675427 653095 675483 653151
rect 675507 653095 675563 653151
rect 675587 653095 675643 653151
rect 675667 653095 675723 653151
rect 675427 652451 675483 652507
rect 675507 652451 675563 652507
rect 675587 652451 675643 652507
rect 675667 652451 675723 652507
rect 675427 651807 675483 651863
rect 675507 651807 675563 651863
rect 675587 651807 675643 651863
rect 675667 651807 675723 651863
rect 675427 649967 675483 650023
rect 675507 649967 675563 650023
rect 675587 649967 675643 650023
rect 675667 649967 675723 650023
rect 675427 649415 675483 649471
rect 675507 649415 675563 649471
rect 675587 649415 675643 649471
rect 675667 649415 675723 649471
rect 675427 648771 675483 648827
rect 675507 648771 675563 648827
rect 675587 648771 675643 648827
rect 675667 648771 675723 648827
rect 675427 648127 675483 648183
rect 675507 648127 675563 648183
rect 675587 648127 675643 648183
rect 675667 648127 675723 648183
rect 675427 645643 675483 645699
rect 675507 645643 675563 645699
rect 675587 645643 675643 645699
rect 675667 645643 675723 645699
rect 675427 645091 675483 645147
rect 675507 645091 675563 645147
rect 675587 645091 675643 645147
rect 675667 645091 675723 645147
rect 675427 644447 675483 644503
rect 675507 644447 675563 644503
rect 675587 644447 675643 644503
rect 675667 644447 675723 644503
rect 675427 643803 675483 643859
rect 675507 643803 675563 643859
rect 675587 643803 675643 643859
rect 675667 643803 675723 643859
rect 675427 642607 675483 642663
rect 675507 642607 675563 642663
rect 675587 642607 675643 642663
rect 675667 642607 675723 642663
rect 675427 641411 675483 641467
rect 675507 641411 675563 641467
rect 675587 641411 675643 641467
rect 675667 641411 675723 641467
rect 675427 640767 675483 640823
rect 675507 640767 675563 640823
rect 675587 640767 675643 640823
rect 675667 640767 675723 640823
rect 675427 640123 675483 640179
rect 675507 640123 675563 640179
rect 675587 640123 675643 640179
rect 675667 640123 675723 640179
rect 675427 638927 675483 638983
rect 675507 638927 675563 638983
rect 675587 638927 675643 638983
rect 675667 638927 675723 638983
rect 41883 626617 41939 626673
rect 41963 626617 42019 626673
rect 42043 626617 42099 626673
rect 42123 626617 42179 626673
rect 41883 625421 41939 625477
rect 41963 625421 42019 625477
rect 42043 625421 42099 625477
rect 42123 625421 42179 625477
rect 41883 624777 41939 624833
rect 41963 624777 42019 624833
rect 42043 624777 42099 624833
rect 42123 624777 42179 624833
rect 41883 624133 41939 624189
rect 41963 624133 42019 624189
rect 42043 624133 42099 624189
rect 42123 624133 42179 624189
rect 41883 622937 41939 622993
rect 41963 622937 42019 622993
rect 42043 622937 42099 622993
rect 42123 622937 42179 622993
rect 41883 621741 41939 621797
rect 41963 621741 42019 621797
rect 42043 621741 42099 621797
rect 42123 621741 42179 621797
rect 41883 621097 41939 621153
rect 41963 621097 42019 621153
rect 42043 621097 42099 621153
rect 42123 621097 42179 621153
rect 41883 620453 41939 620509
rect 41963 620453 42019 620509
rect 42043 620453 42099 620509
rect 42123 620453 42179 620509
rect 41883 619901 41939 619957
rect 41963 619901 42019 619957
rect 42043 619901 42099 619957
rect 42123 619901 42179 619957
rect 41883 617417 41939 617473
rect 41963 617417 42019 617473
rect 42043 617417 42099 617473
rect 42123 617417 42179 617473
rect 41883 616773 41939 616829
rect 41963 616773 42019 616829
rect 42043 616773 42099 616829
rect 42123 616773 42179 616829
rect 41883 616129 41939 616185
rect 41963 616129 42019 616185
rect 42043 616129 42099 616185
rect 42123 616129 42179 616185
rect 41883 615577 41939 615633
rect 41963 615577 42019 615633
rect 42043 615577 42099 615633
rect 42123 615577 42179 615633
rect 41883 613737 41939 613793
rect 41963 613737 42019 613793
rect 42043 613737 42099 613793
rect 42123 613737 42179 613793
rect 41883 613093 41939 613149
rect 41963 613093 42019 613149
rect 42043 613093 42099 613149
rect 42123 613093 42179 613149
rect 41883 612449 41939 612505
rect 41963 612449 42019 612505
rect 42043 612449 42099 612505
rect 42123 612449 42179 612505
rect 675427 608095 675483 608151
rect 675507 608095 675563 608151
rect 675587 608095 675643 608151
rect 675667 608095 675723 608151
rect 675427 607451 675483 607507
rect 675507 607451 675563 607507
rect 675587 607451 675643 607507
rect 675667 607451 675723 607507
rect 675427 606807 675483 606863
rect 675507 606807 675563 606863
rect 675587 606807 675643 606863
rect 675667 606807 675723 606863
rect 675427 604967 675483 605023
rect 675507 604967 675563 605023
rect 675587 604967 675643 605023
rect 675667 604967 675723 605023
rect 675427 604415 675483 604471
rect 675507 604415 675563 604471
rect 675587 604415 675643 604471
rect 675667 604415 675723 604471
rect 675427 603771 675483 603827
rect 675507 603771 675563 603827
rect 675587 603771 675643 603827
rect 675667 603771 675723 603827
rect 675427 603127 675483 603183
rect 675507 603127 675563 603183
rect 675587 603127 675643 603183
rect 675667 603127 675723 603183
rect 675427 600643 675483 600699
rect 675507 600643 675563 600699
rect 675587 600643 675643 600699
rect 675667 600643 675723 600699
rect 675427 600091 675483 600147
rect 675507 600091 675563 600147
rect 675587 600091 675643 600147
rect 675667 600091 675723 600147
rect 675427 599447 675483 599503
rect 675507 599447 675563 599503
rect 675587 599447 675643 599503
rect 675667 599447 675723 599503
rect 675427 598803 675483 598859
rect 675507 598803 675563 598859
rect 675587 598803 675643 598859
rect 675667 598803 675723 598859
rect 675427 597607 675483 597663
rect 675507 597607 675563 597663
rect 675587 597607 675643 597663
rect 675667 597607 675723 597663
rect 675427 596411 675483 596467
rect 675507 596411 675563 596467
rect 675587 596411 675643 596467
rect 675667 596411 675723 596467
rect 675427 595767 675483 595823
rect 675507 595767 675563 595823
rect 675587 595767 675643 595823
rect 675667 595767 675723 595823
rect 675427 595123 675483 595179
rect 675507 595123 675563 595179
rect 675587 595123 675643 595179
rect 675667 595123 675723 595179
rect 675427 593927 675483 593983
rect 675507 593927 675563 593983
rect 675587 593927 675643 593983
rect 675667 593927 675723 593983
rect 41883 583417 41939 583473
rect 41963 583417 42019 583473
rect 42043 583417 42099 583473
rect 42123 583417 42179 583473
rect 41883 582221 41939 582277
rect 41963 582221 42019 582277
rect 42043 582221 42099 582277
rect 42123 582221 42179 582277
rect 41883 581577 41939 581633
rect 41963 581577 42019 581633
rect 42043 581577 42099 581633
rect 42123 581577 42179 581633
rect 41883 580933 41939 580989
rect 41963 580933 42019 580989
rect 42043 580933 42099 580989
rect 42123 580933 42179 580989
rect 41883 579737 41939 579793
rect 41963 579737 42019 579793
rect 42043 579737 42099 579793
rect 42123 579737 42179 579793
rect 41883 578541 41939 578597
rect 41963 578541 42019 578597
rect 42043 578541 42099 578597
rect 42123 578541 42179 578597
rect 41883 577897 41939 577953
rect 41963 577897 42019 577953
rect 42043 577897 42099 577953
rect 42123 577897 42179 577953
rect 41883 577253 41939 577309
rect 41963 577253 42019 577309
rect 42043 577253 42099 577309
rect 42123 577253 42179 577309
rect 41883 576701 41939 576757
rect 41963 576701 42019 576757
rect 42043 576701 42099 576757
rect 42123 576701 42179 576757
rect 41883 574217 41939 574273
rect 41963 574217 42019 574273
rect 42043 574217 42099 574273
rect 42123 574217 42179 574273
rect 41883 573573 41939 573629
rect 41963 573573 42019 573629
rect 42043 573573 42099 573629
rect 42123 573573 42179 573629
rect 41883 572929 41939 572985
rect 41963 572929 42019 572985
rect 42043 572929 42099 572985
rect 42123 572929 42179 572985
rect 41883 572377 41939 572433
rect 41963 572377 42019 572433
rect 42043 572377 42099 572433
rect 42123 572377 42179 572433
rect 41883 570537 41939 570593
rect 41963 570537 42019 570593
rect 42043 570537 42099 570593
rect 42123 570537 42179 570593
rect 41883 569893 41939 569949
rect 41963 569893 42019 569949
rect 42043 569893 42099 569949
rect 42123 569893 42179 569949
rect 41883 569249 41939 569305
rect 41963 569249 42019 569305
rect 42043 569249 42099 569305
rect 42123 569249 42179 569305
rect 675427 562895 675483 562951
rect 675507 562895 675563 562951
rect 675587 562895 675643 562951
rect 675667 562895 675723 562951
rect 675427 562251 675483 562307
rect 675507 562251 675563 562307
rect 675587 562251 675643 562307
rect 675667 562251 675723 562307
rect 675427 561607 675483 561663
rect 675507 561607 675563 561663
rect 675587 561607 675643 561663
rect 675667 561607 675723 561663
rect 675427 559767 675483 559823
rect 675507 559767 675563 559823
rect 675587 559767 675643 559823
rect 675667 559767 675723 559823
rect 675427 559215 675483 559271
rect 675507 559215 675563 559271
rect 675587 559215 675643 559271
rect 675667 559215 675723 559271
rect 675427 558571 675483 558627
rect 675507 558571 675563 558627
rect 675587 558571 675643 558627
rect 675667 558571 675723 558627
rect 675427 557927 675483 557983
rect 675507 557927 675563 557983
rect 675587 557927 675643 557983
rect 675667 557927 675723 557983
rect 675427 555443 675483 555499
rect 675507 555443 675563 555499
rect 675587 555443 675643 555499
rect 675667 555443 675723 555499
rect 675427 554891 675483 554947
rect 675507 554891 675563 554947
rect 675587 554891 675643 554947
rect 675667 554891 675723 554947
rect 675427 554247 675483 554303
rect 675507 554247 675563 554303
rect 675587 554247 675643 554303
rect 675667 554247 675723 554303
rect 675427 553603 675483 553659
rect 675507 553603 675563 553659
rect 675587 553603 675643 553659
rect 675667 553603 675723 553659
rect 675427 552407 675483 552463
rect 675507 552407 675563 552463
rect 675587 552407 675643 552463
rect 675667 552407 675723 552463
rect 675427 551211 675483 551267
rect 675507 551211 675563 551267
rect 675587 551211 675643 551267
rect 675667 551211 675723 551267
rect 675427 550567 675483 550623
rect 675507 550567 675563 550623
rect 675587 550567 675643 550623
rect 675667 550567 675723 550623
rect 675427 549923 675483 549979
rect 675507 549923 675563 549979
rect 675587 549923 675643 549979
rect 675667 549923 675723 549979
rect 675427 548727 675483 548783
rect 675507 548727 675563 548783
rect 675587 548727 675643 548783
rect 675667 548727 675723 548783
rect 41883 540217 41939 540273
rect 41963 540217 42019 540273
rect 42043 540217 42099 540273
rect 42123 540217 42179 540273
rect 41883 539021 41939 539077
rect 41963 539021 42019 539077
rect 42043 539021 42099 539077
rect 42123 539021 42179 539077
rect 41883 538377 41939 538433
rect 41963 538377 42019 538433
rect 42043 538377 42099 538433
rect 42123 538377 42179 538433
rect 41883 537733 41939 537789
rect 41963 537733 42019 537789
rect 42043 537733 42099 537789
rect 42123 537733 42179 537789
rect 41883 536537 41939 536593
rect 41963 536537 42019 536593
rect 42043 536537 42099 536593
rect 42123 536537 42179 536593
rect 41883 535341 41939 535397
rect 41963 535341 42019 535397
rect 42043 535341 42099 535397
rect 42123 535341 42179 535397
rect 41883 534697 41939 534753
rect 41963 534697 42019 534753
rect 42043 534697 42099 534753
rect 42123 534697 42179 534753
rect 41883 534053 41939 534109
rect 41963 534053 42019 534109
rect 42043 534053 42099 534109
rect 42123 534053 42179 534109
rect 41883 533501 41939 533557
rect 41963 533501 42019 533557
rect 42043 533501 42099 533557
rect 42123 533501 42179 533557
rect 41883 531017 41939 531073
rect 41963 531017 42019 531073
rect 42043 531017 42099 531073
rect 42123 531017 42179 531073
rect 41883 530373 41939 530429
rect 41963 530373 42019 530429
rect 42043 530373 42099 530429
rect 42123 530373 42179 530429
rect 41883 529729 41939 529785
rect 41963 529729 42019 529785
rect 42043 529729 42099 529785
rect 42123 529729 42179 529785
rect 41883 529177 41939 529233
rect 41963 529177 42019 529233
rect 42043 529177 42099 529233
rect 42123 529177 42179 529233
rect 41883 527337 41939 527393
rect 41963 527337 42019 527393
rect 42043 527337 42099 527393
rect 42123 527337 42179 527393
rect 41883 526693 41939 526749
rect 41963 526693 42019 526749
rect 42043 526693 42099 526749
rect 42123 526693 42179 526749
rect 41883 526049 41939 526105
rect 41963 526049 42019 526105
rect 42043 526049 42099 526105
rect 42123 526049 42179 526105
rect 41883 412617 41939 412673
rect 41963 412617 42019 412673
rect 42043 412617 42099 412673
rect 42123 412617 42179 412673
rect 41883 411421 41939 411477
rect 41963 411421 42019 411477
rect 42043 411421 42099 411477
rect 42123 411421 42179 411477
rect 41883 410777 41939 410833
rect 41963 410777 42019 410833
rect 42043 410777 42099 410833
rect 42123 410777 42179 410833
rect 41883 410133 41939 410189
rect 41963 410133 42019 410189
rect 42043 410133 42099 410189
rect 42123 410133 42179 410189
rect 41883 408937 41939 408993
rect 41963 408937 42019 408993
rect 42043 408937 42099 408993
rect 42123 408937 42179 408993
rect 41883 407741 41939 407797
rect 41963 407741 42019 407797
rect 42043 407741 42099 407797
rect 42123 407741 42179 407797
rect 41883 407097 41939 407153
rect 41963 407097 42019 407153
rect 42043 407097 42099 407153
rect 42123 407097 42179 407153
rect 41883 406453 41939 406509
rect 41963 406453 42019 406509
rect 42043 406453 42099 406509
rect 42123 406453 42179 406509
rect 41883 405901 41939 405957
rect 41963 405901 42019 405957
rect 42043 405901 42099 405957
rect 42123 405901 42179 405957
rect 41883 403417 41939 403473
rect 41963 403417 42019 403473
rect 42043 403417 42099 403473
rect 42123 403417 42179 403473
rect 41883 402773 41939 402829
rect 41963 402773 42019 402829
rect 42043 402773 42099 402829
rect 42123 402773 42179 402829
rect 41883 402129 41939 402185
rect 41963 402129 42019 402185
rect 42043 402129 42099 402185
rect 42123 402129 42179 402185
rect 41883 401577 41939 401633
rect 41963 401577 42019 401633
rect 42043 401577 42099 401633
rect 42123 401577 42179 401633
rect 41883 399737 41939 399793
rect 41963 399737 42019 399793
rect 42043 399737 42099 399793
rect 42123 399737 42179 399793
rect 41883 399093 41939 399149
rect 41963 399093 42019 399149
rect 42043 399093 42099 399149
rect 42123 399093 42179 399149
rect 41883 398449 41939 398505
rect 41963 398449 42019 398505
rect 42043 398449 42099 398505
rect 42123 398449 42179 398505
rect 675427 385695 675483 385751
rect 675507 385695 675563 385751
rect 675587 385695 675643 385751
rect 675667 385695 675723 385751
rect 675427 385051 675483 385107
rect 675507 385051 675563 385107
rect 675587 385051 675643 385107
rect 675667 385051 675723 385107
rect 675427 384407 675483 384463
rect 675507 384407 675563 384463
rect 675587 384407 675643 384463
rect 675667 384407 675723 384463
rect 675427 382567 675483 382623
rect 675507 382567 675563 382623
rect 675587 382567 675643 382623
rect 675667 382567 675723 382623
rect 675427 382015 675483 382071
rect 675507 382015 675563 382071
rect 675587 382015 675643 382071
rect 675667 382015 675723 382071
rect 675427 381371 675483 381427
rect 675507 381371 675563 381427
rect 675587 381371 675643 381427
rect 675667 381371 675723 381427
rect 675427 380727 675483 380783
rect 675507 380727 675563 380783
rect 675587 380727 675643 380783
rect 675667 380727 675723 380783
rect 675427 378243 675483 378299
rect 675507 378243 675563 378299
rect 675587 378243 675643 378299
rect 675667 378243 675723 378299
rect 675427 377691 675483 377747
rect 675507 377691 675563 377747
rect 675587 377691 675643 377747
rect 675667 377691 675723 377747
rect 675427 377047 675483 377103
rect 675507 377047 675563 377103
rect 675587 377047 675643 377103
rect 675667 377047 675723 377103
rect 675427 376403 675483 376459
rect 675507 376403 675563 376459
rect 675587 376403 675643 376459
rect 675667 376403 675723 376459
rect 675427 375207 675483 375263
rect 675507 375207 675563 375263
rect 675587 375207 675643 375263
rect 675667 375207 675723 375263
rect 675427 373367 675483 373423
rect 675507 373367 675563 373423
rect 675587 373367 675643 373423
rect 675667 373367 675723 373423
rect 675427 372723 675483 372779
rect 675507 372723 675563 372779
rect 675587 372723 675643 372779
rect 675667 372723 675723 372779
rect 675427 371527 675483 371583
rect 675507 371527 675563 371583
rect 675587 371527 675643 371583
rect 675667 371527 675723 371583
rect 41883 369417 41939 369473
rect 41963 369417 42019 369473
rect 42043 369417 42099 369473
rect 42123 369417 42179 369473
rect 41883 368221 41939 368277
rect 41963 368221 42019 368277
rect 42043 368221 42099 368277
rect 42123 368221 42179 368277
rect 41883 367577 41939 367633
rect 41963 367577 42019 367633
rect 42043 367577 42099 367633
rect 42123 367577 42179 367633
rect 41883 366933 41939 366989
rect 41963 366933 42019 366989
rect 42043 366933 42099 366989
rect 42123 366933 42179 366989
rect 41883 365737 41939 365793
rect 41963 365737 42019 365793
rect 42043 365737 42099 365793
rect 42123 365737 42179 365793
rect 41883 364541 41939 364597
rect 41963 364541 42019 364597
rect 42043 364541 42099 364597
rect 42123 364541 42179 364597
rect 41883 363897 41939 363953
rect 41963 363897 42019 363953
rect 42043 363897 42099 363953
rect 42123 363897 42179 363953
rect 41883 363253 41939 363309
rect 41963 363253 42019 363309
rect 42043 363253 42099 363309
rect 42123 363253 42179 363309
rect 41883 362701 41939 362757
rect 41963 362701 42019 362757
rect 42043 362701 42099 362757
rect 42123 362701 42179 362757
rect 41883 360217 41939 360273
rect 41963 360217 42019 360273
rect 42043 360217 42099 360273
rect 42123 360217 42179 360273
rect 41883 359573 41939 359629
rect 41963 359573 42019 359629
rect 42043 359573 42099 359629
rect 42123 359573 42179 359629
rect 41883 358929 41939 358985
rect 41963 358929 42019 358985
rect 42043 358929 42099 358985
rect 42123 358929 42179 358985
rect 41883 358377 41939 358433
rect 41963 358377 42019 358433
rect 42043 358377 42099 358433
rect 42123 358377 42179 358433
rect 41883 356537 41939 356593
rect 41963 356537 42019 356593
rect 42043 356537 42099 356593
rect 42123 356537 42179 356593
rect 41883 355893 41939 355949
rect 41963 355893 42019 355949
rect 42043 355893 42099 355949
rect 42123 355893 42179 355949
rect 41883 355249 41939 355305
rect 41963 355249 42019 355305
rect 42043 355249 42099 355305
rect 42123 355249 42179 355305
rect 675427 340495 675483 340551
rect 675507 340495 675563 340551
rect 675587 340495 675643 340551
rect 675667 340495 675723 340551
rect 675427 339851 675483 339907
rect 675507 339851 675563 339907
rect 675587 339851 675643 339907
rect 675667 339851 675723 339907
rect 675427 339207 675483 339263
rect 675507 339207 675563 339263
rect 675587 339207 675643 339263
rect 675667 339207 675723 339263
rect 675427 337367 675483 337423
rect 675507 337367 675563 337423
rect 675587 337367 675643 337423
rect 675667 337367 675723 337423
rect 675427 336815 675483 336871
rect 675507 336815 675563 336871
rect 675587 336815 675643 336871
rect 675667 336815 675723 336871
rect 675427 336171 675483 336227
rect 675507 336171 675563 336227
rect 675587 336171 675643 336227
rect 675667 336171 675723 336227
rect 675427 335527 675483 335583
rect 675507 335527 675563 335583
rect 675587 335527 675643 335583
rect 675667 335527 675723 335583
rect 675427 333043 675483 333099
rect 675507 333043 675563 333099
rect 675587 333043 675643 333099
rect 675667 333043 675723 333099
rect 675427 332491 675483 332547
rect 675507 332491 675563 332547
rect 675587 332491 675643 332547
rect 675667 332491 675723 332547
rect 675427 331847 675483 331903
rect 675507 331847 675563 331903
rect 675587 331847 675643 331903
rect 675667 331847 675723 331903
rect 675427 331203 675483 331259
rect 675507 331203 675563 331259
rect 675587 331203 675643 331259
rect 675667 331203 675723 331259
rect 675427 330007 675483 330063
rect 675507 330007 675563 330063
rect 675587 330007 675643 330063
rect 675667 330007 675723 330063
rect 675427 328167 675483 328223
rect 675507 328167 675563 328223
rect 675587 328167 675643 328223
rect 675667 328167 675723 328223
rect 675427 327523 675483 327579
rect 675507 327523 675563 327579
rect 675587 327523 675643 327579
rect 675667 327523 675723 327579
rect 675427 326327 675483 326383
rect 675507 326327 675563 326383
rect 675587 326327 675643 326383
rect 675667 326327 675723 326383
rect 41883 326217 41939 326273
rect 41963 326217 42019 326273
rect 42043 326217 42099 326273
rect 42123 326217 42179 326273
rect 41883 325021 41939 325077
rect 41963 325021 42019 325077
rect 42043 325021 42099 325077
rect 42123 325021 42179 325077
rect 41883 324377 41939 324433
rect 41963 324377 42019 324433
rect 42043 324377 42099 324433
rect 42123 324377 42179 324433
rect 41883 323733 41939 323789
rect 41963 323733 42019 323789
rect 42043 323733 42099 323789
rect 42123 323733 42179 323789
rect 41883 322537 41939 322593
rect 41963 322537 42019 322593
rect 42043 322537 42099 322593
rect 42123 322537 42179 322593
rect 41883 321341 41939 321397
rect 41963 321341 42019 321397
rect 42043 321341 42099 321397
rect 42123 321341 42179 321397
rect 41883 320697 41939 320753
rect 41963 320697 42019 320753
rect 42043 320697 42099 320753
rect 42123 320697 42179 320753
rect 41883 320053 41939 320109
rect 41963 320053 42019 320109
rect 42043 320053 42099 320109
rect 42123 320053 42179 320109
rect 41883 319501 41939 319557
rect 41963 319501 42019 319557
rect 42043 319501 42099 319557
rect 42123 319501 42179 319557
rect 41883 317017 41939 317073
rect 41963 317017 42019 317073
rect 42043 317017 42099 317073
rect 42123 317017 42179 317073
rect 41883 316373 41939 316429
rect 41963 316373 42019 316429
rect 42043 316373 42099 316429
rect 42123 316373 42179 316429
rect 41883 315729 41939 315785
rect 41963 315729 42019 315785
rect 42043 315729 42099 315785
rect 42123 315729 42179 315785
rect 41883 315177 41939 315233
rect 41963 315177 42019 315233
rect 42043 315177 42099 315233
rect 42123 315177 42179 315233
rect 41883 313337 41939 313393
rect 41963 313337 42019 313393
rect 42043 313337 42099 313393
rect 42123 313337 42179 313393
rect 41883 312693 41939 312749
rect 41963 312693 42019 312749
rect 42043 312693 42099 312749
rect 42123 312693 42179 312749
rect 41883 312049 41939 312105
rect 41963 312049 42019 312105
rect 42043 312049 42099 312105
rect 42123 312049 42179 312105
rect 675427 295495 675483 295551
rect 675507 295495 675563 295551
rect 675587 295495 675643 295551
rect 675667 295495 675723 295551
rect 675427 294851 675483 294907
rect 675507 294851 675563 294907
rect 675587 294851 675643 294907
rect 675667 294851 675723 294907
rect 675427 294207 675483 294263
rect 675507 294207 675563 294263
rect 675587 294207 675643 294263
rect 675667 294207 675723 294263
rect 675427 292367 675483 292423
rect 675507 292367 675563 292423
rect 675587 292367 675643 292423
rect 675667 292367 675723 292423
rect 675427 291815 675483 291871
rect 675507 291815 675563 291871
rect 675587 291815 675643 291871
rect 675667 291815 675723 291871
rect 675427 291171 675483 291227
rect 675507 291171 675563 291227
rect 675587 291171 675643 291227
rect 675667 291171 675723 291227
rect 675427 290527 675483 290583
rect 675507 290527 675563 290583
rect 675587 290527 675643 290583
rect 675667 290527 675723 290583
rect 675427 288043 675483 288099
rect 675507 288043 675563 288099
rect 675587 288043 675643 288099
rect 675667 288043 675723 288099
rect 675427 287491 675483 287547
rect 675507 287491 675563 287547
rect 675587 287491 675643 287547
rect 675667 287491 675723 287547
rect 675427 286847 675483 286903
rect 675507 286847 675563 286903
rect 675587 286847 675643 286903
rect 675667 286847 675723 286903
rect 675427 286203 675483 286259
rect 675507 286203 675563 286259
rect 675587 286203 675643 286259
rect 675667 286203 675723 286259
rect 675427 285007 675483 285063
rect 675507 285007 675563 285063
rect 675587 285007 675643 285063
rect 675667 285007 675723 285063
rect 675427 283167 675483 283223
rect 675507 283167 675563 283223
rect 675587 283167 675643 283223
rect 675667 283167 675723 283223
rect 41883 283017 41939 283073
rect 41963 283017 42019 283073
rect 42043 283017 42099 283073
rect 42123 283017 42179 283073
rect 675427 282523 675483 282579
rect 675507 282523 675563 282579
rect 675587 282523 675643 282579
rect 675667 282523 675723 282579
rect 41883 281821 41939 281877
rect 41963 281821 42019 281877
rect 42043 281821 42099 281877
rect 42123 281821 42179 281877
rect 675427 281327 675483 281383
rect 675507 281327 675563 281383
rect 675587 281327 675643 281383
rect 675667 281327 675723 281383
rect 41883 281177 41939 281233
rect 41963 281177 42019 281233
rect 42043 281177 42099 281233
rect 42123 281177 42179 281233
rect 41883 280533 41939 280589
rect 41963 280533 42019 280589
rect 42043 280533 42099 280589
rect 42123 280533 42179 280589
rect 41883 279337 41939 279393
rect 41963 279337 42019 279393
rect 42043 279337 42099 279393
rect 42123 279337 42179 279393
rect 41883 278141 41939 278197
rect 41963 278141 42019 278197
rect 42043 278141 42099 278197
rect 42123 278141 42179 278197
rect 41883 277497 41939 277553
rect 41963 277497 42019 277553
rect 42043 277497 42099 277553
rect 42123 277497 42179 277553
rect 41883 276853 41939 276909
rect 41963 276853 42019 276909
rect 42043 276853 42099 276909
rect 42123 276853 42179 276909
rect 41883 276301 41939 276357
rect 41963 276301 42019 276357
rect 42043 276301 42099 276357
rect 42123 276301 42179 276357
rect 41883 273817 41939 273873
rect 41963 273817 42019 273873
rect 42043 273817 42099 273873
rect 42123 273817 42179 273873
rect 41883 273173 41939 273229
rect 41963 273173 42019 273229
rect 42043 273173 42099 273229
rect 42123 273173 42179 273229
rect 41883 272529 41939 272585
rect 41963 272529 42019 272585
rect 42043 272529 42099 272585
rect 42123 272529 42179 272585
rect 41883 271977 41939 272033
rect 41963 271977 42019 272033
rect 42043 271977 42099 272033
rect 42123 271977 42179 272033
rect 41883 270137 41939 270193
rect 41963 270137 42019 270193
rect 42043 270137 42099 270193
rect 42123 270137 42179 270193
rect 41883 269493 41939 269549
rect 41963 269493 42019 269549
rect 42043 269493 42099 269549
rect 42123 269493 42179 269549
rect 41883 268849 41939 268905
rect 41963 268849 42019 268905
rect 42043 268849 42099 268905
rect 42123 268849 42179 268905
rect 675427 250495 675483 250551
rect 675507 250495 675563 250551
rect 675587 250495 675643 250551
rect 675667 250495 675723 250551
rect 675427 249851 675483 249907
rect 675507 249851 675563 249907
rect 675587 249851 675643 249907
rect 675667 249851 675723 249907
rect 675427 249207 675483 249263
rect 675507 249207 675563 249263
rect 675587 249207 675643 249263
rect 675667 249207 675723 249263
rect 675427 247367 675483 247423
rect 675507 247367 675563 247423
rect 675587 247367 675643 247423
rect 675667 247367 675723 247423
rect 675427 246815 675483 246871
rect 675507 246815 675563 246871
rect 675587 246815 675643 246871
rect 675667 246815 675723 246871
rect 675427 246171 675483 246227
rect 675507 246171 675563 246227
rect 675587 246171 675643 246227
rect 675667 246171 675723 246227
rect 675427 245527 675483 245583
rect 675507 245527 675563 245583
rect 675587 245527 675643 245583
rect 675667 245527 675723 245583
rect 675427 243043 675483 243099
rect 675507 243043 675563 243099
rect 675587 243043 675643 243099
rect 675667 243043 675723 243099
rect 675427 242491 675483 242547
rect 675507 242491 675563 242547
rect 675587 242491 675643 242547
rect 675667 242491 675723 242547
rect 675427 241847 675483 241903
rect 675507 241847 675563 241903
rect 675587 241847 675643 241903
rect 675667 241847 675723 241903
rect 675427 241203 675483 241259
rect 675507 241203 675563 241259
rect 675587 241203 675643 241259
rect 675667 241203 675723 241259
rect 675427 240007 675483 240063
rect 675507 240007 675563 240063
rect 675587 240007 675643 240063
rect 675667 240007 675723 240063
rect 41883 239817 41939 239873
rect 41963 239817 42019 239873
rect 42043 239817 42099 239873
rect 42123 239817 42179 239873
rect 41883 238621 41939 238677
rect 41963 238621 42019 238677
rect 42043 238621 42099 238677
rect 42123 238621 42179 238677
rect 675427 238167 675483 238223
rect 675507 238167 675563 238223
rect 675587 238167 675643 238223
rect 675667 238167 675723 238223
rect 41883 237977 41939 238033
rect 41963 237977 42019 238033
rect 42043 237977 42099 238033
rect 42123 237977 42179 238033
rect 675427 237523 675483 237579
rect 675507 237523 675563 237579
rect 675587 237523 675643 237579
rect 675667 237523 675723 237579
rect 675427 236327 675483 236383
rect 675507 236327 675563 236383
rect 675587 236327 675643 236383
rect 675667 236327 675723 236383
rect 41883 236137 41939 236193
rect 41963 236137 42019 236193
rect 42043 236137 42099 236193
rect 42123 236137 42179 236193
rect 41883 234941 41939 234997
rect 41963 234941 42019 234997
rect 42043 234941 42099 234997
rect 42123 234941 42179 234997
rect 41883 234297 41939 234353
rect 41963 234297 42019 234353
rect 42043 234297 42099 234353
rect 42123 234297 42179 234353
rect 41883 233653 41939 233709
rect 41963 233653 42019 233709
rect 42043 233653 42099 233709
rect 42123 233653 42179 233709
rect 41883 233101 41939 233157
rect 41963 233101 42019 233157
rect 42043 233101 42099 233157
rect 42123 233101 42179 233157
rect 41883 230617 41939 230673
rect 41963 230617 42019 230673
rect 42043 230617 42099 230673
rect 42123 230617 42179 230673
rect 41883 229973 41939 230029
rect 41963 229973 42019 230029
rect 42043 229973 42099 230029
rect 42123 229973 42179 230029
rect 41883 229329 41939 229385
rect 41963 229329 42019 229385
rect 42043 229329 42099 229385
rect 42123 229329 42179 229385
rect 41883 228777 41939 228833
rect 41963 228777 42019 228833
rect 42043 228777 42099 228833
rect 42123 228777 42179 228833
rect 41883 226937 41939 226993
rect 41963 226937 42019 226993
rect 42043 226937 42099 226993
rect 42123 226937 42179 226993
rect 41883 226293 41939 226349
rect 41963 226293 42019 226349
rect 42043 226293 42099 226349
rect 42123 226293 42179 226349
rect 41883 225649 41939 225705
rect 41963 225649 42019 225705
rect 42043 225649 42099 225705
rect 42123 225649 42179 225705
rect 675427 205295 675483 205351
rect 675507 205295 675563 205351
rect 675587 205295 675643 205351
rect 675667 205295 675723 205351
rect 675427 204651 675483 204707
rect 675507 204651 675563 204707
rect 675587 204651 675643 204707
rect 675667 204651 675723 204707
rect 675427 204007 675483 204063
rect 675507 204007 675563 204063
rect 675587 204007 675643 204063
rect 675667 204007 675723 204063
rect 675427 202167 675483 202223
rect 675507 202167 675563 202223
rect 675587 202167 675643 202223
rect 675667 202167 675723 202223
rect 675427 201615 675483 201671
rect 675507 201615 675563 201671
rect 675587 201615 675643 201671
rect 675667 201615 675723 201671
rect 675427 200971 675483 201027
rect 675507 200971 675563 201027
rect 675587 200971 675643 201027
rect 675667 200971 675723 201027
rect 675427 200327 675483 200383
rect 675507 200327 675563 200383
rect 675587 200327 675643 200383
rect 675667 200327 675723 200383
rect 675427 197843 675483 197899
rect 675507 197843 675563 197899
rect 675587 197843 675643 197899
rect 675667 197843 675723 197899
rect 675427 197291 675483 197347
rect 675507 197291 675563 197347
rect 675587 197291 675643 197347
rect 675667 197291 675723 197347
rect 41883 196617 41939 196673
rect 41963 196617 42019 196673
rect 42043 196617 42099 196673
rect 42123 196617 42179 196673
rect 675427 196647 675483 196703
rect 675507 196647 675563 196703
rect 675587 196647 675643 196703
rect 675667 196647 675723 196703
rect 675427 196003 675483 196059
rect 675507 196003 675563 196059
rect 675587 196003 675643 196059
rect 675667 196003 675723 196059
rect 41883 195421 41939 195477
rect 41963 195421 42019 195477
rect 42043 195421 42099 195477
rect 42123 195421 42179 195477
rect 41883 194777 41939 194833
rect 41963 194777 42019 194833
rect 42043 194777 42099 194833
rect 42123 194777 42179 194833
rect 675427 194807 675483 194863
rect 675507 194807 675563 194863
rect 675587 194807 675643 194863
rect 675667 194807 675723 194863
rect 41883 192937 41939 192993
rect 41963 192937 42019 192993
rect 42043 192937 42099 192993
rect 42123 192937 42179 192993
rect 675427 192967 675483 193023
rect 675507 192967 675563 193023
rect 675587 192967 675643 193023
rect 675667 192967 675723 193023
rect 675427 192323 675483 192379
rect 675507 192323 675563 192379
rect 675587 192323 675643 192379
rect 675667 192323 675723 192379
rect 41883 191741 41939 191797
rect 41963 191741 42019 191797
rect 42043 191741 42099 191797
rect 42123 191741 42179 191797
rect 41883 191097 41939 191153
rect 41963 191097 42019 191153
rect 42043 191097 42099 191153
rect 42123 191097 42179 191153
rect 675427 191127 675483 191183
rect 675507 191127 675563 191183
rect 675587 191127 675643 191183
rect 675667 191127 675723 191183
rect 41883 190453 41939 190509
rect 41963 190453 42019 190509
rect 42043 190453 42099 190509
rect 42123 190453 42179 190509
rect 41883 189901 41939 189957
rect 41963 189901 42019 189957
rect 42043 189901 42099 189957
rect 42123 189901 42179 189957
rect 41883 187417 41939 187473
rect 41963 187417 42019 187473
rect 42043 187417 42099 187473
rect 42123 187417 42179 187473
rect 41883 186773 41939 186829
rect 41963 186773 42019 186829
rect 42043 186773 42099 186829
rect 42123 186773 42179 186829
rect 41883 186129 41939 186185
rect 41963 186129 42019 186185
rect 42043 186129 42099 186185
rect 42123 186129 42179 186185
rect 41883 185577 41939 185633
rect 41963 185577 42019 185633
rect 42043 185577 42099 185633
rect 42123 185577 42179 185633
rect 41883 183737 41939 183793
rect 41963 183737 42019 183793
rect 42043 183737 42099 183793
rect 42123 183737 42179 183793
rect 41883 183093 41939 183149
rect 41963 183093 42019 183149
rect 42043 183093 42099 183149
rect 42123 183093 42179 183149
rect 41883 182449 41939 182505
rect 41963 182449 42019 182505
rect 42043 182449 42099 182505
rect 42123 182449 42179 182505
rect 675427 160295 675483 160351
rect 675507 160295 675563 160351
rect 675587 160295 675643 160351
rect 675667 160295 675723 160351
rect 675427 159651 675483 159707
rect 675507 159651 675563 159707
rect 675587 159651 675643 159707
rect 675667 159651 675723 159707
rect 675427 159007 675483 159063
rect 675507 159007 675563 159063
rect 675587 159007 675643 159063
rect 675667 159007 675723 159063
rect 675427 157167 675483 157223
rect 675507 157167 675563 157223
rect 675587 157167 675643 157223
rect 675667 157167 675723 157223
rect 675427 156615 675483 156671
rect 675507 156615 675563 156671
rect 675587 156615 675643 156671
rect 675667 156615 675723 156671
rect 675427 155971 675483 156027
rect 675507 155971 675563 156027
rect 675587 155971 675643 156027
rect 675667 155971 675723 156027
rect 675427 155327 675483 155383
rect 675507 155327 675563 155383
rect 675587 155327 675643 155383
rect 675667 155327 675723 155383
rect 675427 152843 675483 152899
rect 675507 152843 675563 152899
rect 675587 152843 675643 152899
rect 675667 152843 675723 152899
rect 675427 152291 675483 152347
rect 675507 152291 675563 152347
rect 675587 152291 675643 152347
rect 675667 152291 675723 152347
rect 675427 151647 675483 151703
rect 675507 151647 675563 151703
rect 675587 151647 675643 151703
rect 675667 151647 675723 151703
rect 675427 151003 675483 151059
rect 675507 151003 675563 151059
rect 675587 151003 675643 151059
rect 675667 151003 675723 151059
rect 675427 149807 675483 149863
rect 675507 149807 675563 149863
rect 675587 149807 675643 149863
rect 675667 149807 675723 149863
rect 675427 147967 675483 148023
rect 675507 147967 675563 148023
rect 675587 147967 675643 148023
rect 675667 147967 675723 148023
rect 675427 147323 675483 147379
rect 675507 147323 675563 147379
rect 675587 147323 675643 147379
rect 675667 147323 675723 147379
rect 675427 146127 675483 146183
rect 675507 146127 675563 146183
rect 675587 146127 675643 146183
rect 675667 146127 675723 146183
rect 675427 115095 675483 115151
rect 675507 115095 675563 115151
rect 675587 115095 675643 115151
rect 675667 115095 675723 115151
rect 675427 114451 675483 114507
rect 675507 114451 675563 114507
rect 675587 114451 675643 114507
rect 675667 114451 675723 114507
rect 675427 113807 675483 113863
rect 675507 113807 675563 113863
rect 675587 113807 675643 113863
rect 675667 113807 675723 113863
rect 675427 111967 675483 112023
rect 675507 111967 675563 112023
rect 675587 111967 675643 112023
rect 675667 111967 675723 112023
rect 675427 111415 675483 111471
rect 675507 111415 675563 111471
rect 675587 111415 675643 111471
rect 675667 111415 675723 111471
rect 675427 110771 675483 110827
rect 675507 110771 675563 110827
rect 675587 110771 675643 110827
rect 675667 110771 675723 110827
rect 675427 110127 675483 110183
rect 675507 110127 675563 110183
rect 675587 110127 675643 110183
rect 675667 110127 675723 110183
rect 675427 107643 675483 107699
rect 675507 107643 675563 107699
rect 675587 107643 675643 107699
rect 675667 107643 675723 107699
rect 675427 107091 675483 107147
rect 675507 107091 675563 107147
rect 675587 107091 675643 107147
rect 675667 107091 675723 107147
rect 675427 106447 675483 106503
rect 675507 106447 675563 106503
rect 675587 106447 675643 106503
rect 675667 106447 675723 106503
rect 675427 105803 675483 105859
rect 675507 105803 675563 105859
rect 675587 105803 675643 105859
rect 675667 105803 675723 105859
rect 675427 104607 675483 104663
rect 675507 104607 675563 104663
rect 675587 104607 675643 104663
rect 675667 104607 675723 104663
rect 675427 102767 675483 102823
rect 675507 102767 675563 102823
rect 675587 102767 675643 102823
rect 675667 102767 675723 102823
rect 675427 102123 675483 102179
rect 675507 102123 675563 102179
rect 675587 102123 675643 102179
rect 675667 102123 675723 102179
rect 675427 100927 675483 100983
rect 675507 100927 675563 100983
rect 675587 100927 675643 100983
rect 675667 100927 675723 100983
rect 143435 40073 143437 40090
rect 143437 40073 143489 40090
rect 143489 40073 143491 40090
rect 143435 40034 143491 40073
rect 145830 40916 145886 40972
rect 202715 40915 202771 40971
rect 205926 40914 205982 40970
rect 311315 40915 311371 40971
rect 315495 40918 315551 40974
rect 366115 40915 366171 40971
rect 370300 40914 370356 40970
rect 420915 40915 420971 40971
rect 425113 40902 425169 40958
rect 475715 40915 475771 40971
rect 479913 40916 479969 40972
rect 530515 40915 530571 40971
rect 534770 40904 534826 40960
rect 145839 40076 145895 40132
<< metal3 >>
rect 41863 969273 42193 969280
rect 41863 969217 41883 969273
rect 41939 969217 41963 969273
rect 42019 969217 42043 969273
rect 42099 969217 42123 969273
rect 42179 969217 42193 969273
rect 41863 969210 42193 969217
rect 41863 968077 42193 968084
rect 41863 968021 41883 968077
rect 41939 968021 41963 968077
rect 42019 968021 42043 968077
rect 42099 968021 42123 968077
rect 42179 968021 42193 968077
rect 41863 968014 42193 968021
rect 41863 967433 42193 967440
rect 41863 967377 41883 967433
rect 41939 967377 41963 967433
rect 42019 967377 42043 967433
rect 42099 967377 42123 967433
rect 42179 967377 42193 967433
rect 41863 967370 42193 967377
rect 41863 966789 42193 966796
rect 41863 966733 41883 966789
rect 41939 966733 41963 966789
rect 42019 966733 42043 966789
rect 42099 966733 42123 966789
rect 42179 966733 42193 966789
rect 41863 966726 42193 966733
rect 675407 966751 675737 966758
rect 675407 966695 675427 966751
rect 675483 966695 675507 966751
rect 675563 966695 675587 966751
rect 675643 966695 675667 966751
rect 675723 966695 675737 966751
rect 675407 966688 675737 966695
rect 675407 966107 675737 966114
rect 675407 966051 675427 966107
rect 675483 966051 675507 966107
rect 675563 966051 675587 966107
rect 675643 966051 675667 966107
rect 675723 966051 675737 966107
rect 675407 966044 675737 966051
rect 41863 965593 42193 965600
rect 41863 965537 41883 965593
rect 41939 965537 41963 965593
rect 42019 965537 42043 965593
rect 42099 965537 42123 965593
rect 42179 965537 42193 965593
rect 41863 965530 42193 965537
rect 675407 965463 675737 965470
rect 675407 965407 675427 965463
rect 675483 965407 675507 965463
rect 675563 965407 675587 965463
rect 675643 965407 675667 965463
rect 675723 965407 675737 965463
rect 675407 965400 675737 965407
rect 41863 964397 42193 964404
rect 41863 964341 41883 964397
rect 41939 964341 41963 964397
rect 42019 964341 42043 964397
rect 42099 964341 42123 964397
rect 42179 964341 42193 964397
rect 41863 964334 42193 964341
rect 41863 963753 42193 963760
rect 41863 963697 41883 963753
rect 41939 963697 41963 963753
rect 42019 963697 42043 963753
rect 42099 963697 42123 963753
rect 42179 963697 42193 963753
rect 41863 963690 42193 963697
rect 675407 963623 675737 963630
rect 675407 963567 675427 963623
rect 675483 963567 675507 963623
rect 675563 963567 675587 963623
rect 675643 963567 675667 963623
rect 675723 963567 675737 963623
rect 675407 963560 675737 963567
rect 41863 963109 42193 963116
rect 41863 963053 41883 963109
rect 41939 963053 41963 963109
rect 42019 963053 42043 963109
rect 42099 963053 42123 963109
rect 42179 963053 42193 963109
rect 41863 963046 42193 963053
rect 675407 963071 675737 963078
rect 675407 963015 675427 963071
rect 675483 963015 675507 963071
rect 675563 963015 675587 963071
rect 675643 963015 675667 963071
rect 675723 963015 675737 963071
rect 675407 963008 675737 963015
rect 41863 962557 42193 962564
rect 41863 962501 41883 962557
rect 41939 962501 41963 962557
rect 42019 962501 42043 962557
rect 42099 962501 42123 962557
rect 42179 962501 42193 962557
rect 41863 962494 42193 962501
rect 675407 962427 675737 962434
rect 675407 962371 675427 962427
rect 675483 962371 675507 962427
rect 675563 962371 675587 962427
rect 675643 962371 675667 962427
rect 675723 962371 675737 962427
rect 675407 962364 675737 962371
rect 675407 961783 675737 961790
rect 675407 961727 675427 961783
rect 675483 961727 675507 961783
rect 675563 961727 675587 961783
rect 675643 961727 675667 961783
rect 675723 961727 675737 961783
rect 675407 961720 675737 961727
rect 41863 960073 42193 960080
rect 41863 960017 41883 960073
rect 41939 960017 41963 960073
rect 42019 960017 42043 960073
rect 42099 960017 42123 960073
rect 42179 960017 42193 960073
rect 41863 960010 42193 960017
rect 41863 959429 42193 959436
rect 41863 959373 41883 959429
rect 41939 959373 41963 959429
rect 42019 959373 42043 959429
rect 42099 959373 42123 959429
rect 42179 959373 42193 959429
rect 41863 959366 42193 959373
rect 675407 959299 675737 959306
rect 675407 959243 675427 959299
rect 675483 959243 675507 959299
rect 675563 959243 675587 959299
rect 675643 959243 675667 959299
rect 675723 959243 675737 959299
rect 675407 959236 675737 959243
rect 41863 958785 42193 958792
rect 41863 958729 41883 958785
rect 41939 958729 41963 958785
rect 42019 958729 42043 958785
rect 42099 958729 42123 958785
rect 42179 958729 42193 958785
rect 41863 958722 42193 958729
rect 675407 958747 675737 958754
rect 675407 958691 675427 958747
rect 675483 958691 675507 958747
rect 675563 958691 675587 958747
rect 675643 958691 675667 958747
rect 675723 958691 675737 958747
rect 675407 958684 675737 958691
rect 41863 958233 42193 958240
rect 41863 958177 41883 958233
rect 41939 958177 41963 958233
rect 42019 958177 42043 958233
rect 42099 958177 42123 958233
rect 42179 958177 42193 958233
rect 41863 958170 42193 958177
rect 675407 958103 675737 958110
rect 675407 958047 675427 958103
rect 675483 958047 675507 958103
rect 675563 958047 675587 958103
rect 675643 958047 675667 958103
rect 675723 958047 675737 958103
rect 675407 958040 675737 958047
rect 675407 957459 675737 957466
rect 675407 957403 675427 957459
rect 675483 957403 675507 957459
rect 675563 957403 675587 957459
rect 675643 957403 675667 957459
rect 675723 957403 675737 957459
rect 675407 957396 675737 957403
rect 41863 956393 42193 956400
rect 41863 956337 41883 956393
rect 41939 956337 41963 956393
rect 42019 956337 42043 956393
rect 42099 956337 42123 956393
rect 42179 956337 42193 956393
rect 41863 956330 42193 956337
rect 675407 956263 675737 956270
rect 675407 956207 675427 956263
rect 675483 956207 675507 956263
rect 675563 956207 675587 956263
rect 675643 956207 675667 956263
rect 675723 956207 675737 956263
rect 675407 956200 675737 956207
rect 41863 955749 42193 955756
rect 41863 955693 41883 955749
rect 41939 955693 41963 955749
rect 42019 955693 42043 955749
rect 42099 955693 42123 955749
rect 42179 955693 42193 955749
rect 41863 955686 42193 955693
rect 41863 955105 42193 955112
rect 41863 955049 41883 955105
rect 41939 955049 41963 955105
rect 42019 955049 42043 955105
rect 42099 955049 42123 955105
rect 42179 955049 42193 955105
rect 41863 955042 42193 955049
rect 675407 955067 675737 955074
rect 675407 955011 675427 955067
rect 675483 955011 675507 955067
rect 675563 955011 675587 955067
rect 675643 955011 675667 955067
rect 675723 955011 675737 955067
rect 675407 955004 675737 955011
rect 675407 954423 675737 954430
rect 675407 954367 675427 954423
rect 675483 954367 675507 954423
rect 675563 954367 675587 954423
rect 675643 954367 675667 954423
rect 675723 954367 675737 954423
rect 675407 954360 675737 954367
rect 675407 953779 675737 953786
rect 675407 953723 675427 953779
rect 675483 953723 675507 953779
rect 675563 953723 675587 953779
rect 675643 953723 675667 953779
rect 675723 953723 675737 953779
rect 675407 953716 675737 953723
rect 675407 952583 675737 952590
rect 675407 952527 675427 952583
rect 675483 952527 675507 952583
rect 675563 952527 675587 952583
rect 675643 952527 675667 952583
rect 675723 952527 675737 952583
rect 675407 952520 675737 952527
rect 675407 877551 675737 877558
rect 675407 877495 675427 877551
rect 675483 877495 675507 877551
rect 675563 877495 675587 877551
rect 675643 877495 675667 877551
rect 675723 877495 675737 877551
rect 675407 877488 675737 877495
rect 675407 876907 675737 876914
rect 675407 876851 675427 876907
rect 675483 876851 675507 876907
rect 675563 876851 675587 876907
rect 675643 876851 675667 876907
rect 675723 876851 675737 876907
rect 675407 876844 675737 876851
rect 675407 876263 675737 876270
rect 675407 876207 675427 876263
rect 675483 876207 675507 876263
rect 675563 876207 675587 876263
rect 675643 876207 675667 876263
rect 675723 876207 675737 876263
rect 675407 876200 675737 876207
rect 675407 874423 675737 874430
rect 675407 874367 675427 874423
rect 675483 874367 675507 874423
rect 675563 874367 675587 874423
rect 675643 874367 675667 874423
rect 675723 874367 675737 874423
rect 675407 874360 675737 874367
rect 675407 873871 675737 873878
rect 675407 873815 675427 873871
rect 675483 873815 675507 873871
rect 675563 873815 675587 873871
rect 675643 873815 675667 873871
rect 675723 873815 675737 873871
rect 675407 873808 675737 873815
rect 675407 873227 675737 873234
rect 675407 873171 675427 873227
rect 675483 873171 675507 873227
rect 675563 873171 675587 873227
rect 675643 873171 675667 873227
rect 675723 873171 675737 873227
rect 675407 873164 675737 873171
rect 675407 872583 675737 872590
rect 675407 872527 675427 872583
rect 675483 872527 675507 872583
rect 675563 872527 675587 872583
rect 675643 872527 675667 872583
rect 675723 872527 675737 872583
rect 675407 872520 675737 872527
rect 675407 870099 675737 870106
rect 675407 870043 675427 870099
rect 675483 870043 675507 870099
rect 675563 870043 675587 870099
rect 675643 870043 675667 870099
rect 675723 870043 675737 870099
rect 675407 870036 675737 870043
rect 675407 869547 675737 869554
rect 675407 869491 675427 869547
rect 675483 869491 675507 869547
rect 675563 869491 675587 869547
rect 675643 869491 675667 869547
rect 675723 869491 675737 869547
rect 675407 869484 675737 869491
rect 675407 868903 675737 868910
rect 675407 868847 675427 868903
rect 675483 868847 675507 868903
rect 675563 868847 675587 868903
rect 675643 868847 675667 868903
rect 675723 868847 675737 868903
rect 675407 868840 675737 868847
rect 675407 868259 675737 868266
rect 675407 868203 675427 868259
rect 675483 868203 675507 868259
rect 675563 868203 675587 868259
rect 675643 868203 675667 868259
rect 675723 868203 675737 868259
rect 675407 868196 675737 868203
rect 675407 867063 675737 867070
rect 675407 867007 675427 867063
rect 675483 867007 675507 867063
rect 675563 867007 675587 867063
rect 675643 867007 675667 867063
rect 675723 867007 675737 867063
rect 675407 867000 675737 867007
rect 675407 865867 675737 865874
rect 675407 865811 675427 865867
rect 675483 865811 675507 865867
rect 675563 865811 675587 865867
rect 675643 865811 675667 865867
rect 675723 865811 675737 865867
rect 675407 865804 675737 865811
rect 675407 865223 675737 865230
rect 675407 865167 675427 865223
rect 675483 865167 675507 865223
rect 675563 865167 675587 865223
rect 675643 865167 675667 865223
rect 675723 865167 675737 865223
rect 675407 865160 675737 865167
rect 675407 864579 675737 864586
rect 675407 864523 675427 864579
rect 675483 864523 675507 864579
rect 675563 864523 675587 864579
rect 675643 864523 675667 864579
rect 675723 864523 675737 864579
rect 675407 864516 675737 864523
rect 675407 863383 675737 863390
rect 675407 863327 675427 863383
rect 675483 863327 675507 863383
rect 675563 863327 675587 863383
rect 675643 863327 675667 863383
rect 675723 863327 675737 863383
rect 675407 863320 675737 863327
rect 41863 799473 42193 799480
rect 41863 799417 41883 799473
rect 41939 799417 41963 799473
rect 42019 799417 42043 799473
rect 42099 799417 42123 799473
rect 42179 799417 42193 799473
rect 41863 799410 42193 799417
rect 41863 798277 42193 798284
rect 41863 798221 41883 798277
rect 41939 798221 41963 798277
rect 42019 798221 42043 798277
rect 42099 798221 42123 798277
rect 42179 798221 42193 798277
rect 41863 798214 42193 798221
rect 41863 797633 42193 797640
rect 41863 797577 41883 797633
rect 41939 797577 41963 797633
rect 42019 797577 42043 797633
rect 42099 797577 42123 797633
rect 42179 797577 42193 797633
rect 41863 797570 42193 797577
rect 41863 796989 42193 796996
rect 41863 796933 41883 796989
rect 41939 796933 41963 796989
rect 42019 796933 42043 796989
rect 42099 796933 42123 796989
rect 42179 796933 42193 796989
rect 41863 796926 42193 796933
rect 41863 795793 42193 795800
rect 41863 795737 41883 795793
rect 41939 795737 41963 795793
rect 42019 795737 42043 795793
rect 42099 795737 42123 795793
rect 42179 795737 42193 795793
rect 41863 795730 42193 795737
rect 41863 794597 42193 794604
rect 41863 794541 41883 794597
rect 41939 794541 41963 794597
rect 42019 794541 42043 794597
rect 42099 794541 42123 794597
rect 42179 794541 42193 794597
rect 41863 794534 42193 794541
rect 41863 793953 42193 793960
rect 41863 793897 41883 793953
rect 41939 793897 41963 793953
rect 42019 793897 42043 793953
rect 42099 793897 42123 793953
rect 42179 793897 42193 793953
rect 41863 793890 42193 793897
rect 41863 793309 42193 793316
rect 41863 793253 41883 793309
rect 41939 793253 41963 793309
rect 42019 793253 42043 793309
rect 42099 793253 42123 793309
rect 42179 793253 42193 793309
rect 41863 793246 42193 793253
rect 41863 792757 42193 792764
rect 41863 792701 41883 792757
rect 41939 792701 41963 792757
rect 42019 792701 42043 792757
rect 42099 792701 42123 792757
rect 42179 792701 42193 792757
rect 41863 792694 42193 792701
rect 41863 790273 42193 790280
rect 41863 790217 41883 790273
rect 41939 790217 41963 790273
rect 42019 790217 42043 790273
rect 42099 790217 42123 790273
rect 42179 790217 42193 790273
rect 41863 790210 42193 790217
rect 41863 789629 42193 789636
rect 41863 789573 41883 789629
rect 41939 789573 41963 789629
rect 42019 789573 42043 789629
rect 42099 789573 42123 789629
rect 42179 789573 42193 789629
rect 41863 789566 42193 789573
rect 41863 788985 42193 788992
rect 41863 788929 41883 788985
rect 41939 788929 41963 788985
rect 42019 788929 42043 788985
rect 42099 788929 42123 788985
rect 42179 788929 42193 788985
rect 41863 788922 42193 788929
rect 41863 788433 42193 788440
rect 41863 788377 41883 788433
rect 41939 788377 41963 788433
rect 42019 788377 42043 788433
rect 42099 788377 42123 788433
rect 42179 788377 42193 788433
rect 41863 788370 42193 788377
rect 675407 788351 675737 788358
rect 675407 788295 675427 788351
rect 675483 788295 675507 788351
rect 675563 788295 675587 788351
rect 675643 788295 675667 788351
rect 675723 788295 675737 788351
rect 675407 788288 675737 788295
rect 675407 787707 675737 787714
rect 675407 787651 675427 787707
rect 675483 787651 675507 787707
rect 675563 787651 675587 787707
rect 675643 787651 675667 787707
rect 675723 787651 675737 787707
rect 675407 787644 675737 787651
rect 675407 787063 675737 787070
rect 675407 787007 675427 787063
rect 675483 787007 675507 787063
rect 675563 787007 675587 787063
rect 675643 787007 675667 787063
rect 675723 787007 675737 787063
rect 675407 787000 675737 787007
rect 41863 786593 42193 786600
rect 41863 786537 41883 786593
rect 41939 786537 41963 786593
rect 42019 786537 42043 786593
rect 42099 786537 42123 786593
rect 42179 786537 42193 786593
rect 41863 786530 42193 786537
rect 41863 785949 42193 785956
rect 41863 785893 41883 785949
rect 41939 785893 41963 785949
rect 42019 785893 42043 785949
rect 42099 785893 42123 785949
rect 42179 785893 42193 785949
rect 41863 785886 42193 785893
rect 41863 785305 42193 785312
rect 41863 785249 41883 785305
rect 41939 785249 41963 785305
rect 42019 785249 42043 785305
rect 42099 785249 42123 785305
rect 42179 785249 42193 785305
rect 41863 785242 42193 785249
rect 675407 785223 675737 785230
rect 675407 785167 675427 785223
rect 675483 785167 675507 785223
rect 675563 785167 675587 785223
rect 675643 785167 675667 785223
rect 675723 785167 675737 785223
rect 675407 785160 675737 785167
rect 675407 784671 675737 784678
rect 675407 784615 675427 784671
rect 675483 784615 675507 784671
rect 675563 784615 675587 784671
rect 675643 784615 675667 784671
rect 675723 784615 675737 784671
rect 675407 784608 675737 784615
rect 675407 784027 675737 784034
rect 675407 783971 675427 784027
rect 675483 783971 675507 784027
rect 675563 783971 675587 784027
rect 675643 783971 675667 784027
rect 675723 783971 675737 784027
rect 675407 783964 675737 783971
rect 675407 783383 675737 783390
rect 675407 783327 675427 783383
rect 675483 783327 675507 783383
rect 675563 783327 675587 783383
rect 675643 783327 675667 783383
rect 675723 783327 675737 783383
rect 675407 783320 675737 783327
rect 675407 780899 675737 780906
rect 675407 780843 675427 780899
rect 675483 780843 675507 780899
rect 675563 780843 675587 780899
rect 675643 780843 675667 780899
rect 675723 780843 675737 780899
rect 675407 780836 675737 780843
rect 675407 780347 675737 780354
rect 675407 780291 675427 780347
rect 675483 780291 675507 780347
rect 675563 780291 675587 780347
rect 675643 780291 675667 780347
rect 675723 780291 675737 780347
rect 675407 780284 675737 780291
rect 675407 779703 675737 779710
rect 675407 779647 675427 779703
rect 675483 779647 675507 779703
rect 675563 779647 675587 779703
rect 675643 779647 675667 779703
rect 675723 779647 675737 779703
rect 675407 779640 675737 779647
rect 675407 779059 675737 779066
rect 675407 779003 675427 779059
rect 675483 779003 675507 779059
rect 675563 779003 675587 779059
rect 675643 779003 675667 779059
rect 675723 779003 675737 779059
rect 675407 778996 675737 779003
rect 675407 777863 675737 777870
rect 675407 777807 675427 777863
rect 675483 777807 675507 777863
rect 675563 777807 675587 777863
rect 675643 777807 675667 777863
rect 675723 777807 675737 777863
rect 675407 777800 675737 777807
rect 675407 776667 675737 776674
rect 675407 776611 675427 776667
rect 675483 776611 675507 776667
rect 675563 776611 675587 776667
rect 675643 776611 675667 776667
rect 675723 776611 675737 776667
rect 675407 776604 675737 776611
rect 675407 776023 675737 776030
rect 675407 775967 675427 776023
rect 675483 775967 675507 776023
rect 675563 775967 675587 776023
rect 675643 775967 675667 776023
rect 675723 775967 675737 776023
rect 675407 775960 675737 775967
rect 675407 775379 675737 775386
rect 675407 775323 675427 775379
rect 675483 775323 675507 775379
rect 675563 775323 675587 775379
rect 675643 775323 675667 775379
rect 675723 775323 675737 775379
rect 675407 775316 675737 775323
rect 675407 774183 675737 774190
rect 675407 774127 675427 774183
rect 675483 774127 675507 774183
rect 675563 774127 675587 774183
rect 675643 774127 675667 774183
rect 675723 774127 675737 774183
rect 675407 774120 675737 774127
rect 41863 756273 42193 756280
rect 41863 756217 41883 756273
rect 41939 756217 41963 756273
rect 42019 756217 42043 756273
rect 42099 756217 42123 756273
rect 42179 756217 42193 756273
rect 41863 756210 42193 756217
rect 41863 755077 42193 755084
rect 41863 755021 41883 755077
rect 41939 755021 41963 755077
rect 42019 755021 42043 755077
rect 42099 755021 42123 755077
rect 42179 755021 42193 755077
rect 41863 755014 42193 755021
rect 41863 754433 42193 754440
rect 41863 754377 41883 754433
rect 41939 754377 41963 754433
rect 42019 754377 42043 754433
rect 42099 754377 42123 754433
rect 42179 754377 42193 754433
rect 41863 754370 42193 754377
rect 41863 753789 42193 753796
rect 41863 753733 41883 753789
rect 41939 753733 41963 753789
rect 42019 753733 42043 753789
rect 42099 753733 42123 753789
rect 42179 753733 42193 753789
rect 41863 753726 42193 753733
rect 41863 752593 42193 752600
rect 41863 752537 41883 752593
rect 41939 752537 41963 752593
rect 42019 752537 42043 752593
rect 42099 752537 42123 752593
rect 42179 752537 42193 752593
rect 41863 752530 42193 752537
rect 41863 751397 42193 751404
rect 41863 751341 41883 751397
rect 41939 751341 41963 751397
rect 42019 751341 42043 751397
rect 42099 751341 42123 751397
rect 42179 751341 42193 751397
rect 41863 751334 42193 751341
rect 41863 750753 42193 750760
rect 41863 750697 41883 750753
rect 41939 750697 41963 750753
rect 42019 750697 42043 750753
rect 42099 750697 42123 750753
rect 42179 750697 42193 750753
rect 41863 750690 42193 750697
rect 41863 750109 42193 750116
rect 41863 750053 41883 750109
rect 41939 750053 41963 750109
rect 42019 750053 42043 750109
rect 42099 750053 42123 750109
rect 42179 750053 42193 750109
rect 41863 750046 42193 750053
rect 41863 749557 42193 749564
rect 41863 749501 41883 749557
rect 41939 749501 41963 749557
rect 42019 749501 42043 749557
rect 42099 749501 42123 749557
rect 42179 749501 42193 749557
rect 41863 749494 42193 749501
rect 41863 747073 42193 747080
rect 41863 747017 41883 747073
rect 41939 747017 41963 747073
rect 42019 747017 42043 747073
rect 42099 747017 42123 747073
rect 42179 747017 42193 747073
rect 41863 747010 42193 747017
rect 41863 746429 42193 746436
rect 41863 746373 41883 746429
rect 41939 746373 41963 746429
rect 42019 746373 42043 746429
rect 42099 746373 42123 746429
rect 42179 746373 42193 746429
rect 41863 746366 42193 746373
rect 41863 745785 42193 745792
rect 41863 745729 41883 745785
rect 41939 745729 41963 745785
rect 42019 745729 42043 745785
rect 42099 745729 42123 745785
rect 42179 745729 42193 745785
rect 41863 745722 42193 745729
rect 41863 745233 42193 745240
rect 41863 745177 41883 745233
rect 41939 745177 41963 745233
rect 42019 745177 42043 745233
rect 42099 745177 42123 745233
rect 42179 745177 42193 745233
rect 41863 745170 42193 745177
rect 41863 743393 42193 743400
rect 41863 743337 41883 743393
rect 41939 743337 41963 743393
rect 42019 743337 42043 743393
rect 42099 743337 42123 743393
rect 42179 743337 42193 743393
rect 41863 743330 42193 743337
rect 675407 743351 675737 743358
rect 675407 743295 675427 743351
rect 675483 743295 675507 743351
rect 675563 743295 675587 743351
rect 675643 743295 675667 743351
rect 675723 743295 675737 743351
rect 675407 743288 675737 743295
rect 41863 742749 42193 742756
rect 41863 742693 41883 742749
rect 41939 742693 41963 742749
rect 42019 742693 42043 742749
rect 42099 742693 42123 742749
rect 42179 742693 42193 742749
rect 41863 742686 42193 742693
rect 675407 742707 675737 742714
rect 675407 742651 675427 742707
rect 675483 742651 675507 742707
rect 675563 742651 675587 742707
rect 675643 742651 675667 742707
rect 675723 742651 675737 742707
rect 675407 742644 675737 742651
rect 41863 742105 42193 742112
rect 41863 742049 41883 742105
rect 41939 742049 41963 742105
rect 42019 742049 42043 742105
rect 42099 742049 42123 742105
rect 42179 742049 42193 742105
rect 41863 742042 42193 742049
rect 675407 742063 675737 742070
rect 675407 742007 675427 742063
rect 675483 742007 675507 742063
rect 675563 742007 675587 742063
rect 675643 742007 675667 742063
rect 675723 742007 675737 742063
rect 675407 742000 675737 742007
rect 675407 740223 675737 740230
rect 675407 740167 675427 740223
rect 675483 740167 675507 740223
rect 675563 740167 675587 740223
rect 675643 740167 675667 740223
rect 675723 740167 675737 740223
rect 675407 740160 675737 740167
rect 675407 739671 675737 739678
rect 675407 739615 675427 739671
rect 675483 739615 675507 739671
rect 675563 739615 675587 739671
rect 675643 739615 675667 739671
rect 675723 739615 675737 739671
rect 675407 739608 675737 739615
rect 675407 739027 675737 739034
rect 675407 738971 675427 739027
rect 675483 738971 675507 739027
rect 675563 738971 675587 739027
rect 675643 738971 675667 739027
rect 675723 738971 675737 739027
rect 675407 738964 675737 738971
rect 675407 738383 675737 738390
rect 675407 738327 675427 738383
rect 675483 738327 675507 738383
rect 675563 738327 675587 738383
rect 675643 738327 675667 738383
rect 675723 738327 675737 738383
rect 675407 738320 675737 738327
rect 675407 735899 675737 735906
rect 675407 735843 675427 735899
rect 675483 735843 675507 735899
rect 675563 735843 675587 735899
rect 675643 735843 675667 735899
rect 675723 735843 675737 735899
rect 675407 735836 675737 735843
rect 675407 735347 675737 735354
rect 675407 735291 675427 735347
rect 675483 735291 675507 735347
rect 675563 735291 675587 735347
rect 675643 735291 675667 735347
rect 675723 735291 675737 735347
rect 675407 735284 675737 735291
rect 675407 734703 675737 734710
rect 675407 734647 675427 734703
rect 675483 734647 675507 734703
rect 675563 734647 675587 734703
rect 675643 734647 675667 734703
rect 675723 734647 675737 734703
rect 675407 734640 675737 734647
rect 675407 734059 675737 734066
rect 675407 734003 675427 734059
rect 675483 734003 675507 734059
rect 675563 734003 675587 734059
rect 675643 734003 675667 734059
rect 675723 734003 675737 734059
rect 675407 733996 675737 734003
rect 675407 732863 675737 732870
rect 675407 732807 675427 732863
rect 675483 732807 675507 732863
rect 675563 732807 675587 732863
rect 675643 732807 675667 732863
rect 675723 732807 675737 732863
rect 675407 732800 675737 732807
rect 675407 731667 675737 731674
rect 675407 731611 675427 731667
rect 675483 731611 675507 731667
rect 675563 731611 675587 731667
rect 675643 731611 675667 731667
rect 675723 731611 675737 731667
rect 675407 731604 675737 731611
rect 675407 731023 675737 731030
rect 675407 730967 675427 731023
rect 675483 730967 675507 731023
rect 675563 730967 675587 731023
rect 675643 730967 675667 731023
rect 675723 730967 675737 731023
rect 675407 730960 675737 730967
rect 675407 730379 675737 730386
rect 675407 730323 675427 730379
rect 675483 730323 675507 730379
rect 675563 730323 675587 730379
rect 675643 730323 675667 730379
rect 675723 730323 675737 730379
rect 675407 730316 675737 730323
rect 675407 729183 675737 729190
rect 675407 729127 675427 729183
rect 675483 729127 675507 729183
rect 675563 729127 675587 729183
rect 675643 729127 675667 729183
rect 675723 729127 675737 729183
rect 675407 729120 675737 729127
rect 41863 713073 42193 713080
rect 41863 713017 41883 713073
rect 41939 713017 41963 713073
rect 42019 713017 42043 713073
rect 42099 713017 42123 713073
rect 42179 713017 42193 713073
rect 41863 713010 42193 713017
rect 41863 711877 42193 711884
rect 41863 711821 41883 711877
rect 41939 711821 41963 711877
rect 42019 711821 42043 711877
rect 42099 711821 42123 711877
rect 42179 711821 42193 711877
rect 41863 711814 42193 711821
rect 41863 711233 42193 711240
rect 41863 711177 41883 711233
rect 41939 711177 41963 711233
rect 42019 711177 42043 711233
rect 42099 711177 42123 711233
rect 42179 711177 42193 711233
rect 41863 711170 42193 711177
rect 41863 710589 42193 710596
rect 41863 710533 41883 710589
rect 41939 710533 41963 710589
rect 42019 710533 42043 710589
rect 42099 710533 42123 710589
rect 42179 710533 42193 710589
rect 41863 710526 42193 710533
rect 41863 709393 42193 709400
rect 41863 709337 41883 709393
rect 41939 709337 41963 709393
rect 42019 709337 42043 709393
rect 42099 709337 42123 709393
rect 42179 709337 42193 709393
rect 41863 709330 42193 709337
rect 41863 708197 42193 708204
rect 41863 708141 41883 708197
rect 41939 708141 41963 708197
rect 42019 708141 42043 708197
rect 42099 708141 42123 708197
rect 42179 708141 42193 708197
rect 41863 708134 42193 708141
rect 41863 707553 42193 707560
rect 41863 707497 41883 707553
rect 41939 707497 41963 707553
rect 42019 707497 42043 707553
rect 42099 707497 42123 707553
rect 42179 707497 42193 707553
rect 41863 707490 42193 707497
rect 41863 706909 42193 706916
rect 41863 706853 41883 706909
rect 41939 706853 41963 706909
rect 42019 706853 42043 706909
rect 42099 706853 42123 706909
rect 42179 706853 42193 706909
rect 41863 706846 42193 706853
rect 41863 706357 42193 706364
rect 41863 706301 41883 706357
rect 41939 706301 41963 706357
rect 42019 706301 42043 706357
rect 42099 706301 42123 706357
rect 42179 706301 42193 706357
rect 41863 706294 42193 706301
rect 41863 703873 42193 703880
rect 41863 703817 41883 703873
rect 41939 703817 41963 703873
rect 42019 703817 42043 703873
rect 42099 703817 42123 703873
rect 42179 703817 42193 703873
rect 41863 703810 42193 703817
rect 41863 703229 42193 703236
rect 41863 703173 41883 703229
rect 41939 703173 41963 703229
rect 42019 703173 42043 703229
rect 42099 703173 42123 703229
rect 42179 703173 42193 703229
rect 41863 703166 42193 703173
rect 41863 702585 42193 702592
rect 41863 702529 41883 702585
rect 41939 702529 41963 702585
rect 42019 702529 42043 702585
rect 42099 702529 42123 702585
rect 42179 702529 42193 702585
rect 41863 702522 42193 702529
rect 41863 702033 42193 702040
rect 41863 701977 41883 702033
rect 41939 701977 41963 702033
rect 42019 701977 42043 702033
rect 42099 701977 42123 702033
rect 42179 701977 42193 702033
rect 41863 701970 42193 701977
rect 41863 700193 42193 700200
rect 41863 700137 41883 700193
rect 41939 700137 41963 700193
rect 42019 700137 42043 700193
rect 42099 700137 42123 700193
rect 42179 700137 42193 700193
rect 41863 700130 42193 700137
rect 41863 699549 42193 699556
rect 41863 699493 41883 699549
rect 41939 699493 41963 699549
rect 42019 699493 42043 699549
rect 42099 699493 42123 699549
rect 42179 699493 42193 699549
rect 41863 699486 42193 699493
rect 41863 698905 42193 698912
rect 41863 698849 41883 698905
rect 41939 698849 41963 698905
rect 42019 698849 42043 698905
rect 42099 698849 42123 698905
rect 42179 698849 42193 698905
rect 41863 698842 42193 698849
rect 675407 698351 675737 698358
rect 675407 698295 675427 698351
rect 675483 698295 675507 698351
rect 675563 698295 675587 698351
rect 675643 698295 675667 698351
rect 675723 698295 675737 698351
rect 675407 698288 675737 698295
rect 675407 697707 675737 697714
rect 675407 697651 675427 697707
rect 675483 697651 675507 697707
rect 675563 697651 675587 697707
rect 675643 697651 675667 697707
rect 675723 697651 675737 697707
rect 675407 697644 675737 697651
rect 675407 697063 675737 697070
rect 675407 697007 675427 697063
rect 675483 697007 675507 697063
rect 675563 697007 675587 697063
rect 675643 697007 675667 697063
rect 675723 697007 675737 697063
rect 675407 697000 675737 697007
rect 675407 695223 675737 695230
rect 675407 695167 675427 695223
rect 675483 695167 675507 695223
rect 675563 695167 675587 695223
rect 675643 695167 675667 695223
rect 675723 695167 675737 695223
rect 675407 695160 675737 695167
rect 675407 694671 675737 694678
rect 675407 694615 675427 694671
rect 675483 694615 675507 694671
rect 675563 694615 675587 694671
rect 675643 694615 675667 694671
rect 675723 694615 675737 694671
rect 675407 694608 675737 694615
rect 675407 694027 675737 694034
rect 675407 693971 675427 694027
rect 675483 693971 675507 694027
rect 675563 693971 675587 694027
rect 675643 693971 675667 694027
rect 675723 693971 675737 694027
rect 675407 693964 675737 693971
rect 675407 693383 675737 693390
rect 675407 693327 675427 693383
rect 675483 693327 675507 693383
rect 675563 693327 675587 693383
rect 675643 693327 675667 693383
rect 675723 693327 675737 693383
rect 675407 693320 675737 693327
rect 675407 690899 675737 690906
rect 675407 690843 675427 690899
rect 675483 690843 675507 690899
rect 675563 690843 675587 690899
rect 675643 690843 675667 690899
rect 675723 690843 675737 690899
rect 675407 690836 675737 690843
rect 675407 690347 675737 690354
rect 675407 690291 675427 690347
rect 675483 690291 675507 690347
rect 675563 690291 675587 690347
rect 675643 690291 675667 690347
rect 675723 690291 675737 690347
rect 675407 690284 675737 690291
rect 675407 689703 675737 689710
rect 675407 689647 675427 689703
rect 675483 689647 675507 689703
rect 675563 689647 675587 689703
rect 675643 689647 675667 689703
rect 675723 689647 675737 689703
rect 675407 689640 675737 689647
rect 675407 689059 675737 689066
rect 675407 689003 675427 689059
rect 675483 689003 675507 689059
rect 675563 689003 675587 689059
rect 675643 689003 675667 689059
rect 675723 689003 675737 689059
rect 675407 688996 675737 689003
rect 675407 687863 675737 687870
rect 675407 687807 675427 687863
rect 675483 687807 675507 687863
rect 675563 687807 675587 687863
rect 675643 687807 675667 687863
rect 675723 687807 675737 687863
rect 675407 687800 675737 687807
rect 675407 686667 675737 686674
rect 675407 686611 675427 686667
rect 675483 686611 675507 686667
rect 675563 686611 675587 686667
rect 675643 686611 675667 686667
rect 675723 686611 675737 686667
rect 675407 686604 675737 686611
rect 675407 686023 675737 686030
rect 675407 685967 675427 686023
rect 675483 685967 675507 686023
rect 675563 685967 675587 686023
rect 675643 685967 675667 686023
rect 675723 685967 675737 686023
rect 675407 685960 675737 685967
rect 675407 685379 675737 685386
rect 675407 685323 675427 685379
rect 675483 685323 675507 685379
rect 675563 685323 675587 685379
rect 675643 685323 675667 685379
rect 675723 685323 675737 685379
rect 675407 685316 675737 685323
rect 675407 684183 675737 684190
rect 675407 684127 675427 684183
rect 675483 684127 675507 684183
rect 675563 684127 675587 684183
rect 675643 684127 675667 684183
rect 675723 684127 675737 684183
rect 675407 684120 675737 684127
rect 41863 669873 42193 669880
rect 41863 669817 41883 669873
rect 41939 669817 41963 669873
rect 42019 669817 42043 669873
rect 42099 669817 42123 669873
rect 42179 669817 42193 669873
rect 41863 669810 42193 669817
rect 41863 668677 42193 668684
rect 41863 668621 41883 668677
rect 41939 668621 41963 668677
rect 42019 668621 42043 668677
rect 42099 668621 42123 668677
rect 42179 668621 42193 668677
rect 41863 668614 42193 668621
rect 41863 668033 42193 668040
rect 41863 667977 41883 668033
rect 41939 667977 41963 668033
rect 42019 667977 42043 668033
rect 42099 667977 42123 668033
rect 42179 667977 42193 668033
rect 41863 667970 42193 667977
rect 41863 667389 42193 667396
rect 41863 667333 41883 667389
rect 41939 667333 41963 667389
rect 42019 667333 42043 667389
rect 42099 667333 42123 667389
rect 42179 667333 42193 667389
rect 41863 667326 42193 667333
rect 41863 666193 42193 666200
rect 41863 666137 41883 666193
rect 41939 666137 41963 666193
rect 42019 666137 42043 666193
rect 42099 666137 42123 666193
rect 42179 666137 42193 666193
rect 41863 666130 42193 666137
rect 41863 664997 42193 665004
rect 41863 664941 41883 664997
rect 41939 664941 41963 664997
rect 42019 664941 42043 664997
rect 42099 664941 42123 664997
rect 42179 664941 42193 664997
rect 41863 664934 42193 664941
rect 41863 664353 42193 664360
rect 41863 664297 41883 664353
rect 41939 664297 41963 664353
rect 42019 664297 42043 664353
rect 42099 664297 42123 664353
rect 42179 664297 42193 664353
rect 41863 664290 42193 664297
rect 41863 663709 42193 663716
rect 41863 663653 41883 663709
rect 41939 663653 41963 663709
rect 42019 663653 42043 663709
rect 42099 663653 42123 663709
rect 42179 663653 42193 663709
rect 41863 663646 42193 663653
rect 41863 663157 42193 663164
rect 41863 663101 41883 663157
rect 41939 663101 41963 663157
rect 42019 663101 42043 663157
rect 42099 663101 42123 663157
rect 42179 663101 42193 663157
rect 41863 663094 42193 663101
rect 41863 660673 42193 660680
rect 41863 660617 41883 660673
rect 41939 660617 41963 660673
rect 42019 660617 42043 660673
rect 42099 660617 42123 660673
rect 42179 660617 42193 660673
rect 41863 660610 42193 660617
rect 41863 660029 42193 660036
rect 41863 659973 41883 660029
rect 41939 659973 41963 660029
rect 42019 659973 42043 660029
rect 42099 659973 42123 660029
rect 42179 659973 42193 660029
rect 41863 659966 42193 659973
rect 41863 659385 42193 659392
rect 41863 659329 41883 659385
rect 41939 659329 41963 659385
rect 42019 659329 42043 659385
rect 42099 659329 42123 659385
rect 42179 659329 42193 659385
rect 41863 659322 42193 659329
rect 41863 658833 42193 658840
rect 41863 658777 41883 658833
rect 41939 658777 41963 658833
rect 42019 658777 42043 658833
rect 42099 658777 42123 658833
rect 42179 658777 42193 658833
rect 41863 658770 42193 658777
rect 41863 656993 42193 657000
rect 41863 656937 41883 656993
rect 41939 656937 41963 656993
rect 42019 656937 42043 656993
rect 42099 656937 42123 656993
rect 42179 656937 42193 656993
rect 41863 656930 42193 656937
rect 41863 656349 42193 656356
rect 41863 656293 41883 656349
rect 41939 656293 41963 656349
rect 42019 656293 42043 656349
rect 42099 656293 42123 656349
rect 42179 656293 42193 656349
rect 41863 656286 42193 656293
rect 41863 655705 42193 655712
rect 41863 655649 41883 655705
rect 41939 655649 41963 655705
rect 42019 655649 42043 655705
rect 42099 655649 42123 655705
rect 42179 655649 42193 655705
rect 41863 655642 42193 655649
rect 675407 653151 675737 653158
rect 675407 653095 675427 653151
rect 675483 653095 675507 653151
rect 675563 653095 675587 653151
rect 675643 653095 675667 653151
rect 675723 653095 675737 653151
rect 675407 653088 675737 653095
rect 675407 652507 675737 652514
rect 675407 652451 675427 652507
rect 675483 652451 675507 652507
rect 675563 652451 675587 652507
rect 675643 652451 675667 652507
rect 675723 652451 675737 652507
rect 675407 652444 675737 652451
rect 675407 651863 675737 651870
rect 675407 651807 675427 651863
rect 675483 651807 675507 651863
rect 675563 651807 675587 651863
rect 675643 651807 675667 651863
rect 675723 651807 675737 651863
rect 675407 651800 675737 651807
rect 675407 650023 675737 650030
rect 675407 649967 675427 650023
rect 675483 649967 675507 650023
rect 675563 649967 675587 650023
rect 675643 649967 675667 650023
rect 675723 649967 675737 650023
rect 675407 649960 675737 649967
rect 675407 649471 675737 649478
rect 675407 649415 675427 649471
rect 675483 649415 675507 649471
rect 675563 649415 675587 649471
rect 675643 649415 675667 649471
rect 675723 649415 675737 649471
rect 675407 649408 675737 649415
rect 675407 648827 675737 648834
rect 675407 648771 675427 648827
rect 675483 648771 675507 648827
rect 675563 648771 675587 648827
rect 675643 648771 675667 648827
rect 675723 648771 675737 648827
rect 675407 648764 675737 648771
rect 675407 648183 675737 648190
rect 675407 648127 675427 648183
rect 675483 648127 675507 648183
rect 675563 648127 675587 648183
rect 675643 648127 675667 648183
rect 675723 648127 675737 648183
rect 675407 648120 675737 648127
rect 675407 645699 675737 645706
rect 675407 645643 675427 645699
rect 675483 645643 675507 645699
rect 675563 645643 675587 645699
rect 675643 645643 675667 645699
rect 675723 645643 675737 645699
rect 675407 645636 675737 645643
rect 675407 645147 675737 645154
rect 675407 645091 675427 645147
rect 675483 645091 675507 645147
rect 675563 645091 675587 645147
rect 675643 645091 675667 645147
rect 675723 645091 675737 645147
rect 675407 645084 675737 645091
rect 675407 644503 675737 644510
rect 675407 644447 675427 644503
rect 675483 644447 675507 644503
rect 675563 644447 675587 644503
rect 675643 644447 675667 644503
rect 675723 644447 675737 644503
rect 675407 644440 675737 644447
rect 675407 643859 675737 643866
rect 675407 643803 675427 643859
rect 675483 643803 675507 643859
rect 675563 643803 675587 643859
rect 675643 643803 675667 643859
rect 675723 643803 675737 643859
rect 675407 643796 675737 643803
rect 675407 642663 675737 642670
rect 675407 642607 675427 642663
rect 675483 642607 675507 642663
rect 675563 642607 675587 642663
rect 675643 642607 675667 642663
rect 675723 642607 675737 642663
rect 675407 642600 675737 642607
rect 675407 641467 675737 641474
rect 675407 641411 675427 641467
rect 675483 641411 675507 641467
rect 675563 641411 675587 641467
rect 675643 641411 675667 641467
rect 675723 641411 675737 641467
rect 675407 641404 675737 641411
rect 675407 640823 675737 640830
rect 675407 640767 675427 640823
rect 675483 640767 675507 640823
rect 675563 640767 675587 640823
rect 675643 640767 675667 640823
rect 675723 640767 675737 640823
rect 675407 640760 675737 640767
rect 675407 640179 675737 640186
rect 675407 640123 675427 640179
rect 675483 640123 675507 640179
rect 675563 640123 675587 640179
rect 675643 640123 675667 640179
rect 675723 640123 675737 640179
rect 675407 640116 675737 640123
rect 675407 638983 675737 638990
rect 675407 638927 675427 638983
rect 675483 638927 675507 638983
rect 675563 638927 675587 638983
rect 675643 638927 675667 638983
rect 675723 638927 675737 638983
rect 675407 638920 675737 638927
rect 41863 626673 42193 626680
rect 41863 626617 41883 626673
rect 41939 626617 41963 626673
rect 42019 626617 42043 626673
rect 42099 626617 42123 626673
rect 42179 626617 42193 626673
rect 41863 626610 42193 626617
rect 41863 625477 42193 625484
rect 41863 625421 41883 625477
rect 41939 625421 41963 625477
rect 42019 625421 42043 625477
rect 42099 625421 42123 625477
rect 42179 625421 42193 625477
rect 41863 625414 42193 625421
rect 41863 624833 42193 624840
rect 41863 624777 41883 624833
rect 41939 624777 41963 624833
rect 42019 624777 42043 624833
rect 42099 624777 42123 624833
rect 42179 624777 42193 624833
rect 41863 624770 42193 624777
rect 41863 624189 42193 624196
rect 41863 624133 41883 624189
rect 41939 624133 41963 624189
rect 42019 624133 42043 624189
rect 42099 624133 42123 624189
rect 42179 624133 42193 624189
rect 41863 624126 42193 624133
rect 41863 622993 42193 623000
rect 41863 622937 41883 622993
rect 41939 622937 41963 622993
rect 42019 622937 42043 622993
rect 42099 622937 42123 622993
rect 42179 622937 42193 622993
rect 41863 622930 42193 622937
rect 41863 621797 42193 621804
rect 41863 621741 41883 621797
rect 41939 621741 41963 621797
rect 42019 621741 42043 621797
rect 42099 621741 42123 621797
rect 42179 621741 42193 621797
rect 41863 621734 42193 621741
rect 41863 621153 42193 621160
rect 41863 621097 41883 621153
rect 41939 621097 41963 621153
rect 42019 621097 42043 621153
rect 42099 621097 42123 621153
rect 42179 621097 42193 621153
rect 41863 621090 42193 621097
rect 41863 620509 42193 620516
rect 41863 620453 41883 620509
rect 41939 620453 41963 620509
rect 42019 620453 42043 620509
rect 42099 620453 42123 620509
rect 42179 620453 42193 620509
rect 41863 620446 42193 620453
rect 41863 619957 42193 619964
rect 41863 619901 41883 619957
rect 41939 619901 41963 619957
rect 42019 619901 42043 619957
rect 42099 619901 42123 619957
rect 42179 619901 42193 619957
rect 41863 619894 42193 619901
rect 41863 617473 42193 617480
rect 41863 617417 41883 617473
rect 41939 617417 41963 617473
rect 42019 617417 42043 617473
rect 42099 617417 42123 617473
rect 42179 617417 42193 617473
rect 41863 617410 42193 617417
rect 41863 616829 42193 616836
rect 41863 616773 41883 616829
rect 41939 616773 41963 616829
rect 42019 616773 42043 616829
rect 42099 616773 42123 616829
rect 42179 616773 42193 616829
rect 41863 616766 42193 616773
rect 41863 616185 42193 616192
rect 41863 616129 41883 616185
rect 41939 616129 41963 616185
rect 42019 616129 42043 616185
rect 42099 616129 42123 616185
rect 42179 616129 42193 616185
rect 41863 616122 42193 616129
rect 41863 615633 42193 615640
rect 41863 615577 41883 615633
rect 41939 615577 41963 615633
rect 42019 615577 42043 615633
rect 42099 615577 42123 615633
rect 42179 615577 42193 615633
rect 41863 615570 42193 615577
rect 41863 613793 42193 613800
rect 41863 613737 41883 613793
rect 41939 613737 41963 613793
rect 42019 613737 42043 613793
rect 42099 613737 42123 613793
rect 42179 613737 42193 613793
rect 41863 613730 42193 613737
rect 41863 613149 42193 613156
rect 41863 613093 41883 613149
rect 41939 613093 41963 613149
rect 42019 613093 42043 613149
rect 42099 613093 42123 613149
rect 42179 613093 42193 613149
rect 41863 613086 42193 613093
rect 41863 612505 42193 612512
rect 41863 612449 41883 612505
rect 41939 612449 41963 612505
rect 42019 612449 42043 612505
rect 42099 612449 42123 612505
rect 42179 612449 42193 612505
rect 41863 612442 42193 612449
rect 675407 608151 675737 608158
rect 675407 608095 675427 608151
rect 675483 608095 675507 608151
rect 675563 608095 675587 608151
rect 675643 608095 675667 608151
rect 675723 608095 675737 608151
rect 675407 608088 675737 608095
rect 675407 607507 675737 607514
rect 675407 607451 675427 607507
rect 675483 607451 675507 607507
rect 675563 607451 675587 607507
rect 675643 607451 675667 607507
rect 675723 607451 675737 607507
rect 675407 607444 675737 607451
rect 675407 606863 675737 606870
rect 675407 606807 675427 606863
rect 675483 606807 675507 606863
rect 675563 606807 675587 606863
rect 675643 606807 675667 606863
rect 675723 606807 675737 606863
rect 675407 606800 675737 606807
rect 675407 605023 675737 605030
rect 675407 604967 675427 605023
rect 675483 604967 675507 605023
rect 675563 604967 675587 605023
rect 675643 604967 675667 605023
rect 675723 604967 675737 605023
rect 675407 604960 675737 604967
rect 675407 604471 675737 604478
rect 675407 604415 675427 604471
rect 675483 604415 675507 604471
rect 675563 604415 675587 604471
rect 675643 604415 675667 604471
rect 675723 604415 675737 604471
rect 675407 604408 675737 604415
rect 675407 603827 675737 603834
rect 675407 603771 675427 603827
rect 675483 603771 675507 603827
rect 675563 603771 675587 603827
rect 675643 603771 675667 603827
rect 675723 603771 675737 603827
rect 675407 603764 675737 603771
rect 675407 603183 675737 603190
rect 675407 603127 675427 603183
rect 675483 603127 675507 603183
rect 675563 603127 675587 603183
rect 675643 603127 675667 603183
rect 675723 603127 675737 603183
rect 675407 603120 675737 603127
rect 675407 600699 675737 600706
rect 675407 600643 675427 600699
rect 675483 600643 675507 600699
rect 675563 600643 675587 600699
rect 675643 600643 675667 600699
rect 675723 600643 675737 600699
rect 675407 600636 675737 600643
rect 675407 600147 675737 600154
rect 675407 600091 675427 600147
rect 675483 600091 675507 600147
rect 675563 600091 675587 600147
rect 675643 600091 675667 600147
rect 675723 600091 675737 600147
rect 675407 600084 675737 600091
rect 675407 599503 675737 599510
rect 675407 599447 675427 599503
rect 675483 599447 675507 599503
rect 675563 599447 675587 599503
rect 675643 599447 675667 599503
rect 675723 599447 675737 599503
rect 675407 599440 675737 599447
rect 675407 598859 675737 598866
rect 675407 598803 675427 598859
rect 675483 598803 675507 598859
rect 675563 598803 675587 598859
rect 675643 598803 675667 598859
rect 675723 598803 675737 598859
rect 675407 598796 675737 598803
rect 675407 597663 675737 597670
rect 675407 597607 675427 597663
rect 675483 597607 675507 597663
rect 675563 597607 675587 597663
rect 675643 597607 675667 597663
rect 675723 597607 675737 597663
rect 675407 597600 675737 597607
rect 675407 596467 675737 596474
rect 675407 596411 675427 596467
rect 675483 596411 675507 596467
rect 675563 596411 675587 596467
rect 675643 596411 675667 596467
rect 675723 596411 675737 596467
rect 675407 596404 675737 596411
rect 675407 595823 675737 595830
rect 675407 595767 675427 595823
rect 675483 595767 675507 595823
rect 675563 595767 675587 595823
rect 675643 595767 675667 595823
rect 675723 595767 675737 595823
rect 675407 595760 675737 595767
rect 675407 595179 675737 595186
rect 675407 595123 675427 595179
rect 675483 595123 675507 595179
rect 675563 595123 675587 595179
rect 675643 595123 675667 595179
rect 675723 595123 675737 595179
rect 675407 595116 675737 595123
rect 675407 593983 675737 593990
rect 675407 593927 675427 593983
rect 675483 593927 675507 593983
rect 675563 593927 675587 593983
rect 675643 593927 675667 593983
rect 675723 593927 675737 593983
rect 675407 593920 675737 593927
rect 41863 583473 42193 583480
rect 41863 583417 41883 583473
rect 41939 583417 41963 583473
rect 42019 583417 42043 583473
rect 42099 583417 42123 583473
rect 42179 583417 42193 583473
rect 41863 583410 42193 583417
rect 41863 582277 42193 582284
rect 41863 582221 41883 582277
rect 41939 582221 41963 582277
rect 42019 582221 42043 582277
rect 42099 582221 42123 582277
rect 42179 582221 42193 582277
rect 41863 582214 42193 582221
rect 41863 581633 42193 581640
rect 41863 581577 41883 581633
rect 41939 581577 41963 581633
rect 42019 581577 42043 581633
rect 42099 581577 42123 581633
rect 42179 581577 42193 581633
rect 41863 581570 42193 581577
rect 41863 580989 42193 580996
rect 41863 580933 41883 580989
rect 41939 580933 41963 580989
rect 42019 580933 42043 580989
rect 42099 580933 42123 580989
rect 42179 580933 42193 580989
rect 41863 580926 42193 580933
rect 41863 579793 42193 579800
rect 41863 579737 41883 579793
rect 41939 579737 41963 579793
rect 42019 579737 42043 579793
rect 42099 579737 42123 579793
rect 42179 579737 42193 579793
rect 41863 579730 42193 579737
rect 41863 578597 42193 578604
rect 41863 578541 41883 578597
rect 41939 578541 41963 578597
rect 42019 578541 42043 578597
rect 42099 578541 42123 578597
rect 42179 578541 42193 578597
rect 41863 578534 42193 578541
rect 41863 577953 42193 577960
rect 41863 577897 41883 577953
rect 41939 577897 41963 577953
rect 42019 577897 42043 577953
rect 42099 577897 42123 577953
rect 42179 577897 42193 577953
rect 41863 577890 42193 577897
rect 41863 577309 42193 577316
rect 41863 577253 41883 577309
rect 41939 577253 41963 577309
rect 42019 577253 42043 577309
rect 42099 577253 42123 577309
rect 42179 577253 42193 577309
rect 41863 577246 42193 577253
rect 41863 576757 42193 576764
rect 41863 576701 41883 576757
rect 41939 576701 41963 576757
rect 42019 576701 42043 576757
rect 42099 576701 42123 576757
rect 42179 576701 42193 576757
rect 41863 576694 42193 576701
rect 41863 574273 42193 574280
rect 41863 574217 41883 574273
rect 41939 574217 41963 574273
rect 42019 574217 42043 574273
rect 42099 574217 42123 574273
rect 42179 574217 42193 574273
rect 41863 574210 42193 574217
rect 41863 573629 42193 573636
rect 41863 573573 41883 573629
rect 41939 573573 41963 573629
rect 42019 573573 42043 573629
rect 42099 573573 42123 573629
rect 42179 573573 42193 573629
rect 41863 573566 42193 573573
rect 41863 572985 42193 572992
rect 41863 572929 41883 572985
rect 41939 572929 41963 572985
rect 42019 572929 42043 572985
rect 42099 572929 42123 572985
rect 42179 572929 42193 572985
rect 41863 572922 42193 572929
rect 41863 572433 42193 572440
rect 41863 572377 41883 572433
rect 41939 572377 41963 572433
rect 42019 572377 42043 572433
rect 42099 572377 42123 572433
rect 42179 572377 42193 572433
rect 41863 572370 42193 572377
rect 41863 570593 42193 570600
rect 41863 570537 41883 570593
rect 41939 570537 41963 570593
rect 42019 570537 42043 570593
rect 42099 570537 42123 570593
rect 42179 570537 42193 570593
rect 41863 570530 42193 570537
rect 41863 569949 42193 569956
rect 41863 569893 41883 569949
rect 41939 569893 41963 569949
rect 42019 569893 42043 569949
rect 42099 569893 42123 569949
rect 42179 569893 42193 569949
rect 41863 569886 42193 569893
rect 41863 569305 42193 569312
rect 41863 569249 41883 569305
rect 41939 569249 41963 569305
rect 42019 569249 42043 569305
rect 42099 569249 42123 569305
rect 42179 569249 42193 569305
rect 41863 569242 42193 569249
rect 675407 562951 675737 562958
rect 675407 562895 675427 562951
rect 675483 562895 675507 562951
rect 675563 562895 675587 562951
rect 675643 562895 675667 562951
rect 675723 562895 675737 562951
rect 675407 562888 675737 562895
rect 675407 562307 675737 562314
rect 675407 562251 675427 562307
rect 675483 562251 675507 562307
rect 675563 562251 675587 562307
rect 675643 562251 675667 562307
rect 675723 562251 675737 562307
rect 675407 562244 675737 562251
rect 675407 561663 675737 561670
rect 675407 561607 675427 561663
rect 675483 561607 675507 561663
rect 675563 561607 675587 561663
rect 675643 561607 675667 561663
rect 675723 561607 675737 561663
rect 675407 561600 675737 561607
rect 675407 559823 675737 559830
rect 675407 559767 675427 559823
rect 675483 559767 675507 559823
rect 675563 559767 675587 559823
rect 675643 559767 675667 559823
rect 675723 559767 675737 559823
rect 675407 559760 675737 559767
rect 675407 559271 675737 559278
rect 675407 559215 675427 559271
rect 675483 559215 675507 559271
rect 675563 559215 675587 559271
rect 675643 559215 675667 559271
rect 675723 559215 675737 559271
rect 675407 559208 675737 559215
rect 675407 558627 675737 558634
rect 675407 558571 675427 558627
rect 675483 558571 675507 558627
rect 675563 558571 675587 558627
rect 675643 558571 675667 558627
rect 675723 558571 675737 558627
rect 675407 558564 675737 558571
rect 675407 557983 675737 557990
rect 675407 557927 675427 557983
rect 675483 557927 675507 557983
rect 675563 557927 675587 557983
rect 675643 557927 675667 557983
rect 675723 557927 675737 557983
rect 675407 557920 675737 557927
rect 675407 555499 675737 555506
rect 675407 555443 675427 555499
rect 675483 555443 675507 555499
rect 675563 555443 675587 555499
rect 675643 555443 675667 555499
rect 675723 555443 675737 555499
rect 675407 555436 675737 555443
rect 675407 554947 675737 554954
rect 675407 554891 675427 554947
rect 675483 554891 675507 554947
rect 675563 554891 675587 554947
rect 675643 554891 675667 554947
rect 675723 554891 675737 554947
rect 675407 554884 675737 554891
rect 675407 554303 675737 554310
rect 675407 554247 675427 554303
rect 675483 554247 675507 554303
rect 675563 554247 675587 554303
rect 675643 554247 675667 554303
rect 675723 554247 675737 554303
rect 675407 554240 675737 554247
rect 675407 553659 675737 553666
rect 675407 553603 675427 553659
rect 675483 553603 675507 553659
rect 675563 553603 675587 553659
rect 675643 553603 675667 553659
rect 675723 553603 675737 553659
rect 675407 553596 675737 553603
rect 675407 552463 675737 552470
rect 675407 552407 675427 552463
rect 675483 552407 675507 552463
rect 675563 552407 675587 552463
rect 675643 552407 675667 552463
rect 675723 552407 675737 552463
rect 675407 552400 675737 552407
rect 675407 551267 675737 551274
rect 675407 551211 675427 551267
rect 675483 551211 675507 551267
rect 675563 551211 675587 551267
rect 675643 551211 675667 551267
rect 675723 551211 675737 551267
rect 675407 551204 675737 551211
rect 675407 550623 675737 550630
rect 675407 550567 675427 550623
rect 675483 550567 675507 550623
rect 675563 550567 675587 550623
rect 675643 550567 675667 550623
rect 675723 550567 675737 550623
rect 675407 550560 675737 550567
rect 675407 549979 675737 549986
rect 675407 549923 675427 549979
rect 675483 549923 675507 549979
rect 675563 549923 675587 549979
rect 675643 549923 675667 549979
rect 675723 549923 675737 549979
rect 675407 549916 675737 549923
rect 675407 548783 675737 548790
rect 675407 548727 675427 548783
rect 675483 548727 675507 548783
rect 675563 548727 675587 548783
rect 675643 548727 675667 548783
rect 675723 548727 675737 548783
rect 675407 548720 675737 548727
rect 41863 540273 42193 540280
rect 41863 540217 41883 540273
rect 41939 540217 41963 540273
rect 42019 540217 42043 540273
rect 42099 540217 42123 540273
rect 42179 540217 42193 540273
rect 41863 540210 42193 540217
rect 41863 539077 42193 539084
rect 41863 539021 41883 539077
rect 41939 539021 41963 539077
rect 42019 539021 42043 539077
rect 42099 539021 42123 539077
rect 42179 539021 42193 539077
rect 41863 539014 42193 539021
rect 41863 538433 42193 538440
rect 41863 538377 41883 538433
rect 41939 538377 41963 538433
rect 42019 538377 42043 538433
rect 42099 538377 42123 538433
rect 42179 538377 42193 538433
rect 41863 538370 42193 538377
rect 41863 537789 42193 537796
rect 41863 537733 41883 537789
rect 41939 537733 41963 537789
rect 42019 537733 42043 537789
rect 42099 537733 42123 537789
rect 42179 537733 42193 537789
rect 41863 537726 42193 537733
rect 41863 536593 42193 536600
rect 41863 536537 41883 536593
rect 41939 536537 41963 536593
rect 42019 536537 42043 536593
rect 42099 536537 42123 536593
rect 42179 536537 42193 536593
rect 41863 536530 42193 536537
rect 41863 535397 42193 535404
rect 41863 535341 41883 535397
rect 41939 535341 41963 535397
rect 42019 535341 42043 535397
rect 42099 535341 42123 535397
rect 42179 535341 42193 535397
rect 41863 535334 42193 535341
rect 41863 534753 42193 534760
rect 41863 534697 41883 534753
rect 41939 534697 41963 534753
rect 42019 534697 42043 534753
rect 42099 534697 42123 534753
rect 42179 534697 42193 534753
rect 41863 534690 42193 534697
rect 41863 534109 42193 534116
rect 41863 534053 41883 534109
rect 41939 534053 41963 534109
rect 42019 534053 42043 534109
rect 42099 534053 42123 534109
rect 42179 534053 42193 534109
rect 41863 534046 42193 534053
rect 41863 533557 42193 533564
rect 41863 533501 41883 533557
rect 41939 533501 41963 533557
rect 42019 533501 42043 533557
rect 42099 533501 42123 533557
rect 42179 533501 42193 533557
rect 41863 533494 42193 533501
rect 41863 531073 42193 531080
rect 41863 531017 41883 531073
rect 41939 531017 41963 531073
rect 42019 531017 42043 531073
rect 42099 531017 42123 531073
rect 42179 531017 42193 531073
rect 41863 531010 42193 531017
rect 41863 530429 42193 530436
rect 41863 530373 41883 530429
rect 41939 530373 41963 530429
rect 42019 530373 42043 530429
rect 42099 530373 42123 530429
rect 42179 530373 42193 530429
rect 41863 530366 42193 530373
rect 41863 529785 42193 529792
rect 41863 529729 41883 529785
rect 41939 529729 41963 529785
rect 42019 529729 42043 529785
rect 42099 529729 42123 529785
rect 42179 529729 42193 529785
rect 41863 529722 42193 529729
rect 41863 529233 42193 529240
rect 41863 529177 41883 529233
rect 41939 529177 41963 529233
rect 42019 529177 42043 529233
rect 42099 529177 42123 529233
rect 42179 529177 42193 529233
rect 41863 529170 42193 529177
rect 41863 527393 42193 527400
rect 41863 527337 41883 527393
rect 41939 527337 41963 527393
rect 42019 527337 42043 527393
rect 42099 527337 42123 527393
rect 42179 527337 42193 527393
rect 41863 527330 42193 527337
rect 41863 526749 42193 526756
rect 41863 526693 41883 526749
rect 41939 526693 41963 526749
rect 42019 526693 42043 526749
rect 42099 526693 42123 526749
rect 42179 526693 42193 526749
rect 41863 526686 42193 526693
rect 41863 526105 42193 526112
rect 41863 526049 41883 526105
rect 41939 526049 41963 526105
rect 42019 526049 42043 526105
rect 42099 526049 42123 526105
rect 42179 526049 42193 526105
rect 41863 526042 42193 526049
rect 41863 412673 42193 412680
rect 41863 412617 41883 412673
rect 41939 412617 41963 412673
rect 42019 412617 42043 412673
rect 42099 412617 42123 412673
rect 42179 412617 42193 412673
rect 41863 412610 42193 412617
rect 41863 411477 42193 411484
rect 41863 411421 41883 411477
rect 41939 411421 41963 411477
rect 42019 411421 42043 411477
rect 42099 411421 42123 411477
rect 42179 411421 42193 411477
rect 41863 411414 42193 411421
rect 41863 410833 42193 410840
rect 41863 410777 41883 410833
rect 41939 410777 41963 410833
rect 42019 410777 42043 410833
rect 42099 410777 42123 410833
rect 42179 410777 42193 410833
rect 41863 410770 42193 410777
rect 41863 410189 42193 410196
rect 41863 410133 41883 410189
rect 41939 410133 41963 410189
rect 42019 410133 42043 410189
rect 42099 410133 42123 410189
rect 42179 410133 42193 410189
rect 41863 410126 42193 410133
rect 41863 408993 42193 409000
rect 41863 408937 41883 408993
rect 41939 408937 41963 408993
rect 42019 408937 42043 408993
rect 42099 408937 42123 408993
rect 42179 408937 42193 408993
rect 41863 408930 42193 408937
rect 41863 407797 42193 407804
rect 41863 407741 41883 407797
rect 41939 407741 41963 407797
rect 42019 407741 42043 407797
rect 42099 407741 42123 407797
rect 42179 407741 42193 407797
rect 41863 407734 42193 407741
rect 41863 407153 42193 407160
rect 41863 407097 41883 407153
rect 41939 407097 41963 407153
rect 42019 407097 42043 407153
rect 42099 407097 42123 407153
rect 42179 407097 42193 407153
rect 41863 407090 42193 407097
rect 41863 406509 42193 406516
rect 41863 406453 41883 406509
rect 41939 406453 41963 406509
rect 42019 406453 42043 406509
rect 42099 406453 42123 406509
rect 42179 406453 42193 406509
rect 41863 406446 42193 406453
rect 41863 405957 42193 405964
rect 41863 405901 41883 405957
rect 41939 405901 41963 405957
rect 42019 405901 42043 405957
rect 42099 405901 42123 405957
rect 42179 405901 42193 405957
rect 41863 405894 42193 405901
rect 41863 403473 42193 403480
rect 41863 403417 41883 403473
rect 41939 403417 41963 403473
rect 42019 403417 42043 403473
rect 42099 403417 42123 403473
rect 42179 403417 42193 403473
rect 41863 403410 42193 403417
rect 41863 402829 42193 402836
rect 41863 402773 41883 402829
rect 41939 402773 41963 402829
rect 42019 402773 42043 402829
rect 42099 402773 42123 402829
rect 42179 402773 42193 402829
rect 41863 402766 42193 402773
rect 41863 402185 42193 402192
rect 41863 402129 41883 402185
rect 41939 402129 41963 402185
rect 42019 402129 42043 402185
rect 42099 402129 42123 402185
rect 42179 402129 42193 402185
rect 41863 402122 42193 402129
rect 41863 401633 42193 401640
rect 41863 401577 41883 401633
rect 41939 401577 41963 401633
rect 42019 401577 42043 401633
rect 42099 401577 42123 401633
rect 42179 401577 42193 401633
rect 41863 401570 42193 401577
rect 41863 399793 42193 399800
rect 41863 399737 41883 399793
rect 41939 399737 41963 399793
rect 42019 399737 42043 399793
rect 42099 399737 42123 399793
rect 42179 399737 42193 399793
rect 41863 399730 42193 399737
rect 41863 399149 42193 399156
rect 41863 399093 41883 399149
rect 41939 399093 41963 399149
rect 42019 399093 42043 399149
rect 42099 399093 42123 399149
rect 42179 399093 42193 399149
rect 41863 399086 42193 399093
rect 41863 398505 42193 398512
rect 41863 398449 41883 398505
rect 41939 398449 41963 398505
rect 42019 398449 42043 398505
rect 42099 398449 42123 398505
rect 42179 398449 42193 398505
rect 41863 398442 42193 398449
rect 675407 385751 675737 385758
rect 675407 385695 675427 385751
rect 675483 385695 675507 385751
rect 675563 385695 675587 385751
rect 675643 385695 675667 385751
rect 675723 385695 675737 385751
rect 675407 385688 675737 385695
rect 675407 385107 675737 385114
rect 675407 385051 675427 385107
rect 675483 385051 675507 385107
rect 675563 385051 675587 385107
rect 675643 385051 675667 385107
rect 675723 385051 675737 385107
rect 675407 385044 675737 385051
rect 675407 384463 675737 384470
rect 675407 384407 675427 384463
rect 675483 384407 675507 384463
rect 675563 384407 675587 384463
rect 675643 384407 675667 384463
rect 675723 384407 675737 384463
rect 675407 384400 675737 384407
rect 675407 382623 675737 382630
rect 675407 382567 675427 382623
rect 675483 382567 675507 382623
rect 675563 382567 675587 382623
rect 675643 382567 675667 382623
rect 675723 382567 675737 382623
rect 675407 382560 675737 382567
rect 675407 382071 675737 382078
rect 675407 382015 675427 382071
rect 675483 382015 675507 382071
rect 675563 382015 675587 382071
rect 675643 382015 675667 382071
rect 675723 382015 675737 382071
rect 675407 382008 675737 382015
rect 675407 381427 675737 381434
rect 675407 381371 675427 381427
rect 675483 381371 675507 381427
rect 675563 381371 675587 381427
rect 675643 381371 675667 381427
rect 675723 381371 675737 381427
rect 675407 381364 675737 381371
rect 675407 380783 675737 380790
rect 675407 380727 675427 380783
rect 675483 380727 675507 380783
rect 675563 380727 675587 380783
rect 675643 380727 675667 380783
rect 675723 380727 675737 380783
rect 675407 380720 675737 380727
rect 675407 378299 675737 378306
rect 675407 378243 675427 378299
rect 675483 378243 675507 378299
rect 675563 378243 675587 378299
rect 675643 378243 675667 378299
rect 675723 378243 675737 378299
rect 675407 378236 675737 378243
rect 675407 377747 675737 377754
rect 675407 377691 675427 377747
rect 675483 377691 675507 377747
rect 675563 377691 675587 377747
rect 675643 377691 675667 377747
rect 675723 377691 675737 377747
rect 675407 377684 675737 377691
rect 675407 377103 675737 377110
rect 675407 377047 675427 377103
rect 675483 377047 675507 377103
rect 675563 377047 675587 377103
rect 675643 377047 675667 377103
rect 675723 377047 675737 377103
rect 675407 377040 675737 377047
rect 675407 376459 675737 376466
rect 675407 376403 675427 376459
rect 675483 376403 675507 376459
rect 675563 376403 675587 376459
rect 675643 376403 675667 376459
rect 675723 376403 675737 376459
rect 675407 376396 675737 376403
rect 675407 375263 675737 375270
rect 675407 375207 675427 375263
rect 675483 375207 675507 375263
rect 675563 375207 675587 375263
rect 675643 375207 675667 375263
rect 675723 375207 675737 375263
rect 675407 375200 675737 375207
rect 675407 373423 675737 373430
rect 675407 373367 675427 373423
rect 675483 373367 675507 373423
rect 675563 373367 675587 373423
rect 675643 373367 675667 373423
rect 675723 373367 675737 373423
rect 675407 373360 675737 373367
rect 675407 372779 675737 372786
rect 675407 372723 675427 372779
rect 675483 372723 675507 372779
rect 675563 372723 675587 372779
rect 675643 372723 675667 372779
rect 675723 372723 675737 372779
rect 675407 372716 675737 372723
rect 675407 371583 675737 371590
rect 675407 371527 675427 371583
rect 675483 371527 675507 371583
rect 675563 371527 675587 371583
rect 675643 371527 675667 371583
rect 675723 371527 675737 371583
rect 675407 371520 675737 371527
rect 41863 369473 42193 369480
rect 41863 369417 41883 369473
rect 41939 369417 41963 369473
rect 42019 369417 42043 369473
rect 42099 369417 42123 369473
rect 42179 369417 42193 369473
rect 41863 369410 42193 369417
rect 41863 368277 42193 368284
rect 41863 368221 41883 368277
rect 41939 368221 41963 368277
rect 42019 368221 42043 368277
rect 42099 368221 42123 368277
rect 42179 368221 42193 368277
rect 41863 368214 42193 368221
rect 41863 367633 42193 367640
rect 41863 367577 41883 367633
rect 41939 367577 41963 367633
rect 42019 367577 42043 367633
rect 42099 367577 42123 367633
rect 42179 367577 42193 367633
rect 41863 367570 42193 367577
rect 41863 366989 42193 366996
rect 41863 366933 41883 366989
rect 41939 366933 41963 366989
rect 42019 366933 42043 366989
rect 42099 366933 42123 366989
rect 42179 366933 42193 366989
rect 41863 366926 42193 366933
rect 41863 365793 42193 365800
rect 41863 365737 41883 365793
rect 41939 365737 41963 365793
rect 42019 365737 42043 365793
rect 42099 365737 42123 365793
rect 42179 365737 42193 365793
rect 41863 365730 42193 365737
rect 41863 364597 42193 364604
rect 41863 364541 41883 364597
rect 41939 364541 41963 364597
rect 42019 364541 42043 364597
rect 42099 364541 42123 364597
rect 42179 364541 42193 364597
rect 41863 364534 42193 364541
rect 41863 363953 42193 363960
rect 41863 363897 41883 363953
rect 41939 363897 41963 363953
rect 42019 363897 42043 363953
rect 42099 363897 42123 363953
rect 42179 363897 42193 363953
rect 41863 363890 42193 363897
rect 41863 363309 42193 363316
rect 41863 363253 41883 363309
rect 41939 363253 41963 363309
rect 42019 363253 42043 363309
rect 42099 363253 42123 363309
rect 42179 363253 42193 363309
rect 41863 363246 42193 363253
rect 41863 362757 42193 362764
rect 41863 362701 41883 362757
rect 41939 362701 41963 362757
rect 42019 362701 42043 362757
rect 42099 362701 42123 362757
rect 42179 362701 42193 362757
rect 41863 362694 42193 362701
rect 41863 360273 42193 360280
rect 41863 360217 41883 360273
rect 41939 360217 41963 360273
rect 42019 360217 42043 360273
rect 42099 360217 42123 360273
rect 42179 360217 42193 360273
rect 41863 360210 42193 360217
rect 41863 359629 42193 359636
rect 41863 359573 41883 359629
rect 41939 359573 41963 359629
rect 42019 359573 42043 359629
rect 42099 359573 42123 359629
rect 42179 359573 42193 359629
rect 41863 359566 42193 359573
rect 41863 358985 42193 358992
rect 41863 358929 41883 358985
rect 41939 358929 41963 358985
rect 42019 358929 42043 358985
rect 42099 358929 42123 358985
rect 42179 358929 42193 358985
rect 41863 358922 42193 358929
rect 41863 358433 42193 358440
rect 41863 358377 41883 358433
rect 41939 358377 41963 358433
rect 42019 358377 42043 358433
rect 42099 358377 42123 358433
rect 42179 358377 42193 358433
rect 41863 358370 42193 358377
rect 41863 356593 42193 356600
rect 41863 356537 41883 356593
rect 41939 356537 41963 356593
rect 42019 356537 42043 356593
rect 42099 356537 42123 356593
rect 42179 356537 42193 356593
rect 41863 356530 42193 356537
rect 41863 355949 42193 355956
rect 41863 355893 41883 355949
rect 41939 355893 41963 355949
rect 42019 355893 42043 355949
rect 42099 355893 42123 355949
rect 42179 355893 42193 355949
rect 41863 355886 42193 355893
rect 41863 355305 42193 355312
rect 41863 355249 41883 355305
rect 41939 355249 41963 355305
rect 42019 355249 42043 355305
rect 42099 355249 42123 355305
rect 42179 355249 42193 355305
rect 41863 355242 42193 355249
rect 675407 340551 675737 340558
rect 675407 340495 675427 340551
rect 675483 340495 675507 340551
rect 675563 340495 675587 340551
rect 675643 340495 675667 340551
rect 675723 340495 675737 340551
rect 675407 340488 675737 340495
rect 675407 339907 675737 339914
rect 675407 339851 675427 339907
rect 675483 339851 675507 339907
rect 675563 339851 675587 339907
rect 675643 339851 675667 339907
rect 675723 339851 675737 339907
rect 675407 339844 675737 339851
rect 675407 339263 675737 339270
rect 675407 339207 675427 339263
rect 675483 339207 675507 339263
rect 675563 339207 675587 339263
rect 675643 339207 675667 339263
rect 675723 339207 675737 339263
rect 675407 339200 675737 339207
rect 675407 337423 675737 337430
rect 675407 337367 675427 337423
rect 675483 337367 675507 337423
rect 675563 337367 675587 337423
rect 675643 337367 675667 337423
rect 675723 337367 675737 337423
rect 675407 337360 675737 337367
rect 675407 336871 675737 336878
rect 675407 336815 675427 336871
rect 675483 336815 675507 336871
rect 675563 336815 675587 336871
rect 675643 336815 675667 336871
rect 675723 336815 675737 336871
rect 675407 336808 675737 336815
rect 675407 336227 675737 336234
rect 675407 336171 675427 336227
rect 675483 336171 675507 336227
rect 675563 336171 675587 336227
rect 675643 336171 675667 336227
rect 675723 336171 675737 336227
rect 675407 336164 675737 336171
rect 675407 335583 675737 335590
rect 675407 335527 675427 335583
rect 675483 335527 675507 335583
rect 675563 335527 675587 335583
rect 675643 335527 675667 335583
rect 675723 335527 675737 335583
rect 675407 335520 675737 335527
rect 675407 333099 675737 333106
rect 675407 333043 675427 333099
rect 675483 333043 675507 333099
rect 675563 333043 675587 333099
rect 675643 333043 675667 333099
rect 675723 333043 675737 333099
rect 675407 333036 675737 333043
rect 675407 332547 675737 332554
rect 675407 332491 675427 332547
rect 675483 332491 675507 332547
rect 675563 332491 675587 332547
rect 675643 332491 675667 332547
rect 675723 332491 675737 332547
rect 675407 332484 675737 332491
rect 675407 331903 675737 331910
rect 675407 331847 675427 331903
rect 675483 331847 675507 331903
rect 675563 331847 675587 331903
rect 675643 331847 675667 331903
rect 675723 331847 675737 331903
rect 675407 331840 675737 331847
rect 675407 331259 675737 331266
rect 675407 331203 675427 331259
rect 675483 331203 675507 331259
rect 675563 331203 675587 331259
rect 675643 331203 675667 331259
rect 675723 331203 675737 331259
rect 675407 331196 675737 331203
rect 675407 330063 675737 330070
rect 675407 330007 675427 330063
rect 675483 330007 675507 330063
rect 675563 330007 675587 330063
rect 675643 330007 675667 330063
rect 675723 330007 675737 330063
rect 675407 330000 675737 330007
rect 675407 328223 675737 328230
rect 675407 328167 675427 328223
rect 675483 328167 675507 328223
rect 675563 328167 675587 328223
rect 675643 328167 675667 328223
rect 675723 328167 675737 328223
rect 675407 328160 675737 328167
rect 675407 327579 675737 327586
rect 675407 327523 675427 327579
rect 675483 327523 675507 327579
rect 675563 327523 675587 327579
rect 675643 327523 675667 327579
rect 675723 327523 675737 327579
rect 675407 327516 675737 327523
rect 675407 326383 675737 326390
rect 675407 326327 675427 326383
rect 675483 326327 675507 326383
rect 675563 326327 675587 326383
rect 675643 326327 675667 326383
rect 675723 326327 675737 326383
rect 675407 326320 675737 326327
rect 41863 326273 42193 326280
rect 41863 326217 41883 326273
rect 41939 326217 41963 326273
rect 42019 326217 42043 326273
rect 42099 326217 42123 326273
rect 42179 326217 42193 326273
rect 41863 326210 42193 326217
rect 41863 325077 42193 325084
rect 41863 325021 41883 325077
rect 41939 325021 41963 325077
rect 42019 325021 42043 325077
rect 42099 325021 42123 325077
rect 42179 325021 42193 325077
rect 41863 325014 42193 325021
rect 41863 324433 42193 324440
rect 41863 324377 41883 324433
rect 41939 324377 41963 324433
rect 42019 324377 42043 324433
rect 42099 324377 42123 324433
rect 42179 324377 42193 324433
rect 41863 324370 42193 324377
rect 41863 323789 42193 323796
rect 41863 323733 41883 323789
rect 41939 323733 41963 323789
rect 42019 323733 42043 323789
rect 42099 323733 42123 323789
rect 42179 323733 42193 323789
rect 41863 323726 42193 323733
rect 41863 322593 42193 322600
rect 41863 322537 41883 322593
rect 41939 322537 41963 322593
rect 42019 322537 42043 322593
rect 42099 322537 42123 322593
rect 42179 322537 42193 322593
rect 41863 322530 42193 322537
rect 41863 321397 42193 321404
rect 41863 321341 41883 321397
rect 41939 321341 41963 321397
rect 42019 321341 42043 321397
rect 42099 321341 42123 321397
rect 42179 321341 42193 321397
rect 41863 321334 42193 321341
rect 41863 320753 42193 320760
rect 41863 320697 41883 320753
rect 41939 320697 41963 320753
rect 42019 320697 42043 320753
rect 42099 320697 42123 320753
rect 42179 320697 42193 320753
rect 41863 320690 42193 320697
rect 41863 320109 42193 320116
rect 41863 320053 41883 320109
rect 41939 320053 41963 320109
rect 42019 320053 42043 320109
rect 42099 320053 42123 320109
rect 42179 320053 42193 320109
rect 41863 320046 42193 320053
rect 41863 319557 42193 319564
rect 41863 319501 41883 319557
rect 41939 319501 41963 319557
rect 42019 319501 42043 319557
rect 42099 319501 42123 319557
rect 42179 319501 42193 319557
rect 41863 319494 42193 319501
rect 41863 317073 42193 317080
rect 41863 317017 41883 317073
rect 41939 317017 41963 317073
rect 42019 317017 42043 317073
rect 42099 317017 42123 317073
rect 42179 317017 42193 317073
rect 41863 317010 42193 317017
rect 41863 316429 42193 316436
rect 41863 316373 41883 316429
rect 41939 316373 41963 316429
rect 42019 316373 42043 316429
rect 42099 316373 42123 316429
rect 42179 316373 42193 316429
rect 41863 316366 42193 316373
rect 41863 315785 42193 315792
rect 41863 315729 41883 315785
rect 41939 315729 41963 315785
rect 42019 315729 42043 315785
rect 42099 315729 42123 315785
rect 42179 315729 42193 315785
rect 41863 315722 42193 315729
rect 41863 315233 42193 315240
rect 41863 315177 41883 315233
rect 41939 315177 41963 315233
rect 42019 315177 42043 315233
rect 42099 315177 42123 315233
rect 42179 315177 42193 315233
rect 41863 315170 42193 315177
rect 41863 313393 42193 313400
rect 41863 313337 41883 313393
rect 41939 313337 41963 313393
rect 42019 313337 42043 313393
rect 42099 313337 42123 313393
rect 42179 313337 42193 313393
rect 41863 313330 42193 313337
rect 41863 312749 42193 312756
rect 41863 312693 41883 312749
rect 41939 312693 41963 312749
rect 42019 312693 42043 312749
rect 42099 312693 42123 312749
rect 42179 312693 42193 312749
rect 41863 312686 42193 312693
rect 41863 312105 42193 312112
rect 41863 312049 41883 312105
rect 41939 312049 41963 312105
rect 42019 312049 42043 312105
rect 42099 312049 42123 312105
rect 42179 312049 42193 312105
rect 41863 312042 42193 312049
rect 675407 295551 675737 295558
rect 675407 295495 675427 295551
rect 675483 295495 675507 295551
rect 675563 295495 675587 295551
rect 675643 295495 675667 295551
rect 675723 295495 675737 295551
rect 675407 295488 675737 295495
rect 675407 294907 675737 294914
rect 675407 294851 675427 294907
rect 675483 294851 675507 294907
rect 675563 294851 675587 294907
rect 675643 294851 675667 294907
rect 675723 294851 675737 294907
rect 675407 294844 675737 294851
rect 675407 294263 675737 294270
rect 675407 294207 675427 294263
rect 675483 294207 675507 294263
rect 675563 294207 675587 294263
rect 675643 294207 675667 294263
rect 675723 294207 675737 294263
rect 675407 294200 675737 294207
rect 675407 292423 675737 292430
rect 675407 292367 675427 292423
rect 675483 292367 675507 292423
rect 675563 292367 675587 292423
rect 675643 292367 675667 292423
rect 675723 292367 675737 292423
rect 675407 292360 675737 292367
rect 675407 291871 675737 291878
rect 675407 291815 675427 291871
rect 675483 291815 675507 291871
rect 675563 291815 675587 291871
rect 675643 291815 675667 291871
rect 675723 291815 675737 291871
rect 675407 291808 675737 291815
rect 675407 291227 675737 291234
rect 675407 291171 675427 291227
rect 675483 291171 675507 291227
rect 675563 291171 675587 291227
rect 675643 291171 675667 291227
rect 675723 291171 675737 291227
rect 675407 291164 675737 291171
rect 675407 290583 675737 290590
rect 675407 290527 675427 290583
rect 675483 290527 675507 290583
rect 675563 290527 675587 290583
rect 675643 290527 675667 290583
rect 675723 290527 675737 290583
rect 675407 290520 675737 290527
rect 675407 288099 675737 288106
rect 675407 288043 675427 288099
rect 675483 288043 675507 288099
rect 675563 288043 675587 288099
rect 675643 288043 675667 288099
rect 675723 288043 675737 288099
rect 675407 288036 675737 288043
rect 675407 287547 675737 287554
rect 675407 287491 675427 287547
rect 675483 287491 675507 287547
rect 675563 287491 675587 287547
rect 675643 287491 675667 287547
rect 675723 287491 675737 287547
rect 675407 287484 675737 287491
rect 675407 286903 675737 286910
rect 675407 286847 675427 286903
rect 675483 286847 675507 286903
rect 675563 286847 675587 286903
rect 675643 286847 675667 286903
rect 675723 286847 675737 286903
rect 675407 286840 675737 286847
rect 675407 286259 675737 286266
rect 675407 286203 675427 286259
rect 675483 286203 675507 286259
rect 675563 286203 675587 286259
rect 675643 286203 675667 286259
rect 675723 286203 675737 286259
rect 675407 286196 675737 286203
rect 675407 285063 675737 285070
rect 675407 285007 675427 285063
rect 675483 285007 675507 285063
rect 675563 285007 675587 285063
rect 675643 285007 675667 285063
rect 675723 285007 675737 285063
rect 675407 285000 675737 285007
rect 675407 283223 675737 283230
rect 675407 283167 675427 283223
rect 675483 283167 675507 283223
rect 675563 283167 675587 283223
rect 675643 283167 675667 283223
rect 675723 283167 675737 283223
rect 675407 283160 675737 283167
rect 41863 283073 42193 283080
rect 41863 283017 41883 283073
rect 41939 283017 41963 283073
rect 42019 283017 42043 283073
rect 42099 283017 42123 283073
rect 42179 283017 42193 283073
rect 41863 283010 42193 283017
rect 675407 282579 675737 282586
rect 675407 282523 675427 282579
rect 675483 282523 675507 282579
rect 675563 282523 675587 282579
rect 675643 282523 675667 282579
rect 675723 282523 675737 282579
rect 675407 282516 675737 282523
rect 41863 281877 42193 281884
rect 41863 281821 41883 281877
rect 41939 281821 41963 281877
rect 42019 281821 42043 281877
rect 42099 281821 42123 281877
rect 42179 281821 42193 281877
rect 41863 281814 42193 281821
rect 675407 281383 675737 281390
rect 675407 281327 675427 281383
rect 675483 281327 675507 281383
rect 675563 281327 675587 281383
rect 675643 281327 675667 281383
rect 675723 281327 675737 281383
rect 675407 281320 675737 281327
rect 41863 281233 42193 281240
rect 41863 281177 41883 281233
rect 41939 281177 41963 281233
rect 42019 281177 42043 281233
rect 42099 281177 42123 281233
rect 42179 281177 42193 281233
rect 41863 281170 42193 281177
rect 41863 280589 42193 280596
rect 41863 280533 41883 280589
rect 41939 280533 41963 280589
rect 42019 280533 42043 280589
rect 42099 280533 42123 280589
rect 42179 280533 42193 280589
rect 41863 280526 42193 280533
rect 41863 279393 42193 279400
rect 41863 279337 41883 279393
rect 41939 279337 41963 279393
rect 42019 279337 42043 279393
rect 42099 279337 42123 279393
rect 42179 279337 42193 279393
rect 41863 279330 42193 279337
rect 41863 278197 42193 278204
rect 41863 278141 41883 278197
rect 41939 278141 41963 278197
rect 42019 278141 42043 278197
rect 42099 278141 42123 278197
rect 42179 278141 42193 278197
rect 41863 278134 42193 278141
rect 41863 277553 42193 277560
rect 41863 277497 41883 277553
rect 41939 277497 41963 277553
rect 42019 277497 42043 277553
rect 42099 277497 42123 277553
rect 42179 277497 42193 277553
rect 41863 277490 42193 277497
rect 41863 276909 42193 276916
rect 41863 276853 41883 276909
rect 41939 276853 41963 276909
rect 42019 276853 42043 276909
rect 42099 276853 42123 276909
rect 42179 276853 42193 276909
rect 41863 276846 42193 276853
rect 41863 276357 42193 276364
rect 41863 276301 41883 276357
rect 41939 276301 41963 276357
rect 42019 276301 42043 276357
rect 42099 276301 42123 276357
rect 42179 276301 42193 276357
rect 41863 276294 42193 276301
rect 41863 273873 42193 273880
rect 41863 273817 41883 273873
rect 41939 273817 41963 273873
rect 42019 273817 42043 273873
rect 42099 273817 42123 273873
rect 42179 273817 42193 273873
rect 41863 273810 42193 273817
rect 41863 273229 42193 273236
rect 41863 273173 41883 273229
rect 41939 273173 41963 273229
rect 42019 273173 42043 273229
rect 42099 273173 42123 273229
rect 42179 273173 42193 273229
rect 41863 273166 42193 273173
rect 41863 272585 42193 272592
rect 41863 272529 41883 272585
rect 41939 272529 41963 272585
rect 42019 272529 42043 272585
rect 42099 272529 42123 272585
rect 42179 272529 42193 272585
rect 41863 272522 42193 272529
rect 41863 272033 42193 272040
rect 41863 271977 41883 272033
rect 41939 271977 41963 272033
rect 42019 271977 42043 272033
rect 42099 271977 42123 272033
rect 42179 271977 42193 272033
rect 41863 271970 42193 271977
rect 41863 270193 42193 270200
rect 41863 270137 41883 270193
rect 41939 270137 41963 270193
rect 42019 270137 42043 270193
rect 42099 270137 42123 270193
rect 42179 270137 42193 270193
rect 41863 270130 42193 270137
rect 41863 269549 42193 269556
rect 41863 269493 41883 269549
rect 41939 269493 41963 269549
rect 42019 269493 42043 269549
rect 42099 269493 42123 269549
rect 42179 269493 42193 269549
rect 41863 269486 42193 269493
rect 41863 268905 42193 268912
rect 41863 268849 41883 268905
rect 41939 268849 41963 268905
rect 42019 268849 42043 268905
rect 42099 268849 42123 268905
rect 42179 268849 42193 268905
rect 41863 268842 42193 268849
rect 675407 250551 675737 250558
rect 675407 250495 675427 250551
rect 675483 250495 675507 250551
rect 675563 250495 675587 250551
rect 675643 250495 675667 250551
rect 675723 250495 675737 250551
rect 675407 250488 675737 250495
rect 675407 249907 675737 249914
rect 675407 249851 675427 249907
rect 675483 249851 675507 249907
rect 675563 249851 675587 249907
rect 675643 249851 675667 249907
rect 675723 249851 675737 249907
rect 675407 249844 675737 249851
rect 675407 249263 675737 249270
rect 675407 249207 675427 249263
rect 675483 249207 675507 249263
rect 675563 249207 675587 249263
rect 675643 249207 675667 249263
rect 675723 249207 675737 249263
rect 675407 249200 675737 249207
rect 675407 247423 675737 247430
rect 675407 247367 675427 247423
rect 675483 247367 675507 247423
rect 675563 247367 675587 247423
rect 675643 247367 675667 247423
rect 675723 247367 675737 247423
rect 675407 247360 675737 247367
rect 675407 246871 675737 246878
rect 675407 246815 675427 246871
rect 675483 246815 675507 246871
rect 675563 246815 675587 246871
rect 675643 246815 675667 246871
rect 675723 246815 675737 246871
rect 675407 246808 675737 246815
rect 675407 246227 675737 246234
rect 675407 246171 675427 246227
rect 675483 246171 675507 246227
rect 675563 246171 675587 246227
rect 675643 246171 675667 246227
rect 675723 246171 675737 246227
rect 675407 246164 675737 246171
rect 675407 245583 675737 245590
rect 675407 245527 675427 245583
rect 675483 245527 675507 245583
rect 675563 245527 675587 245583
rect 675643 245527 675667 245583
rect 675723 245527 675737 245583
rect 675407 245520 675737 245527
rect 675407 243099 675737 243106
rect 675407 243043 675427 243099
rect 675483 243043 675507 243099
rect 675563 243043 675587 243099
rect 675643 243043 675667 243099
rect 675723 243043 675737 243099
rect 675407 243036 675737 243043
rect 675407 242547 675737 242554
rect 675407 242491 675427 242547
rect 675483 242491 675507 242547
rect 675563 242491 675587 242547
rect 675643 242491 675667 242547
rect 675723 242491 675737 242547
rect 675407 242484 675737 242491
rect 675407 241903 675737 241910
rect 675407 241847 675427 241903
rect 675483 241847 675507 241903
rect 675563 241847 675587 241903
rect 675643 241847 675667 241903
rect 675723 241847 675737 241903
rect 675407 241840 675737 241847
rect 675407 241259 675737 241266
rect 675407 241203 675427 241259
rect 675483 241203 675507 241259
rect 675563 241203 675587 241259
rect 675643 241203 675667 241259
rect 675723 241203 675737 241259
rect 675407 241196 675737 241203
rect 675407 240063 675737 240070
rect 675407 240007 675427 240063
rect 675483 240007 675507 240063
rect 675563 240007 675587 240063
rect 675643 240007 675667 240063
rect 675723 240007 675737 240063
rect 675407 240000 675737 240007
rect 41863 239873 42193 239880
rect 41863 239817 41883 239873
rect 41939 239817 41963 239873
rect 42019 239817 42043 239873
rect 42099 239817 42123 239873
rect 42179 239817 42193 239873
rect 41863 239810 42193 239817
rect 41863 238677 42193 238684
rect 41863 238621 41883 238677
rect 41939 238621 41963 238677
rect 42019 238621 42043 238677
rect 42099 238621 42123 238677
rect 42179 238621 42193 238677
rect 41863 238614 42193 238621
rect 675407 238223 675737 238230
rect 675407 238167 675427 238223
rect 675483 238167 675507 238223
rect 675563 238167 675587 238223
rect 675643 238167 675667 238223
rect 675723 238167 675737 238223
rect 675407 238160 675737 238167
rect 41863 238033 42193 238040
rect 41863 237977 41883 238033
rect 41939 237977 41963 238033
rect 42019 237977 42043 238033
rect 42099 237977 42123 238033
rect 42179 237977 42193 238033
rect 41863 237970 42193 237977
rect 675407 237579 675737 237586
rect 675407 237523 675427 237579
rect 675483 237523 675507 237579
rect 675563 237523 675587 237579
rect 675643 237523 675667 237579
rect 675723 237523 675737 237579
rect 675407 237516 675737 237523
rect 675407 236383 675737 236390
rect 675407 236327 675427 236383
rect 675483 236327 675507 236383
rect 675563 236327 675587 236383
rect 675643 236327 675667 236383
rect 675723 236327 675737 236383
rect 675407 236320 675737 236327
rect 41863 236193 42193 236200
rect 41863 236137 41883 236193
rect 41939 236137 41963 236193
rect 42019 236137 42043 236193
rect 42099 236137 42123 236193
rect 42179 236137 42193 236193
rect 41863 236130 42193 236137
rect 41863 234997 42193 235004
rect 41863 234941 41883 234997
rect 41939 234941 41963 234997
rect 42019 234941 42043 234997
rect 42099 234941 42123 234997
rect 42179 234941 42193 234997
rect 41863 234934 42193 234941
rect 41863 234353 42193 234360
rect 41863 234297 41883 234353
rect 41939 234297 41963 234353
rect 42019 234297 42043 234353
rect 42099 234297 42123 234353
rect 42179 234297 42193 234353
rect 41863 234290 42193 234297
rect 41863 233709 42193 233716
rect 41863 233653 41883 233709
rect 41939 233653 41963 233709
rect 42019 233653 42043 233709
rect 42099 233653 42123 233709
rect 42179 233653 42193 233709
rect 41863 233646 42193 233653
rect 41863 233157 42193 233164
rect 41863 233101 41883 233157
rect 41939 233101 41963 233157
rect 42019 233101 42043 233157
rect 42099 233101 42123 233157
rect 42179 233101 42193 233157
rect 41863 233094 42193 233101
rect 41863 230673 42193 230680
rect 41863 230617 41883 230673
rect 41939 230617 41963 230673
rect 42019 230617 42043 230673
rect 42099 230617 42123 230673
rect 42179 230617 42193 230673
rect 41863 230610 42193 230617
rect 41863 230029 42193 230036
rect 41863 229973 41883 230029
rect 41939 229973 41963 230029
rect 42019 229973 42043 230029
rect 42099 229973 42123 230029
rect 42179 229973 42193 230029
rect 41863 229966 42193 229973
rect 41863 229385 42193 229392
rect 41863 229329 41883 229385
rect 41939 229329 41963 229385
rect 42019 229329 42043 229385
rect 42099 229329 42123 229385
rect 42179 229329 42193 229385
rect 41863 229322 42193 229329
rect 41863 228833 42193 228840
rect 41863 228777 41883 228833
rect 41939 228777 41963 228833
rect 42019 228777 42043 228833
rect 42099 228777 42123 228833
rect 42179 228777 42193 228833
rect 41863 228770 42193 228777
rect 41863 226993 42193 227000
rect 41863 226937 41883 226993
rect 41939 226937 41963 226993
rect 42019 226937 42043 226993
rect 42099 226937 42123 226993
rect 42179 226937 42193 226993
rect 41863 226930 42193 226937
rect 41863 226349 42193 226356
rect 41863 226293 41883 226349
rect 41939 226293 41963 226349
rect 42019 226293 42043 226349
rect 42099 226293 42123 226349
rect 42179 226293 42193 226349
rect 41863 226286 42193 226293
rect 41863 225705 42193 225712
rect 41863 225649 41883 225705
rect 41939 225649 41963 225705
rect 42019 225649 42043 225705
rect 42099 225649 42123 225705
rect 42179 225649 42193 225705
rect 41863 225642 42193 225649
rect 675407 205351 675737 205358
rect 675407 205295 675427 205351
rect 675483 205295 675507 205351
rect 675563 205295 675587 205351
rect 675643 205295 675667 205351
rect 675723 205295 675737 205351
rect 675407 205288 675737 205295
rect 675407 204707 675737 204714
rect 675407 204651 675427 204707
rect 675483 204651 675507 204707
rect 675563 204651 675587 204707
rect 675643 204651 675667 204707
rect 675723 204651 675737 204707
rect 675407 204644 675737 204651
rect 675407 204063 675737 204070
rect 675407 204007 675427 204063
rect 675483 204007 675507 204063
rect 675563 204007 675587 204063
rect 675643 204007 675667 204063
rect 675723 204007 675737 204063
rect 675407 204000 675737 204007
rect 675407 202223 675737 202230
rect 675407 202167 675427 202223
rect 675483 202167 675507 202223
rect 675563 202167 675587 202223
rect 675643 202167 675667 202223
rect 675723 202167 675737 202223
rect 675407 202160 675737 202167
rect 675407 201671 675737 201678
rect 675407 201615 675427 201671
rect 675483 201615 675507 201671
rect 675563 201615 675587 201671
rect 675643 201615 675667 201671
rect 675723 201615 675737 201671
rect 675407 201608 675737 201615
rect 675407 201027 675737 201034
rect 675407 200971 675427 201027
rect 675483 200971 675507 201027
rect 675563 200971 675587 201027
rect 675643 200971 675667 201027
rect 675723 200971 675737 201027
rect 675407 200964 675737 200971
rect 675407 200383 675737 200390
rect 675407 200327 675427 200383
rect 675483 200327 675507 200383
rect 675563 200327 675587 200383
rect 675643 200327 675667 200383
rect 675723 200327 675737 200383
rect 675407 200320 675737 200327
rect 675407 197899 675737 197906
rect 675407 197843 675427 197899
rect 675483 197843 675507 197899
rect 675563 197843 675587 197899
rect 675643 197843 675667 197899
rect 675723 197843 675737 197899
rect 675407 197836 675737 197843
rect 675407 197347 675737 197354
rect 675407 197291 675427 197347
rect 675483 197291 675507 197347
rect 675563 197291 675587 197347
rect 675643 197291 675667 197347
rect 675723 197291 675737 197347
rect 675407 197284 675737 197291
rect 675407 196703 675737 196710
rect 41863 196673 42193 196680
rect 41863 196617 41883 196673
rect 41939 196617 41963 196673
rect 42019 196617 42043 196673
rect 42099 196617 42123 196673
rect 42179 196617 42193 196673
rect 675407 196647 675427 196703
rect 675483 196647 675507 196703
rect 675563 196647 675587 196703
rect 675643 196647 675667 196703
rect 675723 196647 675737 196703
rect 675407 196640 675737 196647
rect 41863 196610 42193 196617
rect 675407 196059 675737 196066
rect 675407 196003 675427 196059
rect 675483 196003 675507 196059
rect 675563 196003 675587 196059
rect 675643 196003 675667 196059
rect 675723 196003 675737 196059
rect 675407 195996 675737 196003
rect 41863 195477 42193 195484
rect 41863 195421 41883 195477
rect 41939 195421 41963 195477
rect 42019 195421 42043 195477
rect 42099 195421 42123 195477
rect 42179 195421 42193 195477
rect 41863 195414 42193 195421
rect 675407 194863 675737 194870
rect 41863 194833 42193 194840
rect 41863 194777 41883 194833
rect 41939 194777 41963 194833
rect 42019 194777 42043 194833
rect 42099 194777 42123 194833
rect 42179 194777 42193 194833
rect 675407 194807 675427 194863
rect 675483 194807 675507 194863
rect 675563 194807 675587 194863
rect 675643 194807 675667 194863
rect 675723 194807 675737 194863
rect 675407 194800 675737 194807
rect 41863 194770 42193 194777
rect 675407 193023 675737 193030
rect 41863 192993 42193 193000
rect 41863 192937 41883 192993
rect 41939 192937 41963 192993
rect 42019 192937 42043 192993
rect 42099 192937 42123 192993
rect 42179 192937 42193 192993
rect 675407 192967 675427 193023
rect 675483 192967 675507 193023
rect 675563 192967 675587 193023
rect 675643 192967 675667 193023
rect 675723 192967 675737 193023
rect 675407 192960 675737 192967
rect 41863 192930 42193 192937
rect 675407 192379 675737 192386
rect 675407 192323 675427 192379
rect 675483 192323 675507 192379
rect 675563 192323 675587 192379
rect 675643 192323 675667 192379
rect 675723 192323 675737 192379
rect 675407 192316 675737 192323
rect 41863 191797 42193 191804
rect 41863 191741 41883 191797
rect 41939 191741 41963 191797
rect 42019 191741 42043 191797
rect 42099 191741 42123 191797
rect 42179 191741 42193 191797
rect 41863 191734 42193 191741
rect 675407 191183 675737 191190
rect 41863 191153 42193 191160
rect 41863 191097 41883 191153
rect 41939 191097 41963 191153
rect 42019 191097 42043 191153
rect 42099 191097 42123 191153
rect 42179 191097 42193 191153
rect 675407 191127 675427 191183
rect 675483 191127 675507 191183
rect 675563 191127 675587 191183
rect 675643 191127 675667 191183
rect 675723 191127 675737 191183
rect 675407 191120 675737 191127
rect 41863 191090 42193 191097
rect 41863 190509 42193 190516
rect 41863 190453 41883 190509
rect 41939 190453 41963 190509
rect 42019 190453 42043 190509
rect 42099 190453 42123 190509
rect 42179 190453 42193 190509
rect 41863 190446 42193 190453
rect 41863 189957 42193 189964
rect 41863 189901 41883 189957
rect 41939 189901 41963 189957
rect 42019 189901 42043 189957
rect 42099 189901 42123 189957
rect 42179 189901 42193 189957
rect 41863 189894 42193 189901
rect 41863 187473 42193 187480
rect 41863 187417 41883 187473
rect 41939 187417 41963 187473
rect 42019 187417 42043 187473
rect 42099 187417 42123 187473
rect 42179 187417 42193 187473
rect 41863 187410 42193 187417
rect 41863 186829 42193 186836
rect 41863 186773 41883 186829
rect 41939 186773 41963 186829
rect 42019 186773 42043 186829
rect 42099 186773 42123 186829
rect 42179 186773 42193 186829
rect 41863 186766 42193 186773
rect 41863 186185 42193 186192
rect 41863 186129 41883 186185
rect 41939 186129 41963 186185
rect 42019 186129 42043 186185
rect 42099 186129 42123 186185
rect 42179 186129 42193 186185
rect 41863 186122 42193 186129
rect 41863 185633 42193 185640
rect 41863 185577 41883 185633
rect 41939 185577 41963 185633
rect 42019 185577 42043 185633
rect 42099 185577 42123 185633
rect 42179 185577 42193 185633
rect 41863 185570 42193 185577
rect 41863 183793 42193 183800
rect 41863 183737 41883 183793
rect 41939 183737 41963 183793
rect 42019 183737 42043 183793
rect 42099 183737 42123 183793
rect 42179 183737 42193 183793
rect 41863 183730 42193 183737
rect 41863 183149 42193 183156
rect 41863 183093 41883 183149
rect 41939 183093 41963 183149
rect 42019 183093 42043 183149
rect 42099 183093 42123 183149
rect 42179 183093 42193 183149
rect 41863 183086 42193 183093
rect 41863 182505 42193 182512
rect 41863 182449 41883 182505
rect 41939 182449 41963 182505
rect 42019 182449 42043 182505
rect 42099 182449 42123 182505
rect 42179 182449 42193 182505
rect 41863 182442 42193 182449
rect 675407 160351 675737 160358
rect 675407 160295 675427 160351
rect 675483 160295 675507 160351
rect 675563 160295 675587 160351
rect 675643 160295 675667 160351
rect 675723 160295 675737 160351
rect 675407 160288 675737 160295
rect 675407 159707 675737 159714
rect 675407 159651 675427 159707
rect 675483 159651 675507 159707
rect 675563 159651 675587 159707
rect 675643 159651 675667 159707
rect 675723 159651 675737 159707
rect 675407 159644 675737 159651
rect 675407 159063 675737 159070
rect 675407 159007 675427 159063
rect 675483 159007 675507 159063
rect 675563 159007 675587 159063
rect 675643 159007 675667 159063
rect 675723 159007 675737 159063
rect 675407 159000 675737 159007
rect 675407 157223 675737 157230
rect 675407 157167 675427 157223
rect 675483 157167 675507 157223
rect 675563 157167 675587 157223
rect 675643 157167 675667 157223
rect 675723 157167 675737 157223
rect 675407 157160 675737 157167
rect 675407 156671 675737 156678
rect 675407 156615 675427 156671
rect 675483 156615 675507 156671
rect 675563 156615 675587 156671
rect 675643 156615 675667 156671
rect 675723 156615 675737 156671
rect 675407 156608 675737 156615
rect 675407 156027 675737 156034
rect 675407 155971 675427 156027
rect 675483 155971 675507 156027
rect 675563 155971 675587 156027
rect 675643 155971 675667 156027
rect 675723 155971 675737 156027
rect 675407 155964 675737 155971
rect 675407 155383 675737 155390
rect 675407 155327 675427 155383
rect 675483 155327 675507 155383
rect 675563 155327 675587 155383
rect 675643 155327 675667 155383
rect 675723 155327 675737 155383
rect 675407 155320 675737 155327
rect 675407 152899 675737 152906
rect 675407 152843 675427 152899
rect 675483 152843 675507 152899
rect 675563 152843 675587 152899
rect 675643 152843 675667 152899
rect 675723 152843 675737 152899
rect 675407 152836 675737 152843
rect 675407 152347 675737 152354
rect 675407 152291 675427 152347
rect 675483 152291 675507 152347
rect 675563 152291 675587 152347
rect 675643 152291 675667 152347
rect 675723 152291 675737 152347
rect 675407 152284 675737 152291
rect 675407 151703 675737 151710
rect 675407 151647 675427 151703
rect 675483 151647 675507 151703
rect 675563 151647 675587 151703
rect 675643 151647 675667 151703
rect 675723 151647 675737 151703
rect 675407 151640 675737 151647
rect 675407 151059 675737 151066
rect 675407 151003 675427 151059
rect 675483 151003 675507 151059
rect 675563 151003 675587 151059
rect 675643 151003 675667 151059
rect 675723 151003 675737 151059
rect 675407 150996 675737 151003
rect 675407 149863 675737 149870
rect 675407 149807 675427 149863
rect 675483 149807 675507 149863
rect 675563 149807 675587 149863
rect 675643 149807 675667 149863
rect 675723 149807 675737 149863
rect 675407 149800 675737 149807
rect 675407 148023 675737 148030
rect 675407 147967 675427 148023
rect 675483 147967 675507 148023
rect 675563 147967 675587 148023
rect 675643 147967 675667 148023
rect 675723 147967 675737 148023
rect 675407 147960 675737 147967
rect 675407 147379 675737 147386
rect 675407 147323 675427 147379
rect 675483 147323 675507 147379
rect 675563 147323 675587 147379
rect 675643 147323 675667 147379
rect 675723 147323 675737 147379
rect 675407 147316 675737 147323
rect 675407 146183 675737 146190
rect 675407 146127 675427 146183
rect 675483 146127 675507 146183
rect 675563 146127 675587 146183
rect 675643 146127 675667 146183
rect 675723 146127 675737 146183
rect 675407 146120 675737 146127
rect 675407 115151 675737 115158
rect 675407 115095 675427 115151
rect 675483 115095 675507 115151
rect 675563 115095 675587 115151
rect 675643 115095 675667 115151
rect 675723 115095 675737 115151
rect 675407 115088 675737 115095
rect 675407 114507 675737 114514
rect 675407 114451 675427 114507
rect 675483 114451 675507 114507
rect 675563 114451 675587 114507
rect 675643 114451 675667 114507
rect 675723 114451 675737 114507
rect 675407 114444 675737 114451
rect 675407 113863 675737 113870
rect 675407 113807 675427 113863
rect 675483 113807 675507 113863
rect 675563 113807 675587 113863
rect 675643 113807 675667 113863
rect 675723 113807 675737 113863
rect 675407 113800 675737 113807
rect 675407 112023 675737 112030
rect 675407 111967 675427 112023
rect 675483 111967 675507 112023
rect 675563 111967 675587 112023
rect 675643 111967 675667 112023
rect 675723 111967 675737 112023
rect 675407 111960 675737 111967
rect 675407 111471 675737 111478
rect 675407 111415 675427 111471
rect 675483 111415 675507 111471
rect 675563 111415 675587 111471
rect 675643 111415 675667 111471
rect 675723 111415 675737 111471
rect 675407 111408 675737 111415
rect 675407 110827 675737 110834
rect 675407 110771 675427 110827
rect 675483 110771 675507 110827
rect 675563 110771 675587 110827
rect 675643 110771 675667 110827
rect 675723 110771 675737 110827
rect 675407 110764 675737 110771
rect 675407 110183 675737 110190
rect 675407 110127 675427 110183
rect 675483 110127 675507 110183
rect 675563 110127 675587 110183
rect 675643 110127 675667 110183
rect 675723 110127 675737 110183
rect 675407 110120 675737 110127
rect 675407 107699 675737 107706
rect 675407 107643 675427 107699
rect 675483 107643 675507 107699
rect 675563 107643 675587 107699
rect 675643 107643 675667 107699
rect 675723 107643 675737 107699
rect 675407 107636 675737 107643
rect 675407 107147 675737 107154
rect 675407 107091 675427 107147
rect 675483 107091 675507 107147
rect 675563 107091 675587 107147
rect 675643 107091 675667 107147
rect 675723 107091 675737 107147
rect 675407 107084 675737 107091
rect 675407 106503 675737 106510
rect 675407 106447 675427 106503
rect 675483 106447 675507 106503
rect 675563 106447 675587 106503
rect 675643 106447 675667 106503
rect 675723 106447 675737 106503
rect 675407 106440 675737 106447
rect 675407 105859 675737 105866
rect 675407 105803 675427 105859
rect 675483 105803 675507 105859
rect 675563 105803 675587 105859
rect 675643 105803 675667 105859
rect 675723 105803 675737 105859
rect 675407 105796 675737 105803
rect 675407 104663 675737 104670
rect 675407 104607 675427 104663
rect 675483 104607 675507 104663
rect 675563 104607 675587 104663
rect 675643 104607 675667 104663
rect 675723 104607 675737 104663
rect 675407 104600 675737 104607
rect 675407 102823 675737 102830
rect 675407 102767 675427 102823
rect 675483 102767 675507 102823
rect 675563 102767 675587 102823
rect 675643 102767 675667 102823
rect 675723 102767 675737 102823
rect 675407 102760 675737 102767
rect 675407 102179 675737 102186
rect 675407 102123 675427 102179
rect 675483 102123 675507 102179
rect 675563 102123 675587 102179
rect 675643 102123 675667 102179
rect 675723 102123 675737 102179
rect 675407 102116 675737 102123
rect 675407 100983 675737 100990
rect 675407 100927 675427 100983
rect 675483 100927 675507 100983
rect 675563 100927 675587 100983
rect 675643 100927 675667 100983
rect 675723 100927 675737 100983
rect 675407 100920 675737 100927
rect 145825 40974 145891 40977
rect 145825 40972 148252 40974
rect 145825 40916 145830 40972
rect 145886 40916 148252 40972
rect 145825 40914 148252 40916
rect 202708 40973 202778 40978
rect 202708 40971 203064 40973
rect 202708 40915 202715 40971
rect 202771 40915 203064 40971
rect 205919 40970 205989 40977
rect 145825 40911 145891 40914
rect 202708 40913 203064 40915
rect 205764 40914 205926 40970
rect 205982 40914 205989 40970
rect 202708 40908 202778 40913
rect 205764 40910 205989 40914
rect 205919 40907 205989 40910
rect 311308 40973 311378 40978
rect 315488 40974 315558 40981
rect 315488 40973 315495 40974
rect 311308 40971 312684 40973
rect 311308 40915 311315 40971
rect 311371 40915 312684 40971
rect 311308 40913 312684 40915
rect 315360 40918 315495 40973
rect 315551 40918 315558 40974
rect 315360 40913 315558 40918
rect 311308 40908 311378 40913
rect 315488 40911 315558 40913
rect 366108 40973 366178 40978
rect 366108 40971 367484 40973
rect 366108 40915 366115 40971
rect 366171 40915 367484 40971
rect 370293 40970 370363 40977
rect 370293 40969 370300 40970
rect 366108 40913 367484 40915
rect 370159 40914 370300 40969
rect 370356 40914 370363 40970
rect 366108 40908 366178 40913
rect 370159 40909 370363 40914
rect 370293 40907 370363 40909
rect 420908 40973 420978 40978
rect 475708 40973 475778 40978
rect 420908 40971 422262 40973
rect 420908 40915 420915 40971
rect 420971 40915 422262 40971
rect 475708 40971 477055 40973
rect 425106 40964 425176 40965
rect 420908 40913 422262 40915
rect 424960 40958 425176 40964
rect 420908 40908 420978 40913
rect 424960 40904 425113 40958
rect 425106 40902 425113 40904
rect 425169 40902 425176 40958
rect 475708 40915 475715 40971
rect 475771 40915 477055 40971
rect 479906 40972 479976 40979
rect 479906 40969 479913 40972
rect 475708 40913 477055 40915
rect 479767 40916 479913 40969
rect 479969 40916 479976 40972
rect 475708 40908 475778 40913
rect 479767 40909 479976 40916
rect 530508 40973 530578 40978
rect 530508 40971 531856 40973
rect 530508 40915 530515 40971
rect 530571 40915 531856 40971
rect 534763 40963 534833 40967
rect 530508 40913 531856 40915
rect 534569 40960 534833 40963
rect 530508 40908 530578 40913
rect 534569 40904 534770 40960
rect 534826 40904 534833 40960
rect 534569 40903 534833 40904
rect 425106 40895 425176 40902
rect 534763 40897 534833 40903
rect 133094 40158 144010 40218
rect 133094 39984 133154 40158
rect 143407 40095 143519 40097
rect 143402 40090 143524 40095
rect 143402 40034 143435 40090
rect 143491 40034 143524 40090
rect 143402 39992 143524 40034
rect 143950 39984 144010 40158
rect 145832 40132 145902 40148
rect 145832 40076 145839 40132
rect 145895 40076 145902 40132
rect 145832 39982 145902 40076
rect 148901 40033 149351 40055
rect 148901 39729 149149 40033
rect 149293 39729 149351 40033
rect 148901 31573 149351 39729
rect 149537 40032 149918 40055
rect 149537 39728 149651 40032
rect 149795 39728 149918 40032
rect 149537 38114 149918 39728
rect 149537 37410 149575 38114
rect 149879 37410 149918 38114
rect 149537 37340 149918 37410
rect 203701 40033 204151 40055
rect 203701 39729 203949 40033
rect 204093 39729 204151 40033
rect 148901 30869 148970 31573
rect 149274 30869 149351 31573
rect 148901 30806 149351 30869
rect 203701 31573 204151 39729
rect 204337 40032 204718 40055
rect 204337 39728 204451 40032
rect 204595 39728 204718 40032
rect 204337 38114 204718 39728
rect 204337 37410 204375 38114
rect 204679 37410 204718 38114
rect 204337 37340 204718 37410
rect 313301 40033 313751 40055
rect 313301 39729 313549 40033
rect 313693 39729 313751 40033
rect 203701 30869 203770 31573
rect 204074 30869 204151 31573
rect 203701 30806 204151 30869
rect 313301 31573 313751 39729
rect 313937 40032 314318 40055
rect 313937 39728 314051 40032
rect 314195 39728 314318 40032
rect 313937 38114 314318 39728
rect 313937 37410 313975 38114
rect 314279 37410 314318 38114
rect 313937 37340 314318 37410
rect 368101 40033 368551 40055
rect 368101 39729 368349 40033
rect 368493 39729 368551 40033
rect 313301 30869 313370 31573
rect 313674 30869 313751 31573
rect 313301 30806 313751 30869
rect 368101 31573 368551 39729
rect 368737 40032 369118 40055
rect 368737 39728 368851 40032
rect 368995 39728 369118 40032
rect 368737 38114 369118 39728
rect 368737 37410 368775 38114
rect 369079 37410 369118 38114
rect 368737 37340 369118 37410
rect 422901 40033 423351 40055
rect 422901 39729 423149 40033
rect 423293 39729 423351 40033
rect 368101 30869 368170 31573
rect 368474 30869 368551 31573
rect 368101 30806 368551 30869
rect 422901 31573 423351 39729
rect 423537 40032 423918 40055
rect 423537 39728 423651 40032
rect 423795 39728 423918 40032
rect 423537 38114 423918 39728
rect 423537 37410 423575 38114
rect 423879 37410 423918 38114
rect 423537 37340 423918 37410
rect 477701 40033 478151 40055
rect 477701 39729 477949 40033
rect 478093 39729 478151 40033
rect 422901 30869 422970 31573
rect 423274 30869 423351 31573
rect 422901 30806 423351 30869
rect 477701 31573 478151 39729
rect 478337 40032 478718 40055
rect 478337 39728 478451 40032
rect 478595 39728 478718 40032
rect 478337 38114 478718 39728
rect 478337 37410 478375 38114
rect 478679 37410 478718 38114
rect 478337 37340 478718 37410
rect 532501 40033 532951 40055
rect 532501 39729 532749 40033
rect 532893 39729 532951 40033
rect 477701 30869 477770 31573
rect 478074 30869 478151 31573
rect 477701 30806 478151 30869
rect 532501 31573 532951 39729
rect 533137 40032 533518 40055
rect 533137 39728 533251 40032
rect 533395 39728 533518 40032
rect 533137 38114 533518 39728
rect 533137 37410 533175 38114
rect 533479 37410 533518 38114
rect 533137 37340 533518 37410
rect 532501 30869 532570 31573
rect 532874 30869 532951 31573
rect 532501 30806 532951 30869
<< via3 >>
rect 149149 39729 149293 40033
rect 149651 39728 149795 40032
rect 149575 37410 149879 38114
rect 203949 39729 204093 40033
rect 148970 30869 149274 31573
rect 204451 39728 204595 40032
rect 204375 37410 204679 38114
rect 313549 39729 313693 40033
rect 203770 30869 204074 31573
rect 314051 39728 314195 40032
rect 313975 37410 314279 38114
rect 368349 39729 368493 40033
rect 313370 30869 313674 31573
rect 368851 39728 368995 40032
rect 368775 37410 369079 38114
rect 423149 39729 423293 40033
rect 368170 30869 368474 31573
rect 423651 39728 423795 40032
rect 423575 37410 423879 38114
rect 477949 39729 478093 40033
rect 422970 30869 423274 31573
rect 478451 39728 478595 40032
rect 478375 37410 478679 38114
rect 532749 39729 532893 40033
rect 477770 30869 478074 31573
rect 533251 39728 533395 40032
rect 533175 37410 533479 38114
rect 532570 30869 532874 31573
<< metal4 >>
rect 680587 459800 681277 459993
rect 688881 459800 688947 474800
rect 0 455645 4843 456094
rect 28653 440800 28719 455800
rect 32933 455546 33623 455800
rect 36323 455607 37013 455799
rect 38503 455546 39593 455800
rect 149134 40033 149314 40149
rect 149134 39729 149149 40033
rect 149293 39729 149314 40033
rect 149134 39704 149314 39729
rect 149634 40032 149814 40149
rect 149634 39728 149651 40032
rect 149795 39728 149814 40032
rect 149634 39704 149814 39728
rect 203934 40033 204114 40148
rect 203934 39729 203949 40033
rect 204093 39729 204114 40033
rect 203934 39704 204114 39729
rect 204434 40032 204614 40148
rect 204434 39728 204451 40032
rect 204595 39728 204614 40032
rect 204434 39704 204614 39728
rect 313534 40033 313714 40148
rect 313534 39729 313549 40033
rect 313693 39729 313714 40033
rect 313534 39704 313714 39729
rect 314034 40032 314214 40148
rect 314034 39728 314051 40032
rect 314195 39728 314214 40032
rect 314034 39704 314214 39728
rect 368334 40033 368514 40148
rect 368334 39729 368349 40033
rect 368493 39729 368514 40033
rect 368334 39704 368514 39729
rect 368834 40032 369014 40148
rect 368834 39728 368851 40032
rect 368995 39728 369014 40032
rect 368834 39704 369014 39728
rect 423134 40033 423314 40148
rect 423134 39729 423149 40033
rect 423293 39729 423314 40033
rect 423134 39704 423314 39729
rect 423634 40032 423814 40148
rect 423634 39728 423651 40032
rect 423795 39728 423814 40032
rect 423634 39704 423814 39728
rect 477934 40033 478114 40148
rect 477934 39729 477949 40033
rect 478093 39729 478114 40033
rect 477934 39704 478114 39729
rect 478434 40032 478614 40148
rect 478434 39728 478451 40032
rect 478595 39728 478614 40032
rect 478434 39704 478614 39728
rect 532734 40033 532914 40148
rect 532734 39729 532749 40033
rect 532893 39729 532914 40033
rect 532734 39704 532914 39729
rect 533234 40032 533414 40148
rect 533234 39728 533251 40032
rect 533395 39728 533414 40032
rect 533234 39704 533414 39728
rect 149563 38114 149891 38153
rect 149563 37410 149575 38114
rect 149879 37410 149891 38114
rect 149563 37372 149891 37410
rect 204363 38114 204691 38153
rect 204363 37410 204375 38114
rect 204679 37410 204691 38114
rect 204363 37372 204691 37410
rect 313963 38114 314291 38153
rect 313963 37410 313975 38114
rect 314279 37410 314291 38114
rect 313963 37372 314291 37410
rect 368763 38114 369091 38153
rect 368763 37410 368775 38114
rect 369079 37410 369091 38114
rect 368763 37372 369091 37410
rect 423563 38114 423891 38153
rect 423563 37410 423575 38114
rect 423879 37410 423891 38114
rect 423563 37372 423891 37410
rect 478363 38114 478691 38153
rect 478363 37410 478375 38114
rect 478679 37410 478691 38114
rect 478363 37372 478691 37410
rect 533163 38114 533491 38153
rect 533163 37410 533175 38114
rect 533479 37410 533491 38114
rect 533163 37372 533491 37410
rect 132600 36323 132792 37013
rect 132600 30753 132854 31683
rect 148940 31573 149305 31600
rect 148940 30869 148970 31573
rect 149274 30869 149305 31573
rect 148940 30843 149305 30869
rect 203740 31573 204105 31600
rect 203740 30869 203770 31573
rect 204074 30869 204105 31573
rect 203740 30843 204105 30869
rect 313340 31573 313705 31600
rect 313340 30869 313370 31573
rect 313674 30869 313705 31573
rect 313340 30843 313705 30869
rect 368140 31573 368505 31600
rect 368140 30869 368170 31573
rect 368474 30869 368505 31573
rect 368140 30843 368505 30869
rect 422940 31573 423305 31600
rect 422940 30869 422970 31573
rect 423274 30869 423305 31573
rect 422940 30843 423305 30869
rect 477740 31573 478105 31600
rect 477740 30869 477770 31573
rect 478074 30869 478105 31573
rect 477740 30843 478105 30869
rect 532540 31573 532905 31600
rect 532540 30869 532570 31573
rect 532874 30869 532905 31573
rect 532540 30843 532905 30869
rect 132600 28653 147600 28719
<< metal5 >>
rect 78420 1018512 90960 1031002
rect 129820 1018512 142360 1031002
rect 181220 1018512 193760 1031002
rect 232620 1018512 245160 1031002
rect 284220 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386020 1018512 398560 1031002
rect 475020 1018512 487560 1031002
rect 526420 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628220 1018512 640760 1031002
rect 348400 1007147 348466 1008947
rect 348400 1004968 348466 1005617
rect 348400 1000607 348527 1001257
rect 6598 956420 19088 968960
rect 698512 952840 711002 965380
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876180
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786620 19088 799160
rect 698512 774440 711002 786980
rect 6598 743420 19088 755960
rect 698512 729440 711002 741980
rect 6598 700220 19088 712760
rect 698512 684440 711002 696980
rect 6598 657020 19088 669560
rect 698512 639240 711002 651780
rect 6598 613820 19088 626360
rect 698512 594240 711002 606780
rect 6598 570620 19088 583160
rect 698512 549040 711002 561580
rect 6598 527420 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399820 19088 412360
rect 698512 371840 711002 384380
rect 6598 356620 19088 369160
rect 698512 326640 711002 339180
rect 6598 313420 19088 325960
rect 6598 270220 19088 282760
rect 698512 281640 711002 294180
rect 6598 227020 19088 239560
rect 698512 236640 711002 249180
rect 6598 183820 19088 196360
rect 698512 191440 711002 203980
rect 698512 146440 711002 158980
rect 6811 111610 18975 123778
rect 698512 101240 711002 113780
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19619
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1677077417
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1677077417
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1677077417
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1677077417
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1677077417
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1677077417
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1677077417
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1677077417
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13
timestamp 1677077417
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_14
timestamp 1677077417
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1677077417
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1677077417
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1677077417
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1677077417
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1677077417
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1677077417
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1677077417
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1677077417
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1677077417
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1677077417
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1677077417
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1677077417
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1677077417
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1677077417
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1677077417
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1677077417
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1677077417
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1677077417
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1677077417
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1677077417
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1677077417
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1677077417
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1677077417
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1677077417
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1677077417
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1677077417
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1677077417
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1677077417
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1677077417
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1677077417
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1677077417
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1677077417
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1677077417
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1677077417
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1677077417
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1677077417
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1677077417
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1677077417
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1677077417
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1677077417
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1677077417
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1677077417
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1677077417
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1677077417
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1677077417
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1677077417
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1677077417
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1677077417
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1677077417
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1677077417
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1677077417
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1677077417
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1677077417
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1677077417
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1677077417
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1677077417
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1677077417
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1677077417
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1677077417
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1677077417
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1677077417
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1677077417
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1677077417
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1677077417
transform 1 0 350400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1677077417
transform 1 0 354400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1677077417
transform 1 0 358400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1677077417
transform 1 0 362400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1677077417
transform 1 0 366400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1677077417
transform 1 0 370400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1677077417
transform 1 0 374400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_93
timestamp 1677077417
transform 1 0 378400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_94
timestamp 1677077417
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1677077417
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1677077417
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1677077417
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1677077417
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1677077417
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1677077417
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1677077417
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1677077417
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1677077417
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1677077417
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1677077417
transform 1 0 431800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_107
timestamp 1677077417
transform 1 0 435800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_108
timestamp 1677077417
transform 1 0 439800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_109
timestamp 1677077417
transform 1 0 443800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1677077417
transform 1 0 447800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1677077417
transform 1 0 451800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1677077417
transform 1 0 455800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1677077417
transform 1 0 459800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1677077417
transform 1 0 463800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1677077417
transform 1 0 467800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_116
timestamp 1677077417
transform 1 0 471800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1677077417
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_119
timestamp 1677077417
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_120
timestamp 1677077417
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_121
timestamp 1677077417
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_122
timestamp 1677077417
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1677077417
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1677077417
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1677077417
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_126
timestamp 1677077417
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_127
timestamp 1677077417
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_128
timestamp 1677077417
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_129
timestamp 1677077417
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1677077417
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1677077417
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_133
timestamp 1677077417
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_134
timestamp 1677077417
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1677077417
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1677077417
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1677077417
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1677077417
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_139
timestamp 1677077417
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_140
timestamp 1677077417
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_141
timestamp 1677077417
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_142
timestamp 1677077417
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1677077417
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1677077417
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_146
timestamp 1677077417
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_147
timestamp 1677077417
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_148
timestamp 1677077417
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_149
timestamp 1677077417
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_150
timestamp 1677077417
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1677077417
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_152
timestamp 1677077417
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_153
timestamp 1677077417
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_154
timestamp 1677077417
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_155
timestamp 1677077417
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1677077417
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1677077417
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1677077417
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_160
timestamp 1677077417
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_161
timestamp 1677077417
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_162
timestamp 1677077417
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_163
timestamp 1677077417
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1677077417
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_165
timestamp 1677077417
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_166
timestamp 1677077417
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_167
timestamp 1677077417
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1677077417
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1677077417
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1677077417
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_171
timestamp 1677077417
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_172
timestamp 1677077417
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_173
timestamp 1677077417
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1677077417
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_181
timestamp 1677077417
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_182
timestamp 1677077417
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_183
timestamp 1677077417
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_184
timestamp 1677077417
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1677077417
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_187
timestamp 1677077417
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_188
timestamp 1677077417
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_189
timestamp 1677077417
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_190
timestamp 1677077417
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1677077417
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_198
timestamp 1677077417
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_199
timestamp 1677077417
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_200
timestamp 1677077417
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_201
timestamp 1677077417
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1677077417
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_204
timestamp 1677077417
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_205
timestamp 1677077417
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_206
timestamp 1677077417
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_207
timestamp 1677077417
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1677077417
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_215
timestamp 1677077417
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_216
timestamp 1677077417
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_217
timestamp 1677077417
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_218
timestamp 1677077417
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1677077417
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_221
timestamp 1677077417
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_222
timestamp 1677077417
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_223
timestamp 1677077417
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_224
timestamp 1677077417
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1677077417
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_232
timestamp 1677077417
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_233
timestamp 1677077417
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_234
timestamp 1677077417
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_235
timestamp 1677077417
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1677077417
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_238
timestamp 1677077417
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_239
timestamp 1677077417
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_240
timestamp 1677077417
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_241
timestamp 1677077417
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1677077417
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_249
timestamp 1677077417
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_250
timestamp 1677077417
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_251
timestamp 1677077417
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_252
timestamp 1677077417
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1677077417
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_255
timestamp 1677077417
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_256
timestamp 1677077417
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_257
timestamp 1677077417
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_258
timestamp 1677077417
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1677077417
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_266
timestamp 1677077417
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_267
timestamp 1677077417
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_268
timestamp 1677077417
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_269
timestamp 1677077417
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1677077417
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_272
timestamp 1677077417
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_273
timestamp 1677077417
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_274
timestamp 1677077417
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_275
timestamp 1677077417
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1677077417
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_283
timestamp 1677077417
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_284
timestamp 1677077417
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_285
timestamp 1677077417
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_286
timestamp 1677077417
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1677077417
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_289
timestamp 1677077417
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_290
timestamp 1677077417
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_291
timestamp 1677077417
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_292
timestamp 1677077417
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1677077417
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_300
timestamp 1677077417
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_301
timestamp 1677077417
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_302
timestamp 1677077417
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_303
timestamp 1677077417
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1677077417
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_306
timestamp 1677077417
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_307
timestamp 1677077417
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_308
timestamp 1677077417
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_309
timestamp 1677077417
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1677077417
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_317
timestamp 1677077417
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_318
timestamp 1677077417
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_319
timestamp 1677077417
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_320
timestamp 1677077417
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1677077417
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_323
timestamp 1677077417
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_324
timestamp 1677077417
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_325
timestamp 1677077417
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_326
timestamp 1677077417
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1677077417
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_334
timestamp 1677077417
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_335
timestamp 1677077417
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_336
timestamp 1677077417
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_337
timestamp 1677077417
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1677077417
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_340
timestamp 1677077417
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_341
timestamp 1677077417
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_342
timestamp 1677077417
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_343
timestamp 1677077417
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1677077417
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_351
timestamp 1677077417
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_352
timestamp 1677077417
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_353
timestamp 1677077417
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_354
timestamp 1677077417
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_355
timestamp 1677077417
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1677077417
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_358
timestamp 1677077417
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_359
timestamp 1677077417
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1677077417
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1677077417
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_368
timestamp 1677077417
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_369
timestamp 1677077417
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_370
timestamp 1677077417
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_371
timestamp 1677077417
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_372
timestamp 1677077417
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_373
timestamp 1677077417
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_374
timestamp 1677077417
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1677077417
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1677077417
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1677077417
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1677077417
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1677077417
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_380
timestamp 1677077417
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_381
timestamp 1677077417
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_382
timestamp 1677077417
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1677077417
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1677077417
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1677077417
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_387
timestamp 1677077417
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_388
timestamp 1677077417
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_389
timestamp 1677077417
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_390
timestamp 1677077417
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_391
timestamp 1677077417
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_392
timestamp 1677077417
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1677077417
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1677077417
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1677077417
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_397
timestamp 1677077417
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_398
timestamp 1677077417
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_399
timestamp 1677077417
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_400
timestamp 1677077417
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_401
timestamp 1677077417
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_402
timestamp 1677077417
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1677077417
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1677077417
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_407
timestamp 1677077417
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_408
timestamp 1677077417
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_409
timestamp 1677077417
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_410
timestamp 1677077417
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_411
timestamp 1677077417
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_412
timestamp 1677077417
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_413
timestamp 1677077417
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1677077417
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1677077417
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1677077417
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_418
timestamp 1677077417
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_419
timestamp 1677077417
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_420
timestamp 1677077417
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_421
timestamp 1677077417
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_422
timestamp 1677077417
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_423
timestamp 1677077417
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1677077417
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1677077417
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1677077417
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_428
timestamp 1677077417
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_429
timestamp 1677077417
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_430
timestamp 1677077417
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_431
timestamp 1677077417
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_432
timestamp 1677077417
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_433
timestamp 1677077417
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1677077417
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1677077417
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1677077417
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_438
timestamp 1677077417
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_439
timestamp 1677077417
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_440
timestamp 1677077417
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_441
timestamp 1677077417
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_442
timestamp 1677077417
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_443
timestamp 1677077417
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1677077417
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1677077417
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1677077417
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_448
timestamp 1677077417
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_449
timestamp 1677077417
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_450
timestamp 1677077417
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_451
timestamp 1677077417
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_452
timestamp 1677077417
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_453
timestamp 1677077417
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1677077417
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1677077417
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1677077417
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_458
timestamp 1677077417
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_459
timestamp 1677077417
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_460
timestamp 1677077417
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_461
timestamp 1677077417
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_462
timestamp 1677077417
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_463
timestamp 1677077417
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1677077417
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1677077417
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1677077417
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_468
timestamp 1677077417
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_469
timestamp 1677077417
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_470
timestamp 1677077417
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_471
timestamp 1677077417
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_472
timestamp 1677077417
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_473
timestamp 1677077417
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1677077417
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1677077417
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1677077417
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_478
timestamp 1677077417
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_479
timestamp 1677077417
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_480
timestamp 1677077417
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_481
timestamp 1677077417
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_482
timestamp 1677077417
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_483
timestamp 1677077417
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1677077417
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1677077417
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1677077417
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_488
timestamp 1677077417
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_489
timestamp 1677077417
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_490
timestamp 1677077417
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_491
timestamp 1677077417
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_492
timestamp 1677077417
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_493
timestamp 1677077417
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1677077417
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1677077417
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1677077417
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_498
timestamp 1677077417
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_499
timestamp 1677077417
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_500
timestamp 1677077417
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_501
timestamp 1677077417
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_502
timestamp 1677077417
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_503
timestamp 1677077417
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1677077417
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1677077417
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1677077417
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_508
timestamp 1677077417
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_509
timestamp 1677077417
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_510
timestamp 1677077417
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_511
timestamp 1677077417
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_512
timestamp 1677077417
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_513
timestamp 1677077417
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1677077417
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1677077417
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1677077417
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_518
timestamp 1677077417
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_519
timestamp 1677077417
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_520
timestamp 1677077417
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_521
timestamp 1677077417
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_522
timestamp 1677077417
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_523
timestamp 1677077417
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1677077417
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1677077417
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1677077417
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_528
timestamp 1677077417
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_529
timestamp 1677077417
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_530
timestamp 1677077417
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_531
timestamp 1677077417
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_532
timestamp 1677077417
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_533
timestamp 1677077417
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1677077417
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1677077417
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1677077417
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_538
timestamp 1677077417
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_539
timestamp 1677077417
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_540
timestamp 1677077417
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_541
timestamp 1677077417
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_542
timestamp 1677077417
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_543
timestamp 1677077417
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1677077417
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1677077417
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1677077417
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_548
timestamp 1677077417
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_549
timestamp 1677077417
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_550
timestamp 1677077417
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_551
timestamp 1677077417
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_552
timestamp 1677077417
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_553
timestamp 1677077417
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1677077417
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1677077417
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1677077417
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_558
timestamp 1677077417
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_559
timestamp 1677077417
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_560
timestamp 1677077417
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_561
timestamp 1677077417
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_562
timestamp 1677077417
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_563
timestamp 1677077417
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1677077417
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1677077417
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1677077417
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_568
timestamp 1677077417
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_569
timestamp 1677077417
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1677077417
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_571
timestamp 1677077417
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_572
timestamp 1677077417
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_573
timestamp 1677077417
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1677077417
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1677077417
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1677077417
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_578
timestamp 1677077417
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_579
timestamp 1677077417
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1677077417
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_581
timestamp 1677077417
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_582
timestamp 1677077417
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_583
timestamp 1677077417
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1677077417
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1677077417
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1677077417
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_588
timestamp 1677077417
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_589
timestamp 1677077417
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_590
timestamp 1677077417
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_591
timestamp 1677077417
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_592
timestamp 1677077417
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_593
timestamp 1677077417
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1677077417
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1677077417
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1677077417
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_598
timestamp 1677077417
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1677077417
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1677077417
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_601
timestamp 1677077417
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_602
timestamp 1677077417
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_603
timestamp 1677077417
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_604
timestamp 1677077417
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1677077417
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1677077417
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1677077417
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_608
timestamp 1677077417
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1677077417
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1677077417
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1677077417
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_612
timestamp 1677077417
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1677077417
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1677077417
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1677077417
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1677077417
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1677077417
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1677077417
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1677077417
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_622
timestamp 1677077417
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1677077417
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1677077417
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1677077417
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1677077417
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1677077417
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1677077417
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1677077417
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_631
timestamp 1677077417
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_632
timestamp 1677077417
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1677077417
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1677077417
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1677077417
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1677077417
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1677077417
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1677077417
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1677077417
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_641
timestamp 1677077417
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1677077417
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1677077417
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1677077417
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1677077417
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1677077417
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1677077417
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1677077417
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_650
timestamp 1677077417
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_651
timestamp 1677077417
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1677077417
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1677077417
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1677077417
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1677077417
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_657
timestamp 1677077417
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_658
timestamp 1677077417
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1677077417
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_660
timestamp 1677077417
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1677077417
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1677077417
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1677077417
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1677077417
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1677077417
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1677077417
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1677077417
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_669
timestamp 1677077417
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1677077417
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1677077417
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1677077417
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1677077417
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1677077417
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1677077417
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1677077417
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_678
timestamp 1677077417
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_679
timestamp 1677077417
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1677077417
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1677077417
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1677077417
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1677077417
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_685
timestamp 1677077417
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1677077417
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1677077417
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_688
timestamp 1677077417
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1677077417
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1677077417
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1677077417
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1677077417
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1677077417
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_695
timestamp 1677077417
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_696
timestamp 1677077417
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_697
timestamp 1677077417
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_698
timestamp 1677077417
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1677077417
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1677077417
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1677077417
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1677077417
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1677077417
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1677077417
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1677077417
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_707
timestamp 1677077417
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1677077417
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1677077417
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1677077417
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1677077417
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1677077417
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1677077417
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1677077417
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_716
timestamp 1677077417
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1677077417
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1677077417
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1677077417
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1677077417
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1677077417
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1677077417
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1677077417
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_725
timestamp 1677077417
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_726
timestamp 1677077417
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1677077417
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1677077417
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1677077417
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1677077417
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1677077417
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1677077417
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1677077417
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_735
timestamp 1677077417
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1677077417
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1677077417
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1677077417
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1677077417
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1677077417
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1677077417
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1677077417
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_744
timestamp 1677077417
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_745
timestamp 1677077417
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1677077417
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1677077417
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1677077417
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1677077417
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1677077417
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_752
timestamp 1677077417
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1677077417
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_754
timestamp 1677077417
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1677077417
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1677077417
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1677077417
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1677077417
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1677077417
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1677077417
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1677077417
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_763
timestamp 1677077417
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1677077417
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1677077417
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1677077417
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1677077417
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1677077417
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1677077417
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1677077417
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_772
timestamp 1677077417
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_773
timestamp 1677077417
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1677077417
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1677077417
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1677077417
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1677077417
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_779
timestamp 1677077417
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1677077417
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1677077417
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_782
timestamp 1677077417
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1677077417
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1677077417
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1677077417
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1677077417
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1677077417
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_789
timestamp 1677077417
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_790
timestamp 1677077417
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_791
timestamp 1677077417
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_792
timestamp 1677077417
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1677077417
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1677077417
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1677077417
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1677077417
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_798
timestamp 1677077417
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_799
timestamp 1677077417
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_800
timestamp 1677077417
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_801
timestamp 1677077417
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1677077417
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1677077417
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1677077417
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1677077417
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1677077417
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_808
timestamp 1677077417
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_809
timestamp 1677077417
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_810
timestamp 1677077417
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_811
timestamp 1677077417
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB1
timestamp 1677077417
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB2
timestamp 1677077417
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB3
timestamp 1677077417
transform 1 0 349400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1677077417
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1677077417
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3
timestamp 1677077417
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1677077417
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1677077417
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1677077417
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1677077417
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1677077417
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1677077417
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1677077417
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1677077417
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1677077417
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1677077417
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1677077417
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1677077417
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1677077417
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1677077417
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1677077417
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1677077417
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1677077417
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1677077417
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1677077417
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1677077417
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1677077417
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1677077417
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1677077417
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1677077417
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1677077417
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1677077417
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1677077417
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1677077417
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1677077417
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1677077417
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1677077417
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1677077417
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1677077417
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1677077417
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1677077417
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1677077417
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1677077417
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1677077417
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1677077417
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1677077417
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1677077417
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1677077417
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1677077417
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1677077417
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1677077417
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1677077417
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1677077417
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1677077417
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1677077417
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1677077417
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1677077417
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1677077417
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1677077417
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1677077417
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1677077417
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1677077417
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1677077417
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1677077417
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1677077417
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1677077417
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1677077417
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1677077417
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1677077417
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1677077417
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1677077417
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1677077417
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1677077417
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1677077417
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1677077417
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use chip_io_gpio_connects  chip_io_gpio_connects_0
timestamp 1504095569
transform 0 -1 742000 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_1
timestamp 1504095569
transform 0 -1 640200 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_2
timestamp 1504095569
transform 0 -1 588800 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_3
timestamp 1504095569
transform 0 -1 499800 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_4
timestamp 1504095569
transform 0 -1 398000 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_5
timestamp 1504095569
transform 0 -1 346400 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_6
timestamp 1504095569
transform 0 -1 295000 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_7
timestamp 1504095569
transform 0 -1 243600 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_8
timestamp 1504095569
transform 0 -1 192200 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_9
timestamp 1504095569
transform 1 0 0 0 1 851600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_10
timestamp 1504095569
transform -1 0 717600 0 -1 1070200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_11
timestamp 1504095569
transform 1 0 0 0 1 762400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_12
timestamp 1504095569
transform 1 0 0 0 1 673200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_13
timestamp 1504095569
transform -1 0 717600 0 -1 900400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_14
timestamp 1504095569
transform 1 0 0 0 1 628200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_15
timestamp 1504095569
transform -1 0 717600 0 -1 857200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_16
timestamp 1504095569
transform 1 0 0 0 1 583200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_17
timestamp 1504095569
transform -1 0 717600 0 -1 814000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_18
timestamp 1504095569
transform 1 0 0 0 1 538000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_19
timestamp 1504095569
transform -1 0 717600 0 -1 770800
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_20
timestamp 1504095569
transform 1 0 0 0 1 493000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_21
timestamp 1504095569
transform -1 0 717600 0 -1 727600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_22
timestamp 1504095569
transform -1 0 717600 0 -1 684400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_23
timestamp 1504095569
transform 1 0 0 0 1 447800
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_24
timestamp 1504095569
transform -1 0 717600 0 -1 641200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_25
timestamp 1504095569
transform -1 0 717600 0 -1 513600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_26
timestamp 1504095569
transform 1 0 0 0 1 270600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_27
timestamp 1504095569
transform -1 0 717600 0 -1 470400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_28
timestamp 1504095569
transform 1 0 0 0 1 225400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_29
timestamp 1504095569
transform -1 0 717600 0 -1 427200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_30
timestamp 1504095569
transform 1 0 0 0 1 180400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_31
timestamp 1504095569
transform -1 0 717600 0 -1 384000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_32
timestamp 1504095569
transform 1 0 0 0 1 135400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_33
timestamp 1504095569
transform -1 0 717600 0 -1 340800
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_34
timestamp 1504095569
transform 1 0 0 0 1 90200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_35
timestamp 1504095569
transform -1 0 717600 0 -1 297600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_36
timestamp 1504095569
transform 1 0 0 0 1 45200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_37
timestamp 1504095569
transform 1 0 0 0 1 0
box 675407 99896 675887 115709
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad
timestamp 1677077417
transform -1 0 202400 0 -1 42193
box -143 0 16134 42193
use constant_block  constant_block_0
timestamp 1677077417
transform -1 0 534616 0 1 39652
box 0 496 2800 2224
use constant_block  constant_block_1
timestamp 1677077417
transform -1 0 479816 0 1 39652
box 0 496 2800 2224
use constant_block  constant_block_2
timestamp 1677077417
transform -1 0 425016 0 1 39652
box 0 496 2800 2224
use constant_block  constant_block_3
timestamp 1677077417
transform -1 0 370216 0 1 39652
box 0 496 2800 2224
use constant_block  constant_block_4
timestamp 1677077417
transform -1 0 315416 0 1 39652
box 0 496 2800 2224
use constant_block  constant_block_5
timestamp 1677077417
transform -1 0 205816 0 1 39652
box 0 496 2800 2224
use constant_block  constant_block_6
timestamp 1677077417
transform -1 0 151016 0 1 39652
box 0 496 2800 2224
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1677077417
transform 1 0 348400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1
timestamp 1677077417
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1677077417
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1677077417
transform -1 0 365800 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1677077417
transform -1 0 311000 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1677077417
transform -1 0 420600 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1677077417
transform -1 0 475400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1677077417
transform -1 0 530200 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__corner_pad  mgmt_corner\[0\]
timestamp 1677077417
transform -1 0 40000 0 -1 40800
box -271 -204 40000 40800
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1677077417
transform 0 1 676800 -1 0 40000
box -271 -204 40000 40800
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad
timestamp 1677077417
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad
timestamp 1677077417
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\]
timestamp 1677077417
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1677077417
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad
timestamp 1677077417
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclamp_pad
timestamp 1677077417
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\]
timestamp 1677077417
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1677077417
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1677077417
transform 0 1 675407 -1 0 116000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1677077417
transform 0 1 675407 -1 0 161200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1677077417
transform 0 1 675407 -1 0 206200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1677077417
transform 0 1 675407 -1 0 251400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1677077417
transform 0 1 675407 -1 0 296400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1677077417
transform 0 1 675407 -1 0 341400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1677077417
transform 0 1 675407 -1 0 386600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1677077417
transform 0 1 675407 -1 0 563800
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1677077417
transform 0 1 675407 -1 0 609000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1677077417
transform 0 1 675407 -1 0 654000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1677077417
transform 0 1 675407 -1 0 699200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1677077417
transform 0 1 675407 -1 0 744200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1677077417
transform 0 1 675407 -1 0 789200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1677077417
transform 0 1 675407 -1 0 878400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[14\]
timestamp 1677077417
transform 0 1 675407 -1 0 967600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[15\]
timestamp 1677077417
transform 1 0 626000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[16\]
timestamp 1677077417
transform 1 0 524200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[17\]
timestamp 1677077417
transform 1 0 472800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[18\]
timestamp 1677077417
transform 1 0 383800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1677077417
transform 1 0 282000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1677077417
transform 1 0 230400 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1677077417
transform 1 0 179000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1677077417
transform 1 0 127600 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1677077417
transform 1 0 76200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1677077417
transform 0 -1 42193 1 0 954200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1677077417
transform 0 -1 42193 1 0 784400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1677077417
transform 0 -1 42193 1 0 741200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1677077417
transform 0 -1 42193 1 0 698000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1677077417
transform 0 -1 42193 1 0 654800
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1677077417
transform 0 -1 42193 1 0 611600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1677077417
transform 0 -1 42193 1 0 568400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1677077417
transform 0 -1 42193 1 0 525200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[13\]
timestamp 1677077417
transform 0 -1 42193 1 0 397600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[14\]
timestamp 1677077417
transform 0 -1 42193 1 0 354400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[15\]
timestamp 1677077417
transform 0 -1 42193 1 0 311200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[16\]
timestamp 1677077417
transform 0 -1 42193 1 0 268000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[17\]
timestamp 1677077417
transform 0 -1 42193 1 0 224800
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[18\]
timestamp 1677077417
transform 0 -1 42193 1 0 181600
box -143 0 16134 42193
use sky130_fd_io__top_xres4v2  resetb_pad
timestamp 1677077417
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__corner_pad  user1_corner
timestamp 1677077417
transform 1 0 677600 0 1 996800
box -271 -204 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user1_vccd_lvclamp_pad
timestamp 1677077417
transform 0 1 678007 -1 0 922600
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1677077417
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1677077417
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1677077417
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1677077417
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user1_vssd_lvclamp_pad
timestamp 1677077417
transform 0 1 678007 -1 0 474800
box 0 -2177 17187 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1677077417
transform 0 -1 40800 1 0 997600
box -271 -204 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user2_vccd_lvclamp_pad
timestamp 1677077417
transform 0 -1 39593 1 0 912000
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1677077417
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1677077417
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user2_vssd_lvclamp_pad
timestamp 1677077417
transform 0 -1 39593 1 0 440800
box 0 -2177 17187 39593
<< labels >>
flabel metal2 s 675407 776611 675887 776667 0 FreeSans 400 0 0 0 mprj_analog_io[5]
port 3 nsew
flabel metal2 s 675407 779003 675887 779059 0 FreeSans 400 0 0 0 mprj_io_analog_en[12]
port 5 nsew
flabel metal2 s 675407 780291 675887 780347 0 FreeSans 400 0 0 0 mprj_io_analog_pol[12]
port 7 nsew
flabel metal2 s 675407 783327 675887 783383 0 FreeSans 400 0 0 0 mprj_io_analog_sel[12]
port 9 nsew
flabel metal2 s 675407 779647 675887 779703 0 FreeSans 400 0 0 0 mprj_io_dm[36]
port 11 nsew
flabel metal2 s 675407 777807 675887 777863 0 FreeSans 400 0 0 0 mprj_io_dm[37]
port 13 nsew
flabel metal2 s 675407 783971 675887 784027 0 FreeSans 400 0 0 0 mprj_io_dm[38]
port 15 nsew
flabel metal2 s 675407 784615 675887 784671 0 FreeSans 400 0 0 0 mprj_io_holdover[12]
port 17 nsew
flabel metal2 s 675407 787651 675887 787707 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[12]
port 19 nsew
flabel metal2 s 675407 780843 675887 780899 0 FreeSans 400 0 0 0 mprj_io_inp_dis[12]
port 21 nsew
flabel metal2 s 675407 788295 675887 788351 0 FreeSans 400 0 0 0 mprj_io_oeb[12]
port 23 nsew
flabel metal2 s 675407 785167 675887 785223 0 FreeSans 400 0 0 0 mprj_io_out[12]
port 25 nsew
flabel metal2 s 675407 775967 675887 776023 0 FreeSans 400 0 0 0 mprj_io_slow_sel[12]
port 27 nsew
flabel metal2 s 675407 787007 675887 787063 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[12]
port 29 nsew
flabel metal2 s 675407 774127 675887 774183 0 FreeSans 400 0 0 0 mprj_io_in[12]
port 31 nsew
flabel metal2 s 675407 865811 675887 865867 0 FreeSans 400 0 0 0 mprj_analog_io[6]
port 33 nsew
flabel metal2 s 675407 868203 675887 868259 0 FreeSans 400 0 0 0 mprj_io_analog_en[13]
port 35 nsew
flabel metal2 s 675407 869491 675887 869547 0 FreeSans 400 0 0 0 mprj_io_analog_pol[13]
port 37 nsew
flabel metal2 s 675407 872527 675887 872583 0 FreeSans 400 0 0 0 mprj_io_analog_sel[13]
port 39 nsew
flabel metal2 s 675407 868847 675887 868903 0 FreeSans 400 0 0 0 mprj_io_dm[39]
port 41 nsew
flabel metal2 s 675407 867007 675887 867063 0 FreeSans 400 0 0 0 mprj_io_dm[40]
port 43 nsew
flabel metal2 s 675407 873171 675887 873227 0 FreeSans 400 0 0 0 mprj_io_dm[41]
port 45 nsew
flabel metal2 s 675407 873815 675887 873871 0 FreeSans 400 0 0 0 mprj_io_holdover[13]
port 47 nsew
flabel metal2 s 675407 876851 675887 876907 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[13]
port 49 nsew
flabel metal2 s 675407 870043 675887 870099 0 FreeSans 400 0 0 0 mprj_io_inp_dis[13]
port 51 nsew
flabel metal2 s 675407 877495 675887 877551 0 FreeSans 400 0 0 0 mprj_io_oeb[13]
port 53 nsew
flabel metal2 s 675407 874367 675887 874423 0 FreeSans 400 0 0 0 mprj_io_out[13]
port 55 nsew
flabel metal2 s 675407 865167 675887 865223 0 FreeSans 400 0 0 0 mprj_io_slow_sel[13]
port 57 nsew
flabel metal2 s 675407 876207 675887 876263 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[13]
port 59 nsew
flabel metal2 s 675407 863327 675887 863383 0 FreeSans 400 0 0 0 mprj_io_in[13]
port 61 nsew
flabel metal2 s 675407 955011 675887 955067 0 FreeSans 400 0 0 0 mprj_analog_io[7]
port 63 nsew
flabel metal2 s 675407 957403 675887 957459 0 FreeSans 400 0 0 0 mprj_io_analog_en[14]
port 65 nsew
flabel metal2 s 675407 958691 675887 958747 0 FreeSans 400 0 0 0 mprj_io_analog_pol[14]
port 67 nsew
flabel metal2 s 675407 961727 675887 961783 0 FreeSans 400 0 0 0 mprj_io_analog_sel[14]
port 69 nsew
flabel metal2 s 675407 958047 675887 958103 0 FreeSans 400 0 0 0 mprj_io_dm[42]
port 71 nsew
flabel metal2 s 675407 956207 675887 956263 0 FreeSans 400 0 0 0 mprj_io_dm[43]
port 73 nsew
flabel metal2 s 675407 962371 675887 962427 0 FreeSans 400 0 0 0 mprj_io_dm[44]
port 75 nsew
flabel metal2 s 675407 963015 675887 963071 0 FreeSans 400 0 0 0 mprj_io_holdover[14]
port 77 nsew
flabel metal2 s 675407 966051 675887 966107 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[14]
port 79 nsew
flabel metal2 s 675407 959243 675887 959299 0 FreeSans 400 0 0 0 mprj_io_inp_dis[14]
port 81 nsew
flabel metal2 s 675407 966695 675887 966751 0 FreeSans 400 0 0 0 mprj_io_oeb[14]
port 83 nsew
flabel metal2 s 675407 963567 675887 963623 0 FreeSans 400 0 0 0 mprj_io_out[14]
port 85 nsew
flabel metal2 s 675407 954367 675887 954423 0 FreeSans 400 0 0 0 mprj_io_slow_sel[14]
port 87 nsew
flabel metal2 s 675407 965407 675887 965463 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[14]
port 89 nsew
flabel metal2 s 675407 952527 675887 952583 0 FreeSans 400 0 0 0 mprj_io_in[14]
port 91 nsew
flabel metal2 s 638533 995407 638589 995887 0 FreeSans 400 90 0 0 mprj_analog_io[8]
port 93 nsew
flabel metal2 s 636141 995407 636197 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[15]
port 95 nsew
flabel metal2 s 634853 995407 634909 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[15]
port 97 nsew
flabel metal2 s 631817 995407 631873 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[15]
port 99 nsew
flabel metal2 s 635497 995407 635553 995887 0 FreeSans 400 90 0 0 mprj_io_dm[45]
port 101 nsew
flabel metal2 s 637337 995407 637393 995887 0 FreeSans 400 90 0 0 mprj_io_dm[46]
port 103 nsew
flabel metal2 s 631173 995407 631229 995887 0 FreeSans 400 90 0 0 mprj_io_dm[47]
port 105 nsew
flabel metal2 s 630529 995407 630585 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[15]
port 107 nsew
flabel metal2 s 627493 995407 627549 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[15]
port 109 nsew
flabel metal2 s 634301 995407 634357 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[15]
port 111 nsew
flabel metal2 s 626849 995407 626905 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[15]
port 113 nsew
flabel metal2 s 629977 995407 630033 995887 0 FreeSans 400 90 0 0 mprj_io_out[15]
port 115 nsew
flabel metal2 s 639177 995407 639233 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[15]
port 117 nsew
flabel metal2 s 628137 995407 628193 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[15]
port 119 nsew
flabel metal2 s 641017 995407 641073 995887 0 FreeSans 400 90 0 0 mprj_io_in[15]
port 121 nsew
flabel metal2 s 536733 995407 536789 995887 0 FreeSans 400 90 0 0 mprj_analog_io[9]
port 123 nsew
flabel metal2 s 534341 995407 534397 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[16]
port 125 nsew
flabel metal2 s 533053 995407 533109 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[16]
port 127 nsew
flabel metal2 s 530017 995407 530073 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[16]
port 129 nsew
flabel metal2 s 533697 995407 533753 995887 0 FreeSans 400 90 0 0 mprj_io_dm[48]
port 131 nsew
flabel metal2 s 535537 995407 535593 995887 0 FreeSans 400 90 0 0 mprj_io_dm[49]
port 133 nsew
flabel metal2 s 529373 995407 529429 995887 0 FreeSans 400 90 0 0 mprj_io_dm[50]
port 135 nsew
flabel metal2 s 528729 995407 528785 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[16]
port 137 nsew
flabel metal2 s 525693 995407 525749 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[16]
port 139 nsew
flabel metal2 s 532501 995407 532557 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[16]
port 141 nsew
flabel metal2 s 525049 995407 525105 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[16]
port 143 nsew
flabel metal2 s 528177 995407 528233 995887 0 FreeSans 400 90 0 0 mprj_io_out[16]
port 145 nsew
flabel metal2 s 537377 995407 537433 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[16]
port 147 nsew
flabel metal2 s 526337 995407 526393 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[16]
port 149 nsew
flabel metal2 s 539217 995407 539273 995887 0 FreeSans 400 90 0 0 mprj_io_in[16]
port 151 nsew
flabel metal2 s 675407 775323 675887 775379 0 FreeSans 400 0 0 0 mprj_io_one[12]
port 153 nsew
flabel metal2 s 675407 864523 675887 864579 0 FreeSans 400 0 0 0 mprj_io_one[13]
port 155 nsew
flabel metal2 s 675407 953723 675887 953779 0 FreeSans 400 0 0 0 mprj_io_one[14]
port 157 nsew
flabel metal2 s 639821 995407 639877 995887 0 FreeSans 400 90 0 0 mprj_io_one[15]
port 159 nsew
flabel metal2 s 538021 995407 538077 995887 0 FreeSans 400 90 0 0 mprj_io_one[16]
port 161 nsew
flabel metal2 s 484137 995407 484193 995887 0 FreeSans 400 90 0 0 mprj_io_dm[52]
port 163 nsew
flabel metal2 s 477973 995407 478029 995887 0 FreeSans 400 90 0 0 mprj_io_dm[53]
port 165 nsew
flabel metal2 s 477329 995407 477385 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[17]
port 167 nsew
flabel metal2 s 474293 995407 474349 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[17]
port 169 nsew
flabel metal2 s 481101 995407 481157 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[17]
port 171 nsew
flabel metal2 s 473649 995407 473705 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[17]
port 173 nsew
flabel metal2 s 476777 995407 476833 995887 0 FreeSans 400 90 0 0 mprj_io_out[17]
port 175 nsew
flabel metal2 s 485977 995407 486033 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[17]
port 177 nsew
flabel metal2 s 474937 995407 474993 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[17]
port 179 nsew
flabel metal2 s 487817 995407 487873 995887 0 FreeSans 400 90 0 0 mprj_io_in[17]
port 181 nsew
flabel metal2 s 396333 995407 396389 995887 0 FreeSans 400 90 0 0 mprj_analog_io[11]
port 183 nsew
flabel metal2 s 393941 995407 393997 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[18]
port 185 nsew
flabel metal2 s 392653 995407 392709 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[18]
port 187 nsew
flabel metal2 s 389617 995407 389673 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[18]
port 189 nsew
flabel metal2 s 393297 995407 393353 995887 0 FreeSans 400 90 0 0 mprj_io_dm[54]
port 191 nsew
flabel metal2 s 395137 995407 395193 995887 0 FreeSans 400 90 0 0 mprj_io_dm[55]
port 193 nsew
flabel metal2 s 388973 995407 389029 995887 0 FreeSans 400 90 0 0 mprj_io_dm[56]
port 195 nsew
flabel metal2 s 388329 995407 388385 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[18]
port 197 nsew
flabel metal2 s 385293 995407 385349 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[18]
port 199 nsew
flabel metal2 s 392101 995407 392157 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[18]
port 201 nsew
flabel metal2 s 384649 995407 384705 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[18]
port 203 nsew
flabel metal2 s 387777 995407 387833 995887 0 FreeSans 400 90 0 0 mprj_io_out[18]
port 205 nsew
flabel metal2 s 396977 995407 397033 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[18]
port 207 nsew
flabel metal2 s 385937 995407 385993 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[18]
port 209 nsew
flabel metal2 s 398817 995407 398873 995887 0 FreeSans 400 90 0 0 mprj_io_in[18]
port 211 nsew
flabel metal2 s 485333 995407 485389 995887 0 FreeSans 400 90 0 0 mprj_analog_io[10]
port 213 nsew
flabel metal2 s 482941 995407 482997 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[17]
port 215 nsew
flabel metal2 s 481653 995407 481709 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[17]
port 217 nsew
flabel metal2 s 478617 995407 478673 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[17]
port 219 nsew
flabel metal2 s 482297 995407 482353 995887 0 FreeSans 400 90 0 0 mprj_io_dm[51]
port 221 nsew
flabel metal2 s 486621 995407 486677 995887 0 FreeSans 400 90 0 0 mprj_io_one[17]
port 223 nsew
flabel metal2 s 397621 995407 397677 995887 0 FreeSans 400 90 0 0 mprj_io_one[18]
port 225 nsew
flabel metal2 s 675407 739615 675887 739671 0 FreeSans 400 0 0 0 mprj_io_holdover[11]
port 227 nsew
flabel metal2 s 675407 742651 675887 742707 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[11]
port 229 nsew
flabel metal2 s 675407 735843 675887 735899 0 FreeSans 400 0 0 0 mprj_io_inp_dis[11]
port 231 nsew
flabel metal2 s 675407 743295 675887 743351 0 FreeSans 400 0 0 0 mprj_io_oeb[11]
port 233 nsew
flabel metal2 s 675407 740167 675887 740223 0 FreeSans 400 0 0 0 mprj_io_out[11]
port 235 nsew
flabel metal2 s 675407 730967 675887 731023 0 FreeSans 400 0 0 0 mprj_io_slow_sel[11]
port 237 nsew
flabel metal2 s 675407 742007 675887 742063 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[11]
port 239 nsew
flabel metal2 s 675407 729127 675887 729183 0 FreeSans 400 0 0 0 mprj_io_in[11]
port 241 nsew
flabel metal2 s 675407 686611 675887 686667 0 FreeSans 400 0 0 0 mprj_analog_io[3]
port 243 nsew
flabel metal2 s 675407 689003 675887 689059 0 FreeSans 400 0 0 0 mprj_io_analog_en[10]
port 245 nsew
flabel metal2 s 675407 690291 675887 690347 0 FreeSans 400 0 0 0 mprj_io_analog_pol[10]
port 247 nsew
flabel metal2 s 675407 693327 675887 693383 0 FreeSans 400 0 0 0 mprj_io_analog_sel[10]
port 249 nsew
flabel metal2 s 675407 689647 675887 689703 0 FreeSans 400 0 0 0 mprj_io_dm[30]
port 251 nsew
flabel metal2 s 675407 687807 675887 687863 0 FreeSans 400 0 0 0 mprj_io_dm[31]
port 253 nsew
flabel metal2 s 675407 693971 675887 694027 0 FreeSans 400 0 0 0 mprj_io_dm[32]
port 255 nsew
flabel metal2 s 675407 694615 675887 694671 0 FreeSans 400 0 0 0 mprj_io_holdover[10]
port 257 nsew
flabel metal2 s 675407 697651 675887 697707 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[10]
port 259 nsew
flabel metal2 s 675407 690843 675887 690899 0 FreeSans 400 0 0 0 mprj_io_inp_dis[10]
port 261 nsew
flabel metal2 s 675407 698295 675887 698351 0 FreeSans 400 0 0 0 mprj_io_oeb[10]
port 263 nsew
flabel metal2 s 675407 695167 675887 695223 0 FreeSans 400 0 0 0 mprj_io_out[10]
port 265 nsew
flabel metal2 s 675407 685967 675887 686023 0 FreeSans 400 0 0 0 mprj_io_slow_sel[10]
port 267 nsew
flabel metal2 s 675407 697007 675887 697063 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[10]
port 269 nsew
flabel metal2 s 675407 684127 675887 684183 0 FreeSans 400 0 0 0 mprj_io_in[10]
port 271 nsew
flabel metal2 s 675407 551211 675887 551267 0 FreeSans 400 0 0 0 mprj_analog_io[0]
port 273 nsew
flabel metal2 s 675407 553603 675887 553659 0 FreeSans 400 0 0 0 mprj_io_analog_en[7]
port 275 nsew
flabel metal2 s 675407 554891 675887 554947 0 FreeSans 400 0 0 0 mprj_io_analog_pol[7]
port 277 nsew
flabel metal2 s 675407 557927 675887 557983 0 FreeSans 400 0 0 0 mprj_io_analog_sel[7]
port 279 nsew
flabel metal2 s 675407 554247 675887 554303 0 FreeSans 400 0 0 0 mprj_io_dm[21]
port 281 nsew
flabel metal2 s 675407 552407 675887 552463 0 FreeSans 400 0 0 0 mprj_io_dm[22]
port 283 nsew
flabel metal2 s 675407 558571 675887 558627 0 FreeSans 400 0 0 0 mprj_io_dm[23]
port 285 nsew
flabel metal2 s 675407 559215 675887 559271 0 FreeSans 400 0 0 0 mprj_io_holdover[7]
port 287 nsew
flabel metal2 s 675407 562251 675887 562307 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[7]
port 289 nsew
flabel metal2 s 675407 555443 675887 555499 0 FreeSans 400 0 0 0 mprj_io_inp_dis[7]
port 291 nsew
flabel metal2 s 675407 562895 675887 562951 0 FreeSans 400 0 0 0 mprj_io_oeb[7]
port 293 nsew
flabel metal2 s 675407 559767 675887 559823 0 FreeSans 400 0 0 0 mprj_io_out[7]
port 295 nsew
flabel metal2 s 675407 550567 675887 550623 0 FreeSans 400 0 0 0 mprj_io_slow_sel[7]
port 297 nsew
flabel metal2 s 675407 561607 675887 561663 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[7]
port 299 nsew
flabel metal2 s 675407 548727 675887 548783 0 FreeSans 400 0 0 0 mprj_io_in[7]
port 301 nsew
flabel metal2 s 675407 596411 675887 596467 0 FreeSans 400 0 0 0 mprj_analog_io[1]
port 303 nsew
flabel metal2 s 675407 598803 675887 598859 0 FreeSans 400 0 0 0 mprj_io_analog_en[8]
port 305 nsew
flabel metal2 s 675407 600091 675887 600147 0 FreeSans 400 0 0 0 mprj_io_analog_pol[8]
port 307 nsew
flabel metal2 s 675407 603127 675887 603183 0 FreeSans 400 0 0 0 mprj_io_analog_sel[8]
port 309 nsew
flabel metal2 s 675407 599447 675887 599503 0 FreeSans 400 0 0 0 mprj_io_dm[24]
port 311 nsew
flabel metal2 s 675407 597607 675887 597663 0 FreeSans 400 0 0 0 mprj_io_dm[25]
port 313 nsew
flabel metal2 s 675407 603771 675887 603827 0 FreeSans 400 0 0 0 mprj_io_dm[26]
port 315 nsew
flabel metal2 s 675407 604415 675887 604471 0 FreeSans 400 0 0 0 mprj_io_holdover[8]
port 317 nsew
flabel metal2 s 675407 607451 675887 607507 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[8]
port 319 nsew
flabel metal2 s 675407 600643 675887 600699 0 FreeSans 400 0 0 0 mprj_io_inp_dis[8]
port 321 nsew
flabel metal2 s 675407 608095 675887 608151 0 FreeSans 400 0 0 0 mprj_io_oeb[8]
port 323 nsew
flabel metal2 s 675407 604967 675887 605023 0 FreeSans 400 0 0 0 mprj_io_out[8]
port 325 nsew
flabel metal2 s 675407 595767 675887 595823 0 FreeSans 400 0 0 0 mprj_io_slow_sel[8]
port 327 nsew
flabel metal2 s 675407 606807 675887 606863 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[8]
port 329 nsew
flabel metal2 s 675407 593927 675887 593983 0 FreeSans 400 0 0 0 mprj_io_in[8]
port 331 nsew
flabel metal2 s 675407 641411 675887 641467 0 FreeSans 400 0 0 0 mprj_analog_io[2]
port 333 nsew
flabel metal2 s 675407 643803 675887 643859 0 FreeSans 400 0 0 0 mprj_io_analog_en[9]
port 335 nsew
flabel metal2 s 675407 645091 675887 645147 0 FreeSans 400 0 0 0 mprj_io_analog_pol[9]
port 337 nsew
flabel metal2 s 675407 648127 675887 648183 0 FreeSans 400 0 0 0 mprj_io_analog_sel[9]
port 339 nsew
flabel metal2 s 675407 644447 675887 644503 0 FreeSans 400 0 0 0 mprj_io_dm[27]
port 341 nsew
flabel metal2 s 675407 642607 675887 642663 0 FreeSans 400 0 0 0 mprj_io_dm[28]
port 343 nsew
flabel metal2 s 675407 648771 675887 648827 0 FreeSans 400 0 0 0 mprj_io_dm[29]
port 345 nsew
flabel metal2 s 675407 649415 675887 649471 0 FreeSans 400 0 0 0 mprj_io_holdover[9]
port 347 nsew
flabel metal2 s 675407 652451 675887 652507 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[9]
port 349 nsew
flabel metal2 s 675407 645643 675887 645699 0 FreeSans 400 0 0 0 mprj_io_inp_dis[9]
port 351 nsew
flabel metal2 s 675407 653095 675887 653151 0 FreeSans 400 0 0 0 mprj_io_oeb[9]
port 353 nsew
flabel metal2 s 675407 649967 675887 650023 0 FreeSans 400 0 0 0 mprj_io_out[9]
port 355 nsew
flabel metal2 s 675407 640767 675887 640823 0 FreeSans 400 0 0 0 mprj_io_slow_sel[9]
port 357 nsew
flabel metal2 s 675407 651807 675887 651863 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[9]
port 359 nsew
flabel metal2 s 675407 638927 675887 638983 0 FreeSans 400 0 0 0 mprj_io_in[9]
port 361 nsew
flabel metal2 s 675407 549923 675887 549979 0 FreeSans 400 0 0 0 mprj_io_one[7]
port 363 nsew
flabel metal2 s 675407 595123 675887 595179 0 FreeSans 400 0 0 0 mprj_io_one[8]
port 365 nsew
flabel metal2 s 675407 640123 675887 640179 0 FreeSans 400 0 0 0 mprj_io_one[9]
port 367 nsew
flabel metal2 s 675407 685323 675887 685379 0 FreeSans 400 0 0 0 mprj_io_one[10]
port 369 nsew
flabel metal2 s 675407 730323 675887 730379 0 FreeSans 400 0 0 0 mprj_io_one[11]
port 371 nsew
flabel metal2 s 675407 731611 675887 731667 0 FreeSans 400 0 0 0 mprj_analog_io[4]
port 373 nsew
flabel metal2 s 675407 734003 675887 734059 0 FreeSans 400 0 0 0 mprj_io_analog_en[11]
port 375 nsew
flabel metal2 s 675407 735291 675887 735347 0 FreeSans 400 0 0 0 mprj_io_analog_pol[11]
port 377 nsew
flabel metal2 s 675407 738327 675887 738383 0 FreeSans 400 0 0 0 mprj_io_analog_sel[11]
port 379 nsew
flabel metal2 s 675407 734647 675887 734703 0 FreeSans 400 0 0 0 mprj_io_dm[33]
port 381 nsew
flabel metal2 s 675407 732807 675887 732863 0 FreeSans 400 0 0 0 mprj_io_dm[34]
port 383 nsew
flabel metal2 s 675407 738971 675887 739027 0 FreeSans 400 0 0 0 mprj_io_dm[35]
port 385 nsew
flabel metal2 s 295177 995407 295233 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[19]
port 387 nsew
flabel metal2 s 284137 995407 284193 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[19]
port 389 nsew
flabel metal2 s 297017 995407 297073 995887 0 FreeSans 400 90 0 0 mprj_io_in[19]
port 391 nsew
flabel metal2 s 242933 995407 242989 995887 0 FreeSans 400 90 0 0 mprj_analog_io[13]
port 393 nsew
flabel metal2 s 240541 995407 240597 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[20]
port 395 nsew
flabel metal2 s 239253 995407 239309 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[20]
port 397 nsew
flabel metal2 s 236217 995407 236273 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[20]
port 399 nsew
flabel metal2 s 239897 995407 239953 995887 0 FreeSans 400 90 0 0 mprj_io_dm[60]
port 401 nsew
flabel metal2 s 241737 995407 241793 995887 0 FreeSans 400 90 0 0 mprj_io_dm[61]
port 403 nsew
flabel metal2 s 235573 995407 235629 995887 0 FreeSans 400 90 0 0 mprj_io_dm[62]
port 405 nsew
flabel metal2 s 234929 995407 234985 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[20]
port 407 nsew
flabel metal2 s 231893 995407 231949 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[20]
port 409 nsew
flabel metal2 s 238701 995407 238757 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[20]
port 411 nsew
flabel metal2 s 231249 995407 231305 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[20]
port 413 nsew
flabel metal2 s 234377 995407 234433 995887 0 FreeSans 400 90 0 0 mprj_io_out[20]
port 415 nsew
flabel metal2 s 243577 995407 243633 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[20]
port 417 nsew
flabel metal2 s 232537 995407 232593 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[20]
port 419 nsew
flabel metal2 s 245417 995407 245473 995887 0 FreeSans 400 90 0 0 mprj_io_in[20]
port 421 nsew
flabel metal2 s 294533 995407 294589 995887 0 FreeSans 400 90 0 0 mprj_analog_io[12]
port 423 nsew
flabel metal2 s 292141 995407 292197 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[19]
port 425 nsew
flabel metal2 s 290853 995407 290909 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[19]
port 427 nsew
flabel metal2 s 287817 995407 287873 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[19]
port 429 nsew
flabel metal2 s 291497 995407 291553 995887 0 FreeSans 400 90 0 0 mprj_io_dm[57]
port 431 nsew
flabel metal2 s 293337 995407 293393 995887 0 FreeSans 400 90 0 0 mprj_io_dm[58]
port 433 nsew
flabel metal2 s 287173 995407 287229 995887 0 FreeSans 400 90 0 0 mprj_io_dm[59]
port 435 nsew
flabel metal2 s 286529 995407 286585 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[19]
port 437 nsew
flabel metal2 s 283493 995407 283549 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[19]
port 439 nsew
flabel metal2 s 290301 995407 290357 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[19]
port 441 nsew
flabel metal2 s 282849 995407 282905 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[19]
port 443 nsew
flabel metal2 s 285977 995407 286033 995887 0 FreeSans 400 90 0 0 mprj_io_out[19]
port 445 nsew
flabel metal2 s 295821 995407 295877 995887 0 FreeSans 400 90 0 0 mprj_io_one[19]
port 447 nsew
flabel metal2 s 244221 995407 244277 995887 0 FreeSans 400 90 0 0 mprj_io_one[20]
port 449 nsew
flabel metal2 s 194017 995407 194073 995887 0 FreeSans 400 90 0 0 mprj_io_in[21]
port 451 nsew
flabel metal2 s 140133 995407 140189 995887 0 FreeSans 400 90 0 0 mprj_analog_io[15]
port 453 nsew
flabel metal2 s 137741 995407 137797 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[22]
port 455 nsew
flabel metal2 s 136453 995407 136509 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[22]
port 457 nsew
flabel metal2 s 133417 995407 133473 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[22]
port 459 nsew
flabel metal2 s 137097 995407 137153 995887 0 FreeSans 400 90 0 0 mprj_io_dm[66]
port 461 nsew
flabel metal2 s 138937 995407 138993 995887 0 FreeSans 400 90 0 0 mprj_io_dm[67]
port 463 nsew
flabel metal2 s 132773 995407 132829 995887 0 FreeSans 400 90 0 0 mprj_io_dm[68]
port 465 nsew
flabel metal2 s 132129 995407 132185 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[22]
port 467 nsew
flabel metal2 s 129093 995407 129149 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[22]
port 469 nsew
flabel metal2 s 135901 995407 135957 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[22]
port 471 nsew
flabel metal2 s 128449 995407 128505 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[22]
port 473 nsew
flabel metal2 s 131577 995407 131633 995887 0 FreeSans 400 90 0 0 mprj_io_out[22]
port 475 nsew
flabel metal2 s 140777 995407 140833 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[22]
port 477 nsew
flabel metal2 s 129737 995407 129793 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[22]
port 479 nsew
flabel metal2 s 142617 995407 142673 995887 0 FreeSans 400 90 0 0 mprj_io_in[22]
port 481 nsew
flabel metal2 s 88733 995407 88789 995887 0 FreeSans 400 90 0 0 mprj_analog_io[16]
port 483 nsew
flabel metal2 s 86341 995407 86397 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[23]
port 485 nsew
flabel metal2 s 85053 995407 85109 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[23]
port 487 nsew
flabel metal2 s 82017 995407 82073 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[23]
port 489 nsew
flabel metal2 s 85697 995407 85753 995887 0 FreeSans 400 90 0 0 mprj_io_dm[69]
port 491 nsew
flabel metal2 s 87537 995407 87593 995887 0 FreeSans 400 90 0 0 mprj_io_dm[70]
port 493 nsew
flabel metal2 s 81373 995407 81429 995887 0 FreeSans 400 90 0 0 mprj_io_dm[71]
port 495 nsew
flabel metal2 s 80729 995407 80785 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[23]
port 497 nsew
flabel metal2 s 77693 995407 77749 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[23]
port 499 nsew
flabel metal2 s 84501 995407 84557 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[23]
port 501 nsew
flabel metal2 s 77049 995407 77105 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[23]
port 503 nsew
flabel metal2 s 80177 995407 80233 995887 0 FreeSans 400 90 0 0 mprj_io_out[23]
port 505 nsew
flabel metal2 s 89377 995407 89433 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[23]
port 507 nsew
flabel metal2 s 78337 995407 78393 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[23]
port 509 nsew
flabel metal2 s 91217 995407 91273 995887 0 FreeSans 400 90 0 0 mprj_io_in[23]
port 511 nsew
flabel metal2 s 41713 966733 42193 966789 0 FreeSans 400 0 0 0 mprj_analog_io[17]
port 513 nsew
flabel metal2 s 41713 964341 42193 964397 0 FreeSans 400 0 0 0 mprj_io_analog_en[24]
port 515 nsew
flabel metal2 s 41713 963053 42193 963109 0 FreeSans 400 0 0 0 mprj_io_analog_pol[24]
port 517 nsew
flabel metal2 s 41713 960017 42193 960073 0 FreeSans 400 0 0 0 mprj_io_analog_sel[24]
port 519 nsew
flabel metal2 s 41713 963697 42193 963753 0 FreeSans 400 0 0 0 mprj_io_dm[72]
port 521 nsew
flabel metal2 s 41713 965537 42193 965593 0 FreeSans 400 0 0 0 mprj_io_dm[73]
port 523 nsew
flabel metal2 s 41713 959373 42193 959429 0 FreeSans 400 0 0 0 mprj_io_dm[74]
port 525 nsew
flabel metal2 s 41713 958729 42193 958785 0 FreeSans 400 0 0 0 mprj_io_holdover[24]
port 527 nsew
flabel metal2 s 41713 955693 42193 955749 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[24]
port 529 nsew
flabel metal2 s 41713 962501 42193 962557 0 FreeSans 400 0 0 0 mprj_io_inp_dis[24]
port 531 nsew
flabel metal2 s 41713 955049 42193 955105 0 FreeSans 400 0 0 0 mprj_io_oeb[24]
port 533 nsew
flabel metal2 s 41713 958177 42193 958233 0 FreeSans 400 0 0 0 mprj_io_out[24]
port 535 nsew
flabel metal2 s 41713 967377 42193 967433 0 FreeSans 400 0 0 0 mprj_io_slow_sel[24]
port 537 nsew
flabel metal2 s 41713 956337 42193 956393 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[24]
port 539 nsew
flabel metal2 s 41713 969217 42193 969273 0 FreeSans 400 0 0 0 mprj_io_in[24]
port 541 nsew
flabel metal2 s 41713 796933 42193 796989 0 FreeSans 400 0 0 0 mprj_analog_io[18]
port 543 nsew
flabel metal2 s 41713 794541 42193 794597 0 FreeSans 400 0 0 0 mprj_io_analog_en[25]
port 545 nsew
flabel metal2 s 41713 793253 42193 793309 0 FreeSans 400 0 0 0 mprj_io_analog_pol[25]
port 547 nsew
flabel metal2 s 41713 790217 42193 790273 0 FreeSans 400 0 0 0 mprj_io_analog_sel[25]
port 549 nsew
flabel metal2 s 41713 793897 42193 793953 0 FreeSans 400 0 0 0 mprj_io_dm[75]
port 551 nsew
flabel metal2 s 41713 795737 42193 795793 0 FreeSans 400 0 0 0 mprj_io_dm[76]
port 553 nsew
flabel metal2 s 41713 789573 42193 789629 0 FreeSans 400 0 0 0 mprj_io_dm[77]
port 555 nsew
flabel metal2 s 41713 788929 42193 788985 0 FreeSans 400 0 0 0 mprj_io_holdover[25]
port 557 nsew
flabel metal2 s 41713 785893 42193 785949 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[25]
port 559 nsew
flabel metal2 s 41713 792701 42193 792757 0 FreeSans 400 0 0 0 mprj_io_inp_dis[25]
port 561 nsew
flabel metal2 s 41713 785249 42193 785305 0 FreeSans 400 0 0 0 mprj_io_oeb[25]
port 563 nsew
flabel metal2 s 41713 788377 42193 788433 0 FreeSans 400 0 0 0 mprj_io_out[25]
port 565 nsew
flabel metal2 s 41713 797577 42193 797633 0 FreeSans 400 0 0 0 mprj_io_slow_sel[25]
port 567 nsew
flabel metal2 s 41713 786537 42193 786593 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[25]
port 569 nsew
flabel metal2 s 41713 799417 42193 799473 0 FreeSans 400 0 0 0 mprj_io_in[25]
port 571 nsew
flabel metal2 s 191533 995407 191589 995887 0 FreeSans 400 90 0 0 mprj_analog_io[14]
port 573 nsew
flabel metal2 s 189141 995407 189197 995887 0 FreeSans 400 90 0 0 mprj_io_analog_en[21]
port 575 nsew
flabel metal2 s 187853 995407 187909 995887 0 FreeSans 400 90 0 0 mprj_io_analog_pol[21]
port 577 nsew
flabel metal2 s 184817 995407 184873 995887 0 FreeSans 400 90 0 0 mprj_io_analog_sel[21]
port 579 nsew
flabel metal2 s 188497 995407 188553 995887 0 FreeSans 400 90 0 0 mprj_io_dm[63]
port 581 nsew
flabel metal2 s 190337 995407 190393 995887 0 FreeSans 400 90 0 0 mprj_io_dm[64]
port 583 nsew
flabel metal2 s 184173 995407 184229 995887 0 FreeSans 400 90 0 0 mprj_io_dm[65]
port 585 nsew
flabel metal2 s 183529 995407 183585 995887 0 FreeSans 400 90 0 0 mprj_io_holdover[21]
port 587 nsew
flabel metal2 s 180493 995407 180549 995887 0 FreeSans 400 90 0 0 mprj_io_ib_mode_sel[21]
port 589 nsew
flabel metal2 s 187301 995407 187357 995887 0 FreeSans 400 90 0 0 mprj_io_inp_dis[21]
port 591 nsew
flabel metal2 s 179849 995407 179905 995887 0 FreeSans 400 90 0 0 mprj_io_oeb[21]
port 593 nsew
flabel metal2 s 182977 995407 183033 995887 0 FreeSans 400 90 0 0 mprj_io_out[21]
port 595 nsew
flabel metal2 s 192177 995407 192233 995887 0 FreeSans 400 90 0 0 mprj_io_slow_sel[21]
port 597 nsew
flabel metal2 s 181137 995407 181193 995887 0 FreeSans 400 90 0 0 mprj_io_vtrip_sel[21]
port 599 nsew
flabel metal2 s 192821 995407 192877 995887 0 FreeSans 400 90 0 0 mprj_io_one[21]
port 601 nsew
flabel metal2 s 141421 995407 141477 995887 0 FreeSans 400 90 0 0 mprj_io_one[22]
port 603 nsew
flabel metal2 s 90021 995407 90077 995887 0 FreeSans 400 90 0 0 mprj_io_one[23]
port 605 nsew
flabel metal2 s 41713 968021 42193 968077 0 FreeSans 400 0 0 0 mprj_io_one[24]
port 607 nsew
flabel metal2 s 41713 798221 42193 798277 0 FreeSans 400 0 0 0 mprj_io_one[25]
port 609 nsew
flabel metal2 s 41713 577897 42193 577953 0 FreeSans 400 0 0 0 mprj_io_dm[90]
port 611 nsew
flabel metal2 s 41713 579737 42193 579793 0 FreeSans 400 0 0 0 mprj_io_dm[91]
port 613 nsew
flabel metal2 s 41713 573573 42193 573629 0 FreeSans 400 0 0 0 mprj_io_dm[92]
port 615 nsew
flabel metal2 s 41713 572929 42193 572985 0 FreeSans 400 0 0 0 mprj_io_holdover[30]
port 617 nsew
flabel metal2 s 41713 569893 42193 569949 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[30]
port 619 nsew
flabel metal2 s 41713 576701 42193 576757 0 FreeSans 400 0 0 0 mprj_io_inp_dis[30]
port 621 nsew
flabel metal2 s 41713 569249 42193 569305 0 FreeSans 400 0 0 0 mprj_io_oeb[30]
port 623 nsew
flabel metal2 s 41713 572377 42193 572433 0 FreeSans 400 0 0 0 mprj_io_out[30]
port 625 nsew
flabel metal2 s 41713 581577 42193 581633 0 FreeSans 400 0 0 0 mprj_io_slow_sel[30]
port 627 nsew
flabel metal2 s 41713 570537 42193 570593 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[30]
port 629 nsew
flabel metal2 s 41713 583417 42193 583473 0 FreeSans 400 0 0 0 mprj_io_in[30]
port 631 nsew
flabel metal2 s 41713 537733 42193 537789 0 FreeSans 400 0 0 0 mprj_analog_io[24]
port 633 nsew
flabel metal2 s 41713 535341 42193 535397 0 FreeSans 400 0 0 0 mprj_io_analog_en[31]
port 635 nsew
flabel metal2 s 41713 534053 42193 534109 0 FreeSans 400 0 0 0 mprj_io_analog_pol[31]
port 637 nsew
flabel metal2 s 41713 531017 42193 531073 0 FreeSans 400 0 0 0 mprj_io_analog_sel[31]
port 639 nsew
flabel metal2 s 41713 534697 42193 534753 0 FreeSans 400 0 0 0 mprj_io_dm[93]
port 641 nsew
flabel metal2 s 41713 536537 42193 536593 0 FreeSans 400 0 0 0 mprj_io_dm[94]
port 643 nsew
flabel metal2 s 41713 530373 42193 530429 0 FreeSans 400 0 0 0 mprj_io_dm[95]
port 645 nsew
flabel metal2 s 41713 529729 42193 529785 0 FreeSans 400 0 0 0 mprj_io_holdover[31]
port 647 nsew
flabel metal2 s 41713 526693 42193 526749 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[31]
port 649 nsew
flabel metal2 s 41713 533501 42193 533557 0 FreeSans 400 0 0 0 mprj_io_inp_dis[31]
port 651 nsew
flabel metal2 s 41713 526049 42193 526105 0 FreeSans 400 0 0 0 mprj_io_oeb[31]
port 653 nsew
flabel metal2 s 41713 529177 42193 529233 0 FreeSans 400 0 0 0 mprj_io_out[31]
port 655 nsew
flabel metal2 s 41713 538377 42193 538433 0 FreeSans 400 0 0 0 mprj_io_slow_sel[31]
port 657 nsew
flabel metal2 s 41713 527337 42193 527393 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[31]
port 659 nsew
flabel metal2 s 41713 540217 42193 540273 0 FreeSans 400 0 0 0 mprj_io_in[31]
port 661 nsew
flabel metal2 s 41713 753733 42193 753789 0 FreeSans 400 0 0 0 mprj_analog_io[19]
port 663 nsew
flabel metal2 s 41713 751341 42193 751397 0 FreeSans 400 0 0 0 mprj_io_analog_en[26]
port 665 nsew
flabel metal2 s 41713 750053 42193 750109 0 FreeSans 400 0 0 0 mprj_io_analog_pol[26]
port 667 nsew
flabel metal2 s 41713 747017 42193 747073 0 FreeSans 400 0 0 0 mprj_io_analog_sel[26]
port 669 nsew
flabel metal2 s 41713 750697 42193 750753 0 FreeSans 400 0 0 0 mprj_io_dm[78]
port 671 nsew
flabel metal2 s 41713 752537 42193 752593 0 FreeSans 400 0 0 0 mprj_io_dm[79]
port 673 nsew
flabel metal2 s 41713 746373 42193 746429 0 FreeSans 400 0 0 0 mprj_io_dm[80]
port 675 nsew
flabel metal2 s 41713 745729 42193 745785 0 FreeSans 400 0 0 0 mprj_io_holdover[26]
port 677 nsew
flabel metal2 s 41713 742693 42193 742749 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[26]
port 679 nsew
flabel metal2 s 41713 749501 42193 749557 0 FreeSans 400 0 0 0 mprj_io_inp_dis[26]
port 681 nsew
flabel metal2 s 41713 742049 42193 742105 0 FreeSans 400 0 0 0 mprj_io_oeb[26]
port 683 nsew
flabel metal2 s 41713 745177 42193 745233 0 FreeSans 400 0 0 0 mprj_io_out[26]
port 685 nsew
flabel metal2 s 41713 754377 42193 754433 0 FreeSans 400 0 0 0 mprj_io_slow_sel[26]
port 687 nsew
flabel metal2 s 41713 743337 42193 743393 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[26]
port 689 nsew
flabel metal2 s 41713 756217 42193 756273 0 FreeSans 400 0 0 0 mprj_io_in[26]
port 691 nsew
flabel metal2 s 41713 710533 42193 710589 0 FreeSans 400 0 0 0 mprj_analog_io[20]
port 693 nsew
flabel metal2 s 41713 708141 42193 708197 0 FreeSans 400 0 0 0 mprj_io_analog_en[27]
port 695 nsew
flabel metal2 s 41713 706853 42193 706909 0 FreeSans 400 0 0 0 mprj_io_analog_pol[27]
port 697 nsew
flabel metal2 s 41713 703817 42193 703873 0 FreeSans 400 0 0 0 mprj_io_analog_sel[27]
port 699 nsew
flabel metal2 s 41713 707497 42193 707553 0 FreeSans 400 0 0 0 mprj_io_dm[81]
port 701 nsew
flabel metal2 s 41713 709337 42193 709393 0 FreeSans 400 0 0 0 mprj_io_dm[82]
port 703 nsew
flabel metal2 s 41713 703173 42193 703229 0 FreeSans 400 0 0 0 mprj_io_dm[83]
port 705 nsew
flabel metal2 s 41713 702529 42193 702585 0 FreeSans 400 0 0 0 mprj_io_holdover[27]
port 707 nsew
flabel metal2 s 41713 699493 42193 699549 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[27]
port 709 nsew
flabel metal2 s 41713 706301 42193 706357 0 FreeSans 400 0 0 0 mprj_io_inp_dis[27]
port 711 nsew
flabel metal2 s 41713 698849 42193 698905 0 FreeSans 400 0 0 0 mprj_io_oeb[27]
port 713 nsew
flabel metal2 s 41713 701977 42193 702033 0 FreeSans 400 0 0 0 mprj_io_out[27]
port 715 nsew
flabel metal2 s 41713 711177 42193 711233 0 FreeSans 400 0 0 0 mprj_io_slow_sel[27]
port 717 nsew
flabel metal2 s 41713 700137 42193 700193 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[27]
port 719 nsew
flabel metal2 s 41713 713017 42193 713073 0 FreeSans 400 0 0 0 mprj_io_in[27]
port 721 nsew
flabel metal2 s 41713 667333 42193 667389 0 FreeSans 400 0 0 0 mprj_analog_io[21]
port 723 nsew
flabel metal2 s 41713 664941 42193 664997 0 FreeSans 400 0 0 0 mprj_io_analog_en[28]
port 725 nsew
flabel metal2 s 41713 663653 42193 663709 0 FreeSans 400 0 0 0 mprj_io_analog_pol[28]
port 727 nsew
flabel metal2 s 41713 660617 42193 660673 0 FreeSans 400 0 0 0 mprj_io_analog_sel[28]
port 729 nsew
flabel metal2 s 41713 664297 42193 664353 0 FreeSans 400 0 0 0 mprj_io_dm[84]
port 731 nsew
flabel metal2 s 41713 666137 42193 666193 0 FreeSans 400 0 0 0 mprj_io_dm[85]
port 733 nsew
flabel metal2 s 41713 659973 42193 660029 0 FreeSans 400 0 0 0 mprj_io_dm[86]
port 735 nsew
flabel metal2 s 41713 659329 42193 659385 0 FreeSans 400 0 0 0 mprj_io_holdover[28]
port 737 nsew
flabel metal2 s 41713 656293 42193 656349 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[28]
port 739 nsew
flabel metal2 s 41713 663101 42193 663157 0 FreeSans 400 0 0 0 mprj_io_inp_dis[28]
port 741 nsew
flabel metal2 s 41713 655649 42193 655705 0 FreeSans 400 0 0 0 mprj_io_oeb[28]
port 743 nsew
flabel metal2 s 41713 658777 42193 658833 0 FreeSans 400 0 0 0 mprj_io_out[28]
port 745 nsew
flabel metal2 s 41713 667977 42193 668033 0 FreeSans 400 0 0 0 mprj_io_slow_sel[28]
port 747 nsew
flabel metal2 s 41713 656937 42193 656993 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[28]
port 749 nsew
flabel metal2 s 41713 669817 42193 669873 0 FreeSans 400 0 0 0 mprj_io_in[28]
port 751 nsew
flabel metal2 s 41713 624133 42193 624189 0 FreeSans 400 0 0 0 mprj_analog_io[22]
port 753 nsew
flabel metal2 s 41713 621741 42193 621797 0 FreeSans 400 0 0 0 mprj_io_analog_en[29]
port 755 nsew
flabel metal2 s 41713 620453 42193 620509 0 FreeSans 400 0 0 0 mprj_io_analog_pol[29]
port 757 nsew
flabel metal2 s 41713 617417 42193 617473 0 FreeSans 400 0 0 0 mprj_io_analog_sel[29]
port 759 nsew
flabel metal2 s 41713 621097 42193 621153 0 FreeSans 400 0 0 0 mprj_io_dm[87]
port 761 nsew
flabel metal2 s 41713 622937 42193 622993 0 FreeSans 400 0 0 0 mprj_io_dm[88]
port 763 nsew
flabel metal2 s 41713 616773 42193 616829 0 FreeSans 400 0 0 0 mprj_io_dm[89]
port 765 nsew
flabel metal2 s 41713 616129 42193 616185 0 FreeSans 400 0 0 0 mprj_io_holdover[29]
port 767 nsew
flabel metal2 s 41713 613093 42193 613149 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[29]
port 769 nsew
flabel metal2 s 41713 619901 42193 619957 0 FreeSans 400 0 0 0 mprj_io_inp_dis[29]
port 771 nsew
flabel metal2 s 41713 612449 42193 612505 0 FreeSans 400 0 0 0 mprj_io_oeb[29]
port 773 nsew
flabel metal2 s 41713 615577 42193 615633 0 FreeSans 400 0 0 0 mprj_io_out[29]
port 775 nsew
flabel metal2 s 41713 624777 42193 624833 0 FreeSans 400 0 0 0 mprj_io_slow_sel[29]
port 777 nsew
flabel metal2 s 41713 613737 42193 613793 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[29]
port 779 nsew
flabel metal2 s 41713 626617 42193 626673 0 FreeSans 400 0 0 0 mprj_io_in[29]
port 781 nsew
flabel metal2 s 41713 580933 42193 580989 0 FreeSans 400 0 0 0 mprj_analog_io[23]
port 783 nsew
flabel metal2 s 41713 578541 42193 578597 0 FreeSans 400 0 0 0 mprj_io_analog_en[30]
port 785 nsew
flabel metal2 s 41713 577253 42193 577309 0 FreeSans 400 0 0 0 mprj_io_analog_pol[30]
port 787 nsew
flabel metal2 s 41713 574217 42193 574273 0 FreeSans 400 0 0 0 mprj_io_analog_sel[30]
port 789 nsew
flabel metal2 s 41713 755021 42193 755077 0 FreeSans 400 0 0 0 mprj_io_one[26]
port 791 nsew
flabel metal2 s 41713 711821 42193 711877 0 FreeSans 400 0 0 0 mprj_io_one[27]
port 793 nsew
flabel metal2 s 41713 668621 42193 668677 0 FreeSans 400 0 0 0 mprj_io_one[28]
port 795 nsew
flabel metal2 s 41713 625421 42193 625477 0 FreeSans 400 0 0 0 mprj_io_one[29]
port 797 nsew
flabel metal2 s 41713 582221 42193 582277 0 FreeSans 400 0 0 0 mprj_io_one[30]
port 799 nsew
flabel metal2 s 41713 539021 42193 539077 0 FreeSans 400 0 0 0 mprj_io_one[31]
port 801 nsew
flabel metal2 s 41713 236137 42193 236193 0 FreeSans 400 0 0 0 mprj_io_dm[109]
port 803 nsew
flabel metal2 s 41713 229973 42193 230029 0 FreeSans 400 0 0 0 mprj_io_dm[110]
port 805 nsew
flabel metal2 s 41713 229329 42193 229385 0 FreeSans 400 0 0 0 mprj_io_holdover[36]
port 807 nsew
flabel metal2 s 41713 226293 42193 226349 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[36]
port 809 nsew
flabel metal2 s 41713 233101 42193 233157 0 FreeSans 400 0 0 0 mprj_io_inp_dis[36]
port 811 nsew
flabel metal2 s 41713 225649 42193 225705 0 FreeSans 400 0 0 0 mprj_io_oeb[36]
port 813 nsew
flabel metal2 s 41713 228777 42193 228833 0 FreeSans 400 0 0 0 mprj_io_out[36]
port 815 nsew
flabel metal2 s 41713 237977 42193 238033 0 FreeSans 400 0 0 0 mprj_io_slow_sel[36]
port 817 nsew
flabel metal2 s 41713 226937 42193 226993 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[36]
port 819 nsew
flabel metal2 s 41713 239817 42193 239873 0 FreeSans 400 0 0 0 mprj_io_in[36]
port 821 nsew
flabel metal2 s 41713 191741 42193 191797 0 FreeSans 400 0 0 0 mprj_io_analog_en[37]
port 823 nsew
flabel metal2 s 41713 190453 42193 190509 0 FreeSans 400 0 0 0 mprj_io_analog_pol[37]
port 825 nsew
flabel metal2 s 41713 187417 42193 187473 0 FreeSans 400 0 0 0 mprj_io_analog_sel[37]
port 827 nsew
flabel metal2 s 41713 191097 42193 191153 0 FreeSans 400 0 0 0 mprj_io_dm[111]
port 829 nsew
flabel metal2 s 41713 192937 42193 192993 0 FreeSans 400 0 0 0 mprj_io_dm[112]
port 831 nsew
flabel metal2 s 41713 186773 42193 186829 0 FreeSans 400 0 0 0 mprj_io_dm[113]
port 833 nsew
flabel metal2 s 41713 186129 42193 186185 0 FreeSans 400 0 0 0 mprj_io_holdover[37]
port 835 nsew
flabel metal2 s 41713 183093 42193 183149 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[37]
port 837 nsew
flabel metal2 s 41713 189901 42193 189957 0 FreeSans 400 0 0 0 mprj_io_inp_dis[37]
port 839 nsew
flabel metal2 s 41713 182449 42193 182505 0 FreeSans 400 0 0 0 mprj_io_oeb[37]
port 841 nsew
flabel metal2 s 41713 185577 42193 185633 0 FreeSans 400 0 0 0 mprj_io_out[37]
port 843 nsew
flabel metal2 s 41713 194777 42193 194833 0 FreeSans 400 0 0 0 mprj_io_slow_sel[37]
port 845 nsew
flabel metal2 s 41713 183737 42193 183793 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[37]
port 847 nsew
flabel metal2 s 41713 196617 42193 196673 0 FreeSans 400 0 0 0 mprj_io_in[37]
port 849 nsew
flabel metal2 s 187327 41713 187383 42193 0 FreeSans 400 90 0 0 clock_core
port 851 nsew
flabel metal2 s 194043 41713 194099 42193 0 FreeSans 400 90 0 0 por
port 853 nsew
flabel metal2 s 306967 41713 307023 42193 0 FreeSans 400 90 0 0 flash_csb_core
port 855 nsew
flabel metal2 s 310095 41713 310151 42193 0 FreeSans 400 90 0 0 flash_csb_oeb_core
port 857 nsew
flabel metal2 s 41713 410133 42193 410189 0 FreeSans 400 0 0 0 mprj_analog_io[25]
port 859 nsew
flabel metal2 s 41713 407741 42193 407797 0 FreeSans 400 0 0 0 mprj_io_analog_en[32]
port 861 nsew
flabel metal2 s 41713 406453 42193 406509 0 FreeSans 400 0 0 0 mprj_io_analog_pol[32]
port 863 nsew
flabel metal2 s 41713 403417 42193 403473 0 FreeSans 400 0 0 0 mprj_io_analog_sel[32]
port 865 nsew
flabel metal2 s 41713 407097 42193 407153 0 FreeSans 400 0 0 0 mprj_io_dm[96]
port 867 nsew
flabel metal2 s 41713 408937 42193 408993 0 FreeSans 400 0 0 0 mprj_io_dm[97]
port 869 nsew
flabel metal2 s 41713 402773 42193 402829 0 FreeSans 400 0 0 0 mprj_io_dm[98]
port 871 nsew
flabel metal2 s 41713 402129 42193 402185 0 FreeSans 400 0 0 0 mprj_io_holdover[32]
port 873 nsew
flabel metal2 s 41713 399093 42193 399149 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[32]
port 875 nsew
flabel metal2 s 41713 405901 42193 405957 0 FreeSans 400 0 0 0 mprj_io_inp_dis[32]
port 877 nsew
flabel metal2 s 41713 398449 42193 398505 0 FreeSans 400 0 0 0 mprj_io_oeb[32]
port 879 nsew
flabel metal2 s 41713 401577 42193 401633 0 FreeSans 400 0 0 0 mprj_io_out[32]
port 881 nsew
flabel metal2 s 41713 410777 42193 410833 0 FreeSans 400 0 0 0 mprj_io_slow_sel[32]
port 883 nsew
flabel metal2 s 41713 399737 42193 399793 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[32]
port 885 nsew
flabel metal2 s 41713 412617 42193 412673 0 FreeSans 400 0 0 0 mprj_io_in[32]
port 887 nsew
flabel metal2 s 41713 366933 42193 366989 0 FreeSans 400 0 0 0 mprj_analog_io[26]
port 889 nsew
flabel metal2 s 41713 364541 42193 364597 0 FreeSans 400 0 0 0 mprj_io_analog_en[33]
port 891 nsew
flabel metal2 s 41713 363253 42193 363309 0 FreeSans 400 0 0 0 mprj_io_analog_pol[33]
port 893 nsew
flabel metal2 s 41713 360217 42193 360273 0 FreeSans 400 0 0 0 mprj_io_analog_sel[33]
port 895 nsew
flabel metal2 s 41713 365737 42193 365793 0 FreeSans 400 0 0 0 mprj_io_dm[100]
port 897 nsew
flabel metal2 s 41713 359573 42193 359629 0 FreeSans 400 0 0 0 mprj_io_dm[101]
port 899 nsew
flabel metal2 s 41713 363897 42193 363953 0 FreeSans 400 0 0 0 mprj_io_dm[99]
port 901 nsew
flabel metal2 s 41713 358929 42193 358985 0 FreeSans 400 0 0 0 mprj_io_holdover[33]
port 903 nsew
flabel metal2 s 41713 355893 42193 355949 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[33]
port 905 nsew
flabel metal2 s 41713 362701 42193 362757 0 FreeSans 400 0 0 0 mprj_io_inp_dis[33]
port 907 nsew
flabel metal2 s 41713 355249 42193 355305 0 FreeSans 400 0 0 0 mprj_io_oeb[33]
port 909 nsew
flabel metal2 s 41713 358377 42193 358433 0 FreeSans 400 0 0 0 mprj_io_out[33]
port 911 nsew
flabel metal2 s 41713 367577 42193 367633 0 FreeSans 400 0 0 0 mprj_io_slow_sel[33]
port 913 nsew
flabel metal2 s 41713 356537 42193 356593 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[33]
port 915 nsew
flabel metal2 s 41713 369417 42193 369473 0 FreeSans 400 0 0 0 mprj_io_in[33]
port 917 nsew
flabel metal2 s 41713 323733 42193 323789 0 FreeSans 400 0 0 0 mprj_analog_io[27]
port 919 nsew
flabel metal2 s 41713 321341 42193 321397 0 FreeSans 400 0 0 0 mprj_io_analog_en[34]
port 921 nsew
flabel metal2 s 41713 320053 42193 320109 0 FreeSans 400 0 0 0 mprj_io_analog_pol[34]
port 923 nsew
flabel metal2 s 41713 317017 42193 317073 0 FreeSans 400 0 0 0 mprj_io_analog_sel[34]
port 925 nsew
flabel metal2 s 41713 320697 42193 320753 0 FreeSans 400 0 0 0 mprj_io_dm[102]
port 927 nsew
flabel metal2 s 41713 322537 42193 322593 0 FreeSans 400 0 0 0 mprj_io_dm[103]
port 929 nsew
flabel metal2 s 41713 316373 42193 316429 0 FreeSans 400 0 0 0 mprj_io_dm[104]
port 931 nsew
flabel metal2 s 41713 315729 42193 315785 0 FreeSans 400 0 0 0 mprj_io_holdover[34]
port 933 nsew
flabel metal2 s 41713 312693 42193 312749 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[34]
port 935 nsew
flabel metal2 s 141667 39934 141813 40000 0 FreeSans 400 0 0 0 resetb_core_h
port 937 nsew
flabel metal2 s 41713 319501 42193 319557 0 FreeSans 400 0 0 0 mprj_io_inp_dis[34]
port 939 nsew
flabel metal2 s 41713 312049 42193 312105 0 FreeSans 400 0 0 0 mprj_io_oeb[34]
port 941 nsew
flabel metal2 s 41713 315177 42193 315233 0 FreeSans 400 0 0 0 mprj_io_out[34]
port 943 nsew
flabel metal2 s 41713 324377 42193 324433 0 FreeSans 400 0 0 0 mprj_io_slow_sel[34]
port 945 nsew
flabel metal2 s 41713 313337 42193 313393 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[34]
port 947 nsew
flabel metal2 s 41713 326217 42193 326273 0 FreeSans 400 0 0 0 mprj_io_in[34]
port 949 nsew
flabel metal2 s 41713 280533 42193 280589 0 FreeSans 400 0 0 0 mprj_analog_io[28]
port 951 nsew
flabel metal2 s 41713 278141 42193 278197 0 FreeSans 400 0 0 0 mprj_io_analog_en[35]
port 953 nsew
flabel metal2 s 41713 276853 42193 276909 0 FreeSans 400 0 0 0 mprj_io_analog_pol[35]
port 955 nsew
flabel metal2 s 41713 273817 42193 273873 0 FreeSans 400 0 0 0 mprj_io_analog_sel[35]
port 957 nsew
flabel metal2 s 41713 277497 42193 277553 0 FreeSans 400 0 0 0 mprj_io_dm[105]
port 959 nsew
flabel metal2 s 41713 279337 42193 279393 0 FreeSans 400 0 0 0 mprj_io_dm[106]
port 961 nsew
flabel metal2 s 41713 273173 42193 273229 0 FreeSans 400 0 0 0 mprj_io_dm[107]
port 963 nsew
flabel metal2 s 41713 272529 42193 272585 0 FreeSans 400 0 0 0 mprj_io_holdover[35]
port 965 nsew
flabel metal2 s 41713 269493 42193 269549 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[35]
port 967 nsew
flabel metal2 s 41713 276301 42193 276357 0 FreeSans 400 0 0 0 mprj_io_inp_dis[35]
port 969 nsew
flabel metal2 s 41713 268849 42193 268905 0 FreeSans 400 0 0 0 mprj_io_oeb[35]
port 971 nsew
flabel metal2 s 41713 271977 42193 272033 0 FreeSans 400 0 0 0 mprj_io_out[35]
port 973 nsew
flabel metal2 s 41713 281177 42193 281233 0 FreeSans 400 0 0 0 mprj_io_slow_sel[35]
port 975 nsew
flabel metal2 s 41713 270137 42193 270193 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[35]
port 977 nsew
flabel metal2 s 41713 283017 42193 283073 0 FreeSans 400 0 0 0 mprj_io_in[35]
port 979 nsew
flabel metal2 s 41713 234941 42193 234997 0 FreeSans 400 0 0 0 mprj_io_analog_en[36]
port 981 nsew
flabel metal2 s 41713 233653 42193 233709 0 FreeSans 400 0 0 0 mprj_io_analog_pol[36]
port 983 nsew
flabel metal2 s 41713 230617 42193 230673 0 FreeSans 400 0 0 0 mprj_io_analog_sel[36]
port 985 nsew
flabel metal2 s 41713 234297 42193 234353 0 FreeSans 400 0 0 0 mprj_io_dm[108]
port 987 nsew
flabel metal2 s 41713 411421 42193 411477 0 FreeSans 400 0 0 0 mprj_io_one[32]
port 989 nsew
flabel metal2 s 41713 368221 42193 368277 0 FreeSans 400 0 0 0 mprj_io_one[33]
port 991 nsew
flabel metal2 s 41713 325021 42193 325077 0 FreeSans 400 0 0 0 mprj_io_one[34]
port 993 nsew
flabel metal2 s 41713 281821 42193 281877 0 FreeSans 400 0 0 0 mprj_io_one[35]
port 995 nsew
flabel metal2 s 41713 238621 42193 238677 0 FreeSans 400 0 0 0 mprj_io_one[36]
port 997 nsew
flabel metal2 s 41713 195421 42193 195477 0 FreeSans 400 0 0 0 mprj_io_one[37]
port 999 nsew
flabel metal2 s 308255 41713 308311 42193 0 FreeSans 400 90 0 0 porb_h
port 1001 nsew
flabel metal2 s 675407 286203 675887 286259 0 FreeSans 400 0 0 0 mprj_io_analog_en[4]
port 1003 nsew
flabel metal2 s 675407 287491 675887 287547 0 FreeSans 400 0 0 0 mprj_io_analog_pol[4]
port 1005 nsew
flabel metal2 s 675407 290527 675887 290583 0 FreeSans 400 0 0 0 mprj_io_analog_sel[4]
port 1007 nsew
flabel metal2 s 675407 286847 675887 286903 0 FreeSans 400 0 0 0 mprj_io_dm[12]
port 1009 nsew
flabel metal2 s 675407 285007 675887 285063 0 FreeSans 400 0 0 0 mprj_io_dm[13]
port 1011 nsew
flabel metal2 s 675407 291171 675887 291227 0 FreeSans 400 0 0 0 mprj_io_dm[14]
port 1013 nsew
flabel metal2 s 675407 291815 675887 291871 0 FreeSans 400 0 0 0 mprj_io_holdover[4]
port 1015 nsew
flabel metal2 s 675407 294851 675887 294907 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[4]
port 1017 nsew
flabel metal2 s 675407 288043 675887 288099 0 FreeSans 400 0 0 0 mprj_io_inp_dis[4]
port 1019 nsew
flabel metal2 s 675407 295495 675887 295551 0 FreeSans 400 0 0 0 mprj_io_oeb[4]
port 1021 nsew
flabel metal2 s 675407 292367 675887 292423 0 FreeSans 400 0 0 0 mprj_io_out[4]
port 1023 nsew
flabel metal2 s 675407 283167 675887 283223 0 FreeSans 400 0 0 0 mprj_io_slow_sel[4]
port 1025 nsew
flabel metal2 s 675407 294207 675887 294263 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[4]
port 1027 nsew
flabel metal2 s 675407 281327 675887 281383 0 FreeSans 400 0 0 0 mprj_io_in[4]
port 1029 nsew
flabel metal2 s 675407 331203 675887 331259 0 FreeSans 400 0 0 0 mprj_io_analog_en[5]
port 1031 nsew
flabel metal2 s 675407 332491 675887 332547 0 FreeSans 400 0 0 0 mprj_io_analog_pol[5]
port 1033 nsew
flabel metal2 s 675407 335527 675887 335583 0 FreeSans 400 0 0 0 mprj_io_analog_sel[5]
port 1035 nsew
flabel metal2 s 675407 331847 675887 331903 0 FreeSans 400 0 0 0 mprj_io_dm[15]
port 1037 nsew
flabel metal2 s 675407 330007 675887 330063 0 FreeSans 400 0 0 0 mprj_io_dm[16]
port 1039 nsew
flabel metal2 s 675407 336171 675887 336227 0 FreeSans 400 0 0 0 mprj_io_dm[17]
port 1041 nsew
flabel metal2 s 675407 336815 675887 336871 0 FreeSans 400 0 0 0 mprj_io_holdover[5]
port 1043 nsew
flabel metal2 s 675407 339851 675887 339907 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[5]
port 1045 nsew
flabel metal2 s 675407 333043 675887 333099 0 FreeSans 400 0 0 0 mprj_io_inp_dis[5]
port 1047 nsew
flabel metal2 s 675407 340495 675887 340551 0 FreeSans 400 0 0 0 mprj_io_oeb[5]
port 1049 nsew
flabel metal2 s 675407 337367 675887 337423 0 FreeSans 400 0 0 0 mprj_io_out[5]
port 1051 nsew
flabel metal2 s 675407 328167 675887 328223 0 FreeSans 400 0 0 0 mprj_io_slow_sel[5]
port 1053 nsew
flabel metal2 s 675407 339207 675887 339263 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[5]
port 1055 nsew
flabel metal2 s 675407 326327 675887 326383 0 FreeSans 400 0 0 0 mprj_io_in[5]
port 1057 nsew
flabel metal2 s 675407 376403 675887 376459 0 FreeSans 400 0 0 0 mprj_io_analog_en[6]
port 1059 nsew
flabel metal2 s 675407 282523 675887 282579 0 FreeSans 400 0 0 0 mprj_io_one[4]
port 1061 nsew
flabel metal2 s 675407 327523 675887 327579 0 FreeSans 400 0 0 0 mprj_io_one[5]
port 1063 nsew
flabel metal2 s 675407 372723 675887 372779 0 FreeSans 400 0 0 0 mprj_io_one[6]
port 1065 nsew
flabel metal2 s 675407 377691 675887 377747 0 FreeSans 400 0 0 0 mprj_io_analog_pol[6]
port 1067 nsew
flabel metal2 s 675407 380727 675887 380783 0 FreeSans 400 0 0 0 mprj_io_analog_sel[6]
port 1069 nsew
flabel metal2 s 675407 377047 675887 377103 0 FreeSans 400 0 0 0 mprj_io_dm[18]
port 1071 nsew
flabel metal2 s 675407 375207 675887 375263 0 FreeSans 400 0 0 0 mprj_io_dm[19]
port 1073 nsew
flabel metal2 s 675407 381371 675887 381427 0 FreeSans 400 0 0 0 mprj_io_dm[20]
port 1075 nsew
flabel metal2 s 675407 382015 675887 382071 0 FreeSans 400 0 0 0 mprj_io_holdover[6]
port 1077 nsew
flabel metal2 s 675407 385051 675887 385107 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[6]
port 1079 nsew
flabel metal2 s 675407 378243 675887 378299 0 FreeSans 400 0 0 0 mprj_io_inp_dis[6]
port 1081 nsew
flabel metal2 s 675407 385695 675887 385751 0 FreeSans 400 0 0 0 mprj_io_oeb[6]
port 1083 nsew
flabel metal2 s 675407 382567 675887 382623 0 FreeSans 400 0 0 0 mprj_io_out[6]
port 1085 nsew
flabel metal2 s 675407 373367 675887 373423 0 FreeSans 400 0 0 0 mprj_io_slow_sel[6]
port 1087 nsew
flabel metal2 s 675407 384407 675887 384463 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[6]
port 1089 nsew
flabel metal2 s 675407 371527 675887 371583 0 FreeSans 400 0 0 0 mprj_io_in[6]
port 1091 nsew
flabel metal2 s 471367 41713 471423 42193 0 FreeSans 400 90 0 0 flash_io1_do_core
port 1093 nsew
flabel metal2 s 467043 41713 467099 42193 0 FreeSans 400 90 0 0 flash_io1_ieb_core
port 1095 nsew
flabel metal2 s 474495 41713 474551 42193 0 FreeSans 400 90 0 0 flash_io1_oeb_core
port 1097 nsew
flabel metal2 s 515127 41713 515183 42193 0 FreeSans 400 90 0 0 gpio_in_core
port 1099 nsew
flabel metal2 s 412243 41713 412299 42193 0 FreeSans 400 90 0 0 flash_io0_ieb_core
port 1101 nsew
flabel metal2 s 419695 41713 419751 42193 0 FreeSans 400 90 0 0 flash_io0_oeb_core
port 1103 nsew
flabel metal2 s 460327 41713 460383 42193 0 FreeSans 400 90 0 0 flash_io1_di_core
port 1105 nsew
flabel metal2 s 361767 41713 361823 42193 0 FreeSans 400 90 0 0 flash_clk_core
port 1107 nsew
flabel metal2 s 364895 41713 364951 42193 0 FreeSans 400 90 0 0 flash_clk_oeb_core
port 1109 nsew
flabel metal2 s 405527 41713 405583 42193 0 FreeSans 400 90 0 0 flash_io0_di_core
port 1111 nsew
flabel metal2 s 416567 41713 416623 42193 0 FreeSans 400 90 0 0 flash_io0_do_core
port 1113 nsew
flabel metal2 s 526167 41713 526223 42193 0 FreeSans 400 90 0 0 gpio_out_core
port 1115 nsew
flabel metal2 s 675407 151003 675887 151059 0 FreeSans 400 0 0 0 mprj_io_analog_en[1]
port 1117 nsew
flabel metal2 s 675407 152291 675887 152347 0 FreeSans 400 0 0 0 mprj_io_analog_pol[1]
port 1119 nsew
flabel metal2 s 675407 155327 675887 155383 0 FreeSans 400 0 0 0 mprj_io_analog_sel[1]
port 1121 nsew
flabel metal2 s 675407 151647 675887 151703 0 FreeSans 400 0 0 0 mprj_io_dm[3]
port 1123 nsew
flabel metal2 s 675407 149807 675887 149863 0 FreeSans 400 0 0 0 mprj_io_dm[4]
port 1125 nsew
flabel metal2 s 675407 155971 675887 156027 0 FreeSans 400 0 0 0 mprj_io_dm[5]
port 1127 nsew
flabel metal2 s 675407 156615 675887 156671 0 FreeSans 400 0 0 0 mprj_io_holdover[1]
port 1129 nsew
flabel metal2 s 675407 159651 675887 159707 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[1]
port 1131 nsew
flabel metal2 s 675407 152843 675887 152899 0 FreeSans 400 0 0 0 mprj_io_inp_dis[1]
port 1133 nsew
flabel metal2 s 675407 160295 675887 160351 0 FreeSans 400 0 0 0 mprj_io_oeb[1]
port 1135 nsew
flabel metal2 s 675407 157167 675887 157223 0 FreeSans 400 0 0 0 mprj_io_out[1]
port 1137 nsew
flabel metal2 s 675407 147967 675887 148023 0 FreeSans 400 0 0 0 mprj_io_slow_sel[1]
port 1139 nsew
flabel metal2 s 675407 159007 675887 159063 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[1]
port 1141 nsew
flabel metal2 s 675407 146127 675887 146183 0 FreeSans 400 0 0 0 mprj_io_in[1]
port 1143 nsew
flabel metal2 s 675407 196003 675887 196059 0 FreeSans 400 0 0 0 mprj_io_analog_en[2]
port 1145 nsew
flabel metal2 s 675407 197291 675887 197347 0 FreeSans 400 0 0 0 mprj_io_analog_pol[2]
port 1147 nsew
flabel metal2 s 675407 200327 675887 200383 0 FreeSans 400 0 0 0 mprj_io_analog_sel[2]
port 1149 nsew
flabel metal2 s 675407 196647 675887 196703 0 FreeSans 400 0 0 0 mprj_io_dm[6]
port 1151 nsew
flabel metal2 s 675407 194807 675887 194863 0 FreeSans 400 0 0 0 mprj_io_dm[7]
port 1153 nsew
flabel metal2 s 675407 200971 675887 201027 0 FreeSans 400 0 0 0 mprj_io_dm[8]
port 1155 nsew
flabel metal2 s 675407 201615 675887 201671 0 FreeSans 400 0 0 0 mprj_io_holdover[2]
port 1157 nsew
flabel metal2 s 675407 204651 675887 204707 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[2]
port 1159 nsew
flabel metal2 s 675407 197843 675887 197899 0 FreeSans 400 0 0 0 mprj_io_inp_dis[2]
port 1161 nsew
flabel metal2 s 675407 205295 675887 205351 0 FreeSans 400 0 0 0 mprj_io_oeb[2]
port 1163 nsew
flabel metal2 s 675407 202167 675887 202223 0 FreeSans 400 0 0 0 mprj_io_out[2]
port 1165 nsew
flabel metal2 s 675407 102123 675887 102179 0 FreeSans 400 0 0 0 mprj_io_one[0]
port 1167 nsew
flabel metal2 s 675407 147323 675887 147379 0 FreeSans 400 0 0 0 mprj_io_one[1]
port 1169 nsew
flabel metal2 s 675407 192323 675887 192379 0 FreeSans 400 0 0 0 mprj_io_one[2]
port 1171 nsew
flabel metal2 s 675407 237523 675887 237579 0 FreeSans 400 0 0 0 mprj_io_one[3]
port 1173 nsew
flabel metal2 s 675407 192967 675887 193023 0 FreeSans 400 0 0 0 mprj_io_slow_sel[2]
port 1175 nsew
flabel metal2 s 675407 204007 675887 204063 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[2]
port 1177 nsew
flabel metal2 s 675407 191127 675887 191183 0 FreeSans 400 0 0 0 mprj_io_in[2]
port 1179 nsew
flabel metal2 s 675407 241203 675887 241259 0 FreeSans 400 0 0 0 mprj_io_analog_en[3]
port 1181 nsew
flabel metal2 s 675407 242491 675887 242547 0 FreeSans 400 0 0 0 mprj_io_analog_pol[3]
port 1183 nsew
flabel metal2 s 675407 245527 675887 245583 0 FreeSans 400 0 0 0 mprj_io_analog_sel[3]
port 1185 nsew
flabel metal2 s 675407 240007 675887 240063 0 FreeSans 400 0 0 0 mprj_io_dm[10]
port 1187 nsew
flabel metal2 s 675407 246171 675887 246227 0 FreeSans 400 0 0 0 mprj_io_dm[11]
port 1189 nsew
flabel metal2 s 675407 241847 675887 241903 0 FreeSans 400 0 0 0 mprj_io_dm[9]
port 1191 nsew
flabel metal2 s 675407 246815 675887 246871 0 FreeSans 400 0 0 0 mprj_io_holdover[3]
port 1193 nsew
flabel metal2 s 675407 249851 675887 249907 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[3]
port 1195 nsew
flabel metal2 s 675407 243043 675887 243099 0 FreeSans 400 0 0 0 mprj_io_inp_dis[3]
port 1197 nsew
flabel metal2 s 675407 250495 675887 250551 0 FreeSans 400 0 0 0 mprj_io_oeb[3]
port 1199 nsew
flabel metal2 s 675407 247367 675887 247423 0 FreeSans 400 0 0 0 mprj_io_out[3]
port 1201 nsew
flabel metal2 s 675407 238167 675887 238223 0 FreeSans 400 0 0 0 mprj_io_slow_sel[3]
port 1203 nsew
flabel metal2 s 675407 249207 675887 249263 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[3]
port 1205 nsew
flabel metal2 s 529295 41713 529351 42193 0 FreeSans 400 90 0 0 gpio_outenb_core
port 1207 nsew
flabel metal2 s 675407 105803 675887 105859 0 FreeSans 400 0 0 0 mprj_io_analog_en[0]
port 1209 nsew
flabel metal2 s 675407 107091 675887 107147 0 FreeSans 400 0 0 0 mprj_io_analog_pol[0]
port 1211 nsew
flabel metal2 s 675407 110127 675887 110183 0 FreeSans 400 0 0 0 mprj_io_analog_sel[0]
port 1213 nsew
flabel metal2 s 675407 106447 675887 106503 0 FreeSans 400 0 0 0 mprj_io_dm[0]
port 1215 nsew
flabel metal2 s 675407 104607 675887 104663 0 FreeSans 400 0 0 0 mprj_io_dm[1]
port 1217 nsew
flabel metal2 s 675407 110771 675887 110827 0 FreeSans 400 0 0 0 mprj_io_dm[2]
port 1219 nsew
flabel metal2 s 675407 111415 675887 111471 0 FreeSans 400 0 0 0 mprj_io_holdover[0]
port 1221 nsew
flabel metal2 s 675407 114451 675887 114507 0 FreeSans 400 0 0 0 mprj_io_ib_mode_sel[0]
port 1223 nsew
flabel metal2 s 675407 107643 675887 107699 0 FreeSans 400 0 0 0 mprj_io_inp_dis[0]
port 1225 nsew
flabel metal2 s 675407 115095 675887 115151 0 FreeSans 400 0 0 0 mprj_io_oeb[0]
port 1227 nsew
flabel metal2 s 675407 111967 675887 112023 0 FreeSans 400 0 0 0 mprj_io_out[0]
port 1229 nsew
flabel metal2 s 675407 102767 675887 102823 0 FreeSans 400 0 0 0 mprj_io_slow_sel[0]
port 1231 nsew
flabel metal2 s 675407 113807 675887 113863 0 FreeSans 400 0 0 0 mprj_io_vtrip_sel[0]
port 1233 nsew
flabel metal2 s 675407 100927 675887 100983 0 FreeSans 400 0 0 0 mprj_io_in[0]
port 1235 nsew
flabel metal2 s 675407 236327 675887 236383 0 FreeSans 400 0 0 0 mprj_io_in[3]
port 1237 nsew
flabel metal2 s 521843 41713 521899 42193 0 FreeSans 400 90 0 0 gpio_inenb_core
port 1239 nsew
flabel metal2 s 520647 41713 520703 42193 0 FreeSans 400 90 0 0 gpio_mode0_core
port 1241 nsew
flabel metal2 s 524971 41713 525027 42193 0 FreeSans 400 90 0 0 gpio_mode1_core
port 1243 nsew
rlabel metal1 s 142538 40100 142538 40100 4 xres_vss_loop
flabel metal4 s 132600 36323 132792 37013 6 FreeSans 400 0 0 0 vdda
port 1246 nsew
flabel metal4 s 36323 455607 37013 455799 6 FreeSans 400 0 0 0 vdda2
port 1248 nsew
flabel metal4 s 28653 440800 28719 455800 6 FreeSans 400 0 0 0 vssa2
port 1250 nsew
flabel metal4 s 38503 455546 39593 455800 0 FreeSans 400 0 0 0 vccd
port 1252 nsew
flabel metal4 s 680587 459800 681277 459993 0 FreeSans 400 0 0 0 vdda1
port 1254 nsew
flabel metal4 s 32933 455546 33623 455800 0 FreeSans 400 0 0 0 vddio
port 1256 nsew
flabel metal4 s 132600 28653 147600 28719 0 FreeSans 400 0 0 0 vssa
port 1258 nsew
flabel metal4 s 688881 459800 688947 474800 0 FreeSans 400 0 0 0 vssa1
port 1260 nsew
flabel metal4 s 132600 30753 132854 31683 0 FreeSans 400 0 0 0 vssd
port 1262 nsew
flabel metal4 s 0 455645 4843 456094 0 FreeSans 400 0 0 0 vssio
port 1264 nsew
flabel metal5 s 187640 6598 200180 19088 6 FreeSans 400 0 0 0 clock
port 1267 nsew
flabel metal5 s 351040 6598 363580 19088 6 FreeSans 400 0 0 0 flash_clk
port 1269 nsew
flabel metal5 s 296240 6598 308780 19088 6 FreeSans 400 0 0 0 flash_csb
port 1271 nsew
flabel metal5 s 405840 6598 418380 19088 6 FreeSans 400 0 0 0 flash_io0
port 1273 nsew
flabel metal5 s 460640 6598 473180 19088 6 FreeSans 400 0 0 0 flash_io1
port 1275 nsew
flabel metal5 s 515440 6598 527980 19088 6 FreeSans 400 0 0 0 gpio
port 1277 nsew
flabel metal5 s 6167 70054 19619 80934 6 FreeSans 400 0 0 0 vccd_pad
port 1279 nsew
flabel metal5 s 624222 6811 636390 18975 6 FreeSans 400 0 0 0 vdda_pad
port 1281 nsew
flabel metal5 s 6811 111610 18975 123778 6 FreeSans 400 0 0 0 vddio_pad
port 1283 nsew
flabel metal5 s 6811 871210 18975 883378 6 FreeSans 400 0 0 0 vddio_pad2
port 1285 nsew
flabel metal5 s 80222 6811 92390 18975 6 FreeSans 400 0 0 0 vssa_pad
port 1287 nsew
flabel metal5 s 243266 6167 254146 19619 6 FreeSans 400 0 0 0 vssd_pad
port 1289 nsew
flabel metal5 s 570422 6811 582590 18975 6 FreeSans 400 0 0 0 vssio_pad
port 1291 nsew
flabel metal5 s 334810 1018624 346978 1030788 6 FreeSans 400 0 0 0 vssio_pad2
port 1293 nsew
flabel metal5 s 698512 101240 711002 113780 6 FreeSans 400 0 0 0 mprj_io[0]
port 1295 nsew
flabel metal5 s 698512 684440 711002 696980 6 FreeSans 400 0 0 0 mprj_io[10]
port 1297 nsew
flabel metal5 s 698512 729440 711002 741980 6 FreeSans 400 0 0 0 mprj_io[11]
port 1299 nsew
flabel metal5 s 698512 774440 711002 786980 6 FreeSans 400 0 0 0 mprj_io[12]
port 1301 nsew
flabel metal5 s 698512 863640 711002 876180 6 FreeSans 400 0 0 0 mprj_io[13]
port 1303 nsew
flabel metal5 s 698512 952840 711002 965380 6 FreeSans 400 0 0 0 mprj_io[14]
port 1305 nsew
flabel metal5 s 628220 1018512 640760 1031002 6 FreeSans 400 0 0 0 mprj_io[15]
port 1307 nsew
flabel metal5 s 526420 1018512 538960 1031002 6 FreeSans 400 0 0 0 mprj_io[16]
port 1309 nsew
flabel metal5 s 475020 1018512 487560 1031002 6 FreeSans 400 0 0 0 mprj_io[17]
port 1311 nsew
flabel metal5 s 386020 1018512 398560 1031002 6 FreeSans 400 0 0 0 mprj_io[18]
port 1313 nsew
flabel metal5 s 698512 146440 711002 158980 6 FreeSans 400 0 0 0 mprj_io[1]
port 1315 nsew
flabel metal5 s 698512 191440 711002 203980 6 FreeSans 400 0 0 0 mprj_io[2]
port 1317 nsew
flabel metal5 s 698512 236640 711002 249180 6 FreeSans 400 0 0 0 mprj_io[3]
port 1319 nsew
flabel metal5 s 698512 281640 711002 294180 6 FreeSans 400 0 0 0 mprj_io[4]
port 1321 nsew
flabel metal5 s 698512 326640 711002 339180 6 FreeSans 400 0 0 0 mprj_io[5]
port 1323 nsew
flabel metal5 s 698512 371840 711002 384380 6 FreeSans 400 0 0 0 mprj_io[6]
port 1325 nsew
flabel metal5 s 698512 549040 711002 561580 6 FreeSans 400 0 0 0 mprj_io[7]
port 1327 nsew
flabel metal5 s 698512 594240 711002 606780 6 FreeSans 400 0 0 0 mprj_io[8]
port 1329 nsew
flabel metal5 s 698512 639240 711002 651780 6 FreeSans 400 0 0 0 mprj_io[9]
port 1331 nsew
flabel metal5 s 284220 1018512 296760 1031002 6 FreeSans 400 0 0 0 mprj_io[19]
port 1333 nsew
flabel metal5 s 6598 613820 19088 626360 6 FreeSans 400 0 0 0 mprj_io[29]
port 1335 nsew
flabel metal5 s 6598 570620 19088 583160 6 FreeSans 400 0 0 0 mprj_io[30]
port 1337 nsew
flabel metal5 s 6598 527420 19088 539960 6 FreeSans 400 0 0 0 mprj_io[31]
port 1339 nsew
flabel metal5 s 6598 399820 19088 412360 6 FreeSans 400 0 0 0 mprj_io[32]
port 1341 nsew
flabel metal5 s 6598 356620 19088 369160 6 FreeSans 400 0 0 0 mprj_io[33]
port 1343 nsew
flabel metal5 s 6598 313420 19088 325960 6 FreeSans 400 0 0 0 mprj_io[34]
port 1345 nsew
flabel metal5 s 6598 270220 19088 282760 6 FreeSans 400 0 0 0 mprj_io[35]
port 1347 nsew
flabel metal5 s 6598 227020 19088 239560 6 FreeSans 400 0 0 0 mprj_io[36]
port 1349 nsew
flabel metal5 s 6598 183820 19088 196360 6 FreeSans 400 0 0 0 mprj_io[37]
port 1351 nsew
flabel metal5 s 232620 1018512 245160 1031002 6 FreeSans 400 0 0 0 mprj_io[20]
port 1353 nsew
flabel metal5 s 181220 1018512 193760 1031002 6 FreeSans 400 0 0 0 mprj_io[21]
port 1355 nsew
flabel metal5 s 129820 1018512 142360 1031002 6 FreeSans 400 0 0 0 mprj_io[22]
port 1357 nsew
flabel metal5 s 78420 1018512 90960 1031002 6 FreeSans 400 0 0 0 mprj_io[23]
port 1359 nsew
flabel metal5 s 6598 956420 19088 968960 6 FreeSans 400 0 0 0 mprj_io[24]
port 1361 nsew
flabel metal5 s 6598 786620 19088 799160 6 FreeSans 400 0 0 0 mprj_io[25]
port 1363 nsew
flabel metal5 s 6598 743420 19088 755960 6 FreeSans 400 0 0 0 mprj_io[26]
port 1365 nsew
flabel metal5 s 6598 700220 19088 712760 6 FreeSans 400 0 0 0 mprj_io[27]
port 1367 nsew
flabel metal5 s 6598 657020 19088 669560 6 FreeSans 400 0 0 0 mprj_io[28]
port 1369 nsew
flabel metal5 s 136713 7143 144149 18309 6 FreeSans 400 0 0 0 resetb
port 1371 nsew
flabel metal5 s 697980 909666 711432 920546 6 FreeSans 400 0 0 0 vccd1_pad
port 1373 nsew
flabel metal5 s 698624 819822 710788 831990 6 FreeSans 400 0 0 0 vdda1_pad
port 1375 nsew
flabel metal5 s 698624 505222 710788 517390 6 FreeSans 400 0 0 0 vdda1_pad2
port 1377 nsew
flabel metal5 s 577010 1018624 589178 1030788 6 FreeSans 400 0 0 0 vssa1_pad
port 1379 nsew
flabel metal5 s 698624 417022 710788 429190 6 FreeSans 400 0 0 0 vssa1_pad2
port 1381 nsew
flabel metal5 s 697980 461866 711432 472746 6 FreeSans 400 0 0 0 vssd1_pad
port 1383 nsew
flabel metal5 s 6167 914054 19619 924934 6 FreeSans 400 0 0 0 vccd2_pad
port 1385 nsew
flabel metal5 s 6811 484410 18975 496578 6 FreeSans 400 0 0 0 vdda2_pad
port 1387 nsew
flabel metal5 s 6811 829010 18975 841178 6 FreeSans 400 0 0 0 vssa2_pad
port 1389 nsew
flabel metal5 s 6167 442854 19619 453734 6 FreeSans 400 0 0 0 vssd2_pad
port 1391 nsew
rlabel metal3 s 140494 40183 140494 40183 4 xresloop
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
