VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO housekeeping_alt
  CLASS BLOCK ;
  FOREIGN housekeeping_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END housekeeping_alt
END LIBRARY

