VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect
  CLASS BLOCK ;
  FOREIGN mgmt_protect ;
  ORIGIN 0.000 0.000 ;
  SIZE 2120.000 BY 160.000 ;
  PIN caravel_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 -2.000 979.710 4.000 ;
    END
  END caravel_clk
  PIN caravel_clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 41.520 2122.000 42.120 ;
    END
  END caravel_clk2
  PIN caravel_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 -2.000 982.930 4.000 ;
    END
  END caravel_rstn
  PIN la_data_in_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 156.000 484.750 162.000 ;
    END
  END la_data_in_core[0]
  PIN la_data_in_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.470 156.000 1726.750 162.000 ;
    END
  END la_data_in_core[100]
  PIN la_data_in_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 156.000 1739.170 162.000 ;
    END
  END la_data_in_core[101]
  PIN la_data_in_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.310 156.000 1751.590 162.000 ;
    END
  END la_data_in_core[102]
  PIN la_data_in_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.730 156.000 1764.010 162.000 ;
    END
  END la_data_in_core[103]
  PIN la_data_in_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.150 156.000 1776.430 162.000 ;
    END
  END la_data_in_core[104]
  PIN la_data_in_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1788.570 156.000 1788.850 162.000 ;
    END
  END la_data_in_core[105]
  PIN la_data_in_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.990 156.000 1801.270 162.000 ;
    END
  END la_data_in_core[106]
  PIN la_data_in_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.410 156.000 1813.690 162.000 ;
    END
  END la_data_in_core[107]
  PIN la_data_in_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 156.000 1826.110 162.000 ;
    END
  END la_data_in_core[108]
  PIN la_data_in_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.250 156.000 1838.530 162.000 ;
    END
  END la_data_in_core[109]
  PIN la_data_in_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 156.000 608.950 162.000 ;
    END
  END la_data_in_core[10]
  PIN la_data_in_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.670 156.000 1850.950 162.000 ;
    END
  END la_data_in_core[110]
  PIN la_data_in_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.090 156.000 1863.370 162.000 ;
    END
  END la_data_in_core[111]
  PIN la_data_in_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.510 156.000 1875.790 162.000 ;
    END
  END la_data_in_core[112]
  PIN la_data_in_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.930 156.000 1888.210 162.000 ;
    END
  END la_data_in_core[113]
  PIN la_data_in_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.350 156.000 1900.630 162.000 ;
    END
  END la_data_in_core[114]
  PIN la_data_in_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 156.000 1913.050 162.000 ;
    END
  END la_data_in_core[115]
  PIN la_data_in_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.190 156.000 1925.470 162.000 ;
    END
  END la_data_in_core[116]
  PIN la_data_in_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.610 156.000 1937.890 162.000 ;
    END
  END la_data_in_core[117]
  PIN la_data_in_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.030 156.000 1950.310 162.000 ;
    END
  END la_data_in_core[118]
  PIN la_data_in_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.450 156.000 1962.730 162.000 ;
    END
  END la_data_in_core[119]
  PIN la_data_in_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 156.000 621.370 162.000 ;
    END
  END la_data_in_core[11]
  PIN la_data_in_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.870 156.000 1975.150 162.000 ;
    END
  END la_data_in_core[120]
  PIN la_data_in_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.290 156.000 1987.570 162.000 ;
    END
  END la_data_in_core[121]
  PIN la_data_in_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.710 156.000 1999.990 162.000 ;
    END
  END la_data_in_core[122]
  PIN la_data_in_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.130 156.000 2012.410 162.000 ;
    END
  END la_data_in_core[123]
  PIN la_data_in_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.550 156.000 2024.830 162.000 ;
    END
  END la_data_in_core[124]
  PIN la_data_in_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.970 156.000 2037.250 162.000 ;
    END
  END la_data_in_core[125]
  PIN la_data_in_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2049.390 156.000 2049.670 162.000 ;
    END
  END la_data_in_core[126]
  PIN la_data_in_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2061.810 156.000 2062.090 162.000 ;
    END
  END la_data_in_core[127]
  PIN la_data_in_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 156.000 633.790 162.000 ;
    END
  END la_data_in_core[12]
  PIN la_data_in_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 156.000 646.210 162.000 ;
    END
  END la_data_in_core[13]
  PIN la_data_in_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 156.000 658.630 162.000 ;
    END
  END la_data_in_core[14]
  PIN la_data_in_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 156.000 671.050 162.000 ;
    END
  END la_data_in_core[15]
  PIN la_data_in_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 156.000 683.470 162.000 ;
    END
  END la_data_in_core[16]
  PIN la_data_in_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 156.000 695.890 162.000 ;
    END
  END la_data_in_core[17]
  PIN la_data_in_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 156.000 708.310 162.000 ;
    END
  END la_data_in_core[18]
  PIN la_data_in_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 156.000 720.730 162.000 ;
    END
  END la_data_in_core[19]
  PIN la_data_in_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 156.000 497.170 162.000 ;
    END
  END la_data_in_core[1]
  PIN la_data_in_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 156.000 733.150 162.000 ;
    END
  END la_data_in_core[20]
  PIN la_data_in_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 156.000 745.570 162.000 ;
    END
  END la_data_in_core[21]
  PIN la_data_in_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 156.000 757.990 162.000 ;
    END
  END la_data_in_core[22]
  PIN la_data_in_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 156.000 770.410 162.000 ;
    END
  END la_data_in_core[23]
  PIN la_data_in_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 156.000 782.830 162.000 ;
    END
  END la_data_in_core[24]
  PIN la_data_in_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 156.000 795.250 162.000 ;
    END
  END la_data_in_core[25]
  PIN la_data_in_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 156.000 807.670 162.000 ;
    END
  END la_data_in_core[26]
  PIN la_data_in_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 156.000 820.090 162.000 ;
    END
  END la_data_in_core[27]
  PIN la_data_in_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 156.000 832.510 162.000 ;
    END
  END la_data_in_core[28]
  PIN la_data_in_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 156.000 844.930 162.000 ;
    END
  END la_data_in_core[29]
  PIN la_data_in_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 156.000 509.590 162.000 ;
    END
  END la_data_in_core[2]
  PIN la_data_in_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 156.000 857.350 162.000 ;
    END
  END la_data_in_core[30]
  PIN la_data_in_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 156.000 869.770 162.000 ;
    END
  END la_data_in_core[31]
  PIN la_data_in_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 156.000 882.190 162.000 ;
    END
  END la_data_in_core[32]
  PIN la_data_in_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 156.000 894.610 162.000 ;
    END
  END la_data_in_core[33]
  PIN la_data_in_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 156.000 907.030 162.000 ;
    END
  END la_data_in_core[34]
  PIN la_data_in_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 156.000 919.450 162.000 ;
    END
  END la_data_in_core[35]
  PIN la_data_in_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 156.000 931.870 162.000 ;
    END
  END la_data_in_core[36]
  PIN la_data_in_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 156.000 944.290 162.000 ;
    END
  END la_data_in_core[37]
  PIN la_data_in_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 156.000 956.710 162.000 ;
    END
  END la_data_in_core[38]
  PIN la_data_in_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 156.000 969.130 162.000 ;
    END
  END la_data_in_core[39]
  PIN la_data_in_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 156.000 522.010 162.000 ;
    END
  END la_data_in_core[3]
  PIN la_data_in_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 156.000 981.550 162.000 ;
    END
  END la_data_in_core[40]
  PIN la_data_in_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 156.000 993.970 162.000 ;
    END
  END la_data_in_core[41]
  PIN la_data_in_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.110 156.000 1006.390 162.000 ;
    END
  END la_data_in_core[42]
  PIN la_data_in_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 156.000 1018.810 162.000 ;
    END
  END la_data_in_core[43]
  PIN la_data_in_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 156.000 1031.230 162.000 ;
    END
  END la_data_in_core[44]
  PIN la_data_in_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 156.000 1043.650 162.000 ;
    END
  END la_data_in_core[45]
  PIN la_data_in_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 156.000 1056.070 162.000 ;
    END
  END la_data_in_core[46]
  PIN la_data_in_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 156.000 1068.490 162.000 ;
    END
  END la_data_in_core[47]
  PIN la_data_in_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 156.000 1080.910 162.000 ;
    END
  END la_data_in_core[48]
  PIN la_data_in_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 156.000 1093.330 162.000 ;
    END
  END la_data_in_core[49]
  PIN la_data_in_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 156.000 534.430 162.000 ;
    END
  END la_data_in_core[4]
  PIN la_data_in_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 156.000 1105.750 162.000 ;
    END
  END la_data_in_core[50]
  PIN la_data_in_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 156.000 1118.170 162.000 ;
    END
  END la_data_in_core[51]
  PIN la_data_in_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 156.000 1130.590 162.000 ;
    END
  END la_data_in_core[52]
  PIN la_data_in_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.730 156.000 1143.010 162.000 ;
    END
  END la_data_in_core[53]
  PIN la_data_in_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.150 156.000 1155.430 162.000 ;
    END
  END la_data_in_core[54]
  PIN la_data_in_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 156.000 1167.850 162.000 ;
    END
  END la_data_in_core[55]
  PIN la_data_in_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.990 156.000 1180.270 162.000 ;
    END
  END la_data_in_core[56]
  PIN la_data_in_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.410 156.000 1192.690 162.000 ;
    END
  END la_data_in_core[57]
  PIN la_data_in_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.830 156.000 1205.110 162.000 ;
    END
  END la_data_in_core[58]
  PIN la_data_in_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 156.000 1217.530 162.000 ;
    END
  END la_data_in_core[59]
  PIN la_data_in_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 156.000 546.850 162.000 ;
    END
  END la_data_in_core[5]
  PIN la_data_in_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.670 156.000 1229.950 162.000 ;
    END
  END la_data_in_core[60]
  PIN la_data_in_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.090 156.000 1242.370 162.000 ;
    END
  END la_data_in_core[61]
  PIN la_data_in_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.510 156.000 1254.790 162.000 ;
    END
  END la_data_in_core[62]
  PIN la_data_in_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 156.000 1267.210 162.000 ;
    END
  END la_data_in_core[63]
  PIN la_data_in_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.350 156.000 1279.630 162.000 ;
    END
  END la_data_in_core[64]
  PIN la_data_in_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 156.000 1292.050 162.000 ;
    END
  END la_data_in_core[65]
  PIN la_data_in_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 156.000 1304.470 162.000 ;
    END
  END la_data_in_core[66]
  PIN la_data_in_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.610 156.000 1316.890 162.000 ;
    END
  END la_data_in_core[67]
  PIN la_data_in_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.030 156.000 1329.310 162.000 ;
    END
  END la_data_in_core[68]
  PIN la_data_in_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.450 156.000 1341.730 162.000 ;
    END
  END la_data_in_core[69]
  PIN la_data_in_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 156.000 559.270 162.000 ;
    END
  END la_data_in_core[6]
  PIN la_data_in_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.870 156.000 1354.150 162.000 ;
    END
  END la_data_in_core[70]
  PIN la_data_in_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.290 156.000 1366.570 162.000 ;
    END
  END la_data_in_core[71]
  PIN la_data_in_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 156.000 1378.990 162.000 ;
    END
  END la_data_in_core[72]
  PIN la_data_in_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 156.000 1391.410 162.000 ;
    END
  END la_data_in_core[73]
  PIN la_data_in_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.550 156.000 1403.830 162.000 ;
    END
  END la_data_in_core[74]
  PIN la_data_in_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.970 156.000 1416.250 162.000 ;
    END
  END la_data_in_core[75]
  PIN la_data_in_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 156.000 1428.670 162.000 ;
    END
  END la_data_in_core[76]
  PIN la_data_in_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.810 156.000 1441.090 162.000 ;
    END
  END la_data_in_core[77]
  PIN la_data_in_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.230 156.000 1453.510 162.000 ;
    END
  END la_data_in_core[78]
  PIN la_data_in_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.650 156.000 1465.930 162.000 ;
    END
  END la_data_in_core[79]
  PIN la_data_in_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 156.000 571.690 162.000 ;
    END
  END la_data_in_core[7]
  PIN la_data_in_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 156.000 1478.350 162.000 ;
    END
  END la_data_in_core[80]
  PIN la_data_in_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 156.000 1490.770 162.000 ;
    END
  END la_data_in_core[81]
  PIN la_data_in_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.910 156.000 1503.190 162.000 ;
    END
  END la_data_in_core[82]
  PIN la_data_in_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 156.000 1515.610 162.000 ;
    END
  END la_data_in_core[83]
  PIN la_data_in_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.750 156.000 1528.030 162.000 ;
    END
  END la_data_in_core[84]
  PIN la_data_in_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.170 156.000 1540.450 162.000 ;
    END
  END la_data_in_core[85]
  PIN la_data_in_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.590 156.000 1552.870 162.000 ;
    END
  END la_data_in_core[86]
  PIN la_data_in_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 156.000 1565.290 162.000 ;
    END
  END la_data_in_core[87]
  PIN la_data_in_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.430 156.000 1577.710 162.000 ;
    END
  END la_data_in_core[88]
  PIN la_data_in_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 156.000 1590.130 162.000 ;
    END
  END la_data_in_core[89]
  PIN la_data_in_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 156.000 584.110 162.000 ;
    END
  END la_data_in_core[8]
  PIN la_data_in_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.270 156.000 1602.550 162.000 ;
    END
  END la_data_in_core[90]
  PIN la_data_in_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.690 156.000 1614.970 162.000 ;
    END
  END la_data_in_core[91]
  PIN la_data_in_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.110 156.000 1627.390 162.000 ;
    END
  END la_data_in_core[92]
  PIN la_data_in_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 156.000 1639.810 162.000 ;
    END
  END la_data_in_core[93]
  PIN la_data_in_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 156.000 1652.230 162.000 ;
    END
  END la_data_in_core[94]
  PIN la_data_in_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 156.000 1664.650 162.000 ;
    END
  END la_data_in_core[95]
  PIN la_data_in_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.790 156.000 1677.070 162.000 ;
    END
  END la_data_in_core[96]
  PIN la_data_in_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.210 156.000 1689.490 162.000 ;
    END
  END la_data_in_core[97]
  PIN la_data_in_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.630 156.000 1701.910 162.000 ;
    END
  END la_data_in_core[98]
  PIN la_data_in_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.050 156.000 1714.330 162.000 ;
    END
  END la_data_in_core[99]
  PIN la_data_in_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 156.000 596.530 162.000 ;
    END
  END la_data_in_core[9]
  PIN la_data_in_mprj[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 -2.000 65.230 4.000 ;
    END
  END la_data_in_mprj[0]
  PIN la_data_in_mprj[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 -2.000 1359.670 4.000 ;
    END
  END la_data_in_mprj[100]
  PIN la_data_in_mprj[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.270 -2.000 1372.550 4.000 ;
    END
  END la_data_in_mprj[101]
  PIN la_data_in_mprj[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 -2.000 1385.430 4.000 ;
    END
  END la_data_in_mprj[102]
  PIN la_data_in_mprj[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.030 -2.000 1398.310 4.000 ;
    END
  END la_data_in_mprj[103]
  PIN la_data_in_mprj[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 -2.000 1411.190 4.000 ;
    END
  END la_data_in_mprj[104]
  PIN la_data_in_mprj[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.790 -2.000 1424.070 4.000 ;
    END
  END la_data_in_mprj[105]
  PIN la_data_in_mprj[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.670 -2.000 1436.950 4.000 ;
    END
  END la_data_in_mprj[106]
  PIN la_data_in_mprj[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 -2.000 1449.830 4.000 ;
    END
  END la_data_in_mprj[107]
  PIN la_data_in_mprj[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 -2.000 1462.710 4.000 ;
    END
  END la_data_in_mprj[108]
  PIN la_data_in_mprj[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 -2.000 1475.590 4.000 ;
    END
  END la_data_in_mprj[109]
  PIN la_data_in_mprj[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 -2.000 194.030 4.000 ;
    END
  END la_data_in_mprj[10]
  PIN la_data_in_mprj[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.190 -2.000 1488.470 4.000 ;
    END
  END la_data_in_mprj[110]
  PIN la_data_in_mprj[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.070 -2.000 1501.350 4.000 ;
    END
  END la_data_in_mprj[111]
  PIN la_data_in_mprj[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.950 -2.000 1514.230 4.000 ;
    END
  END la_data_in_mprj[112]
  PIN la_data_in_mprj[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.830 -2.000 1527.110 4.000 ;
    END
  END la_data_in_mprj[113]
  PIN la_data_in_mprj[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.710 -2.000 1539.990 4.000 ;
    END
  END la_data_in_mprj[114]
  PIN la_data_in_mprj[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.590 -2.000 1552.870 4.000 ;
    END
  END la_data_in_mprj[115]
  PIN la_data_in_mprj[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.470 -2.000 1565.750 4.000 ;
    END
  END la_data_in_mprj[116]
  PIN la_data_in_mprj[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.350 -2.000 1578.630 4.000 ;
    END
  END la_data_in_mprj[117]
  PIN la_data_in_mprj[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 -2.000 1591.510 4.000 ;
    END
  END la_data_in_mprj[118]
  PIN la_data_in_mprj[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.110 -2.000 1604.390 4.000 ;
    END
  END la_data_in_mprj[119]
  PIN la_data_in_mprj[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 -2.000 206.910 4.000 ;
    END
  END la_data_in_mprj[11]
  PIN la_data_in_mprj[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 -2.000 1617.270 4.000 ;
    END
  END la_data_in_mprj[120]
  PIN la_data_in_mprj[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.870 -2.000 1630.150 4.000 ;
    END
  END la_data_in_mprj[121]
  PIN la_data_in_mprj[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.750 -2.000 1643.030 4.000 ;
    END
  END la_data_in_mprj[122]
  PIN la_data_in_mprj[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.630 -2.000 1655.910 4.000 ;
    END
  END la_data_in_mprj[123]
  PIN la_data_in_mprj[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.510 -2.000 1668.790 4.000 ;
    END
  END la_data_in_mprj[124]
  PIN la_data_in_mprj[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.390 -2.000 1681.670 4.000 ;
    END
  END la_data_in_mprj[125]
  PIN la_data_in_mprj[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.270 -2.000 1694.550 4.000 ;
    END
  END la_data_in_mprj[126]
  PIN la_data_in_mprj[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.150 -2.000 1707.430 4.000 ;
    END
  END la_data_in_mprj[127]
  PIN la_data_in_mprj[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 -2.000 219.790 4.000 ;
    END
  END la_data_in_mprj[12]
  PIN la_data_in_mprj[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 -2.000 232.670 4.000 ;
    END
  END la_data_in_mprj[13]
  PIN la_data_in_mprj[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 -2.000 245.550 4.000 ;
    END
  END la_data_in_mprj[14]
  PIN la_data_in_mprj[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 -2.000 258.430 4.000 ;
    END
  END la_data_in_mprj[15]
  PIN la_data_in_mprj[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 -2.000 271.310 4.000 ;
    END
  END la_data_in_mprj[16]
  PIN la_data_in_mprj[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 -2.000 284.190 4.000 ;
    END
  END la_data_in_mprj[17]
  PIN la_data_in_mprj[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 -2.000 297.070 4.000 ;
    END
  END la_data_in_mprj[18]
  PIN la_data_in_mprj[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 -2.000 309.950 4.000 ;
    END
  END la_data_in_mprj[19]
  PIN la_data_in_mprj[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 -2.000 78.110 4.000 ;
    END
  END la_data_in_mprj[1]
  PIN la_data_in_mprj[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 -2.000 322.830 4.000 ;
    END
  END la_data_in_mprj[20]
  PIN la_data_in_mprj[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 -2.000 335.710 4.000 ;
    END
  END la_data_in_mprj[21]
  PIN la_data_in_mprj[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 -2.000 348.590 4.000 ;
    END
  END la_data_in_mprj[22]
  PIN la_data_in_mprj[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 -2.000 361.470 4.000 ;
    END
  END la_data_in_mprj[23]
  PIN la_data_in_mprj[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 -2.000 374.350 4.000 ;
    END
  END la_data_in_mprj[24]
  PIN la_data_in_mprj[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 -2.000 387.230 4.000 ;
    END
  END la_data_in_mprj[25]
  PIN la_data_in_mprj[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 -2.000 400.110 4.000 ;
    END
  END la_data_in_mprj[26]
  PIN la_data_in_mprj[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 -2.000 412.990 4.000 ;
    END
  END la_data_in_mprj[27]
  PIN la_data_in_mprj[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 -2.000 425.870 4.000 ;
    END
  END la_data_in_mprj[28]
  PIN la_data_in_mprj[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 -2.000 438.750 4.000 ;
    END
  END la_data_in_mprj[29]
  PIN la_data_in_mprj[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 -2.000 90.990 4.000 ;
    END
  END la_data_in_mprj[2]
  PIN la_data_in_mprj[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 -2.000 451.630 4.000 ;
    END
  END la_data_in_mprj[30]
  PIN la_data_in_mprj[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 -2.000 464.510 4.000 ;
    END
  END la_data_in_mprj[31]
  PIN la_data_in_mprj[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 -2.000 477.390 4.000 ;
    END
  END la_data_in_mprj[32]
  PIN la_data_in_mprj[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 -2.000 490.270 4.000 ;
    END
  END la_data_in_mprj[33]
  PIN la_data_in_mprj[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 -2.000 503.150 4.000 ;
    END
  END la_data_in_mprj[34]
  PIN la_data_in_mprj[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 -2.000 516.030 4.000 ;
    END
  END la_data_in_mprj[35]
  PIN la_data_in_mprj[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 -2.000 528.910 4.000 ;
    END
  END la_data_in_mprj[36]
  PIN la_data_in_mprj[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 -2.000 541.790 4.000 ;
    END
  END la_data_in_mprj[37]
  PIN la_data_in_mprj[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 -2.000 554.670 4.000 ;
    END
  END la_data_in_mprj[38]
  PIN la_data_in_mprj[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 -2.000 567.550 4.000 ;
    END
  END la_data_in_mprj[39]
  PIN la_data_in_mprj[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 -2.000 103.870 4.000 ;
    END
  END la_data_in_mprj[3]
  PIN la_data_in_mprj[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 -2.000 580.430 4.000 ;
    END
  END la_data_in_mprj[40]
  PIN la_data_in_mprj[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 -2.000 593.310 4.000 ;
    END
  END la_data_in_mprj[41]
  PIN la_data_in_mprj[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 -2.000 606.190 4.000 ;
    END
  END la_data_in_mprj[42]
  PIN la_data_in_mprj[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 -2.000 619.070 4.000 ;
    END
  END la_data_in_mprj[43]
  PIN la_data_in_mprj[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 -2.000 631.950 4.000 ;
    END
  END la_data_in_mprj[44]
  PIN la_data_in_mprj[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 -2.000 644.830 4.000 ;
    END
  END la_data_in_mprj[45]
  PIN la_data_in_mprj[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 -2.000 657.710 4.000 ;
    END
  END la_data_in_mprj[46]
  PIN la_data_in_mprj[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 -2.000 670.590 4.000 ;
    END
  END la_data_in_mprj[47]
  PIN la_data_in_mprj[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 -2.000 683.470 4.000 ;
    END
  END la_data_in_mprj[48]
  PIN la_data_in_mprj[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 -2.000 696.350 4.000 ;
    END
  END la_data_in_mprj[49]
  PIN la_data_in_mprj[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 -2.000 116.750 4.000 ;
    END
  END la_data_in_mprj[4]
  PIN la_data_in_mprj[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 -2.000 709.230 4.000 ;
    END
  END la_data_in_mprj[50]
  PIN la_data_in_mprj[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 -2.000 722.110 4.000 ;
    END
  END la_data_in_mprj[51]
  PIN la_data_in_mprj[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 -2.000 734.990 4.000 ;
    END
  END la_data_in_mprj[52]
  PIN la_data_in_mprj[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 -2.000 747.870 4.000 ;
    END
  END la_data_in_mprj[53]
  PIN la_data_in_mprj[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 -2.000 760.750 4.000 ;
    END
  END la_data_in_mprj[54]
  PIN la_data_in_mprj[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 -2.000 773.630 4.000 ;
    END
  END la_data_in_mprj[55]
  PIN la_data_in_mprj[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 -2.000 786.510 4.000 ;
    END
  END la_data_in_mprj[56]
  PIN la_data_in_mprj[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 -2.000 799.390 4.000 ;
    END
  END la_data_in_mprj[57]
  PIN la_data_in_mprj[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 -2.000 812.270 4.000 ;
    END
  END la_data_in_mprj[58]
  PIN la_data_in_mprj[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 -2.000 825.150 4.000 ;
    END
  END la_data_in_mprj[59]
  PIN la_data_in_mprj[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 -2.000 129.630 4.000 ;
    END
  END la_data_in_mprj[5]
  PIN la_data_in_mprj[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 -2.000 838.030 4.000 ;
    END
  END la_data_in_mprj[60]
  PIN la_data_in_mprj[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 -2.000 850.910 4.000 ;
    END
  END la_data_in_mprj[61]
  PIN la_data_in_mprj[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 -2.000 863.790 4.000 ;
    END
  END la_data_in_mprj[62]
  PIN la_data_in_mprj[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 -2.000 876.670 4.000 ;
    END
  END la_data_in_mprj[63]
  PIN la_data_in_mprj[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 -2.000 889.550 4.000 ;
    END
  END la_data_in_mprj[64]
  PIN la_data_in_mprj[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.150 -2.000 902.430 4.000 ;
    END
  END la_data_in_mprj[65]
  PIN la_data_in_mprj[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 -2.000 915.310 4.000 ;
    END
  END la_data_in_mprj[66]
  PIN la_data_in_mprj[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 -2.000 928.190 4.000 ;
    END
  END la_data_in_mprj[67]
  PIN la_data_in_mprj[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 -2.000 941.070 4.000 ;
    END
  END la_data_in_mprj[68]
  PIN la_data_in_mprj[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 -2.000 953.950 4.000 ;
    END
  END la_data_in_mprj[69]
  PIN la_data_in_mprj[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 -2.000 142.510 4.000 ;
    END
  END la_data_in_mprj[6]
  PIN la_data_in_mprj[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 -2.000 966.830 4.000 ;
    END
  END la_data_in_mprj[70]
  PIN la_data_in_mprj[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 -2.000 986.150 4.000 ;
    END
  END la_data_in_mprj[71]
  PIN la_data_in_mprj[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 -2.000 999.030 4.000 ;
    END
  END la_data_in_mprj[72]
  PIN la_data_in_mprj[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 -2.000 1011.910 4.000 ;
    END
  END la_data_in_mprj[73]
  PIN la_data_in_mprj[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 -2.000 1024.790 4.000 ;
    END
  END la_data_in_mprj[74]
  PIN la_data_in_mprj[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 -2.000 1037.670 4.000 ;
    END
  END la_data_in_mprj[75]
  PIN la_data_in_mprj[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 -2.000 1050.550 4.000 ;
    END
  END la_data_in_mprj[76]
  PIN la_data_in_mprj[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 -2.000 1063.430 4.000 ;
    END
  END la_data_in_mprj[77]
  PIN la_data_in_mprj[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 -2.000 1076.310 4.000 ;
    END
  END la_data_in_mprj[78]
  PIN la_data_in_mprj[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 -2.000 1089.190 4.000 ;
    END
  END la_data_in_mprj[79]
  PIN la_data_in_mprj[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 -2.000 155.390 4.000 ;
    END
  END la_data_in_mprj[7]
  PIN la_data_in_mprj[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 -2.000 1102.070 4.000 ;
    END
  END la_data_in_mprj[80]
  PIN la_data_in_mprj[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 -2.000 1114.950 4.000 ;
    END
  END la_data_in_mprj[81]
  PIN la_data_in_mprj[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.550 -2.000 1127.830 4.000 ;
    END
  END la_data_in_mprj[82]
  PIN la_data_in_mprj[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.430 -2.000 1140.710 4.000 ;
    END
  END la_data_in_mprj[83]
  PIN la_data_in_mprj[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.310 -2.000 1153.590 4.000 ;
    END
  END la_data_in_mprj[84]
  PIN la_data_in_mprj[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.190 -2.000 1166.470 4.000 ;
    END
  END la_data_in_mprj[85]
  PIN la_data_in_mprj[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.070 -2.000 1179.350 4.000 ;
    END
  END la_data_in_mprj[86]
  PIN la_data_in_mprj[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 -2.000 1192.230 4.000 ;
    END
  END la_data_in_mprj[87]
  PIN la_data_in_mprj[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.830 -2.000 1205.110 4.000 ;
    END
  END la_data_in_mprj[88]
  PIN la_data_in_mprj[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.710 -2.000 1217.990 4.000 ;
    END
  END la_data_in_mprj[89]
  PIN la_data_in_mprj[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 -2.000 168.270 4.000 ;
    END
  END la_data_in_mprj[8]
  PIN la_data_in_mprj[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.590 -2.000 1230.870 4.000 ;
    END
  END la_data_in_mprj[90]
  PIN la_data_in_mprj[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 -2.000 1243.750 4.000 ;
    END
  END la_data_in_mprj[91]
  PIN la_data_in_mprj[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 -2.000 1256.630 4.000 ;
    END
  END la_data_in_mprj[92]
  PIN la_data_in_mprj[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.230 -2.000 1269.510 4.000 ;
    END
  END la_data_in_mprj[93]
  PIN la_data_in_mprj[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 -2.000 1282.390 4.000 ;
    END
  END la_data_in_mprj[94]
  PIN la_data_in_mprj[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 -2.000 1295.270 4.000 ;
    END
  END la_data_in_mprj[95]
  PIN la_data_in_mprj[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 -2.000 1308.150 4.000 ;
    END
  END la_data_in_mprj[96]
  PIN la_data_in_mprj[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 -2.000 1321.030 4.000 ;
    END
  END la_data_in_mprj[97]
  PIN la_data_in_mprj[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 -2.000 1333.910 4.000 ;
    END
  END la_data_in_mprj[98]
  PIN la_data_in_mprj[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 -2.000 1346.790 4.000 ;
    END
  END la_data_in_mprj[99]
  PIN la_data_in_mprj[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 -2.000 181.150 4.000 ;
    END
  END la_data_in_mprj[9]
  PIN la_data_out_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 156.000 488.890 162.000 ;
    END
  END la_data_out_core[0]
  PIN la_data_out_core[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.610 156.000 1730.890 162.000 ;
    END
  END la_data_out_core[100]
  PIN la_data_out_core[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.030 156.000 1743.310 162.000 ;
    END
  END la_data_out_core[101]
  PIN la_data_out_core[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.450 156.000 1755.730 162.000 ;
    END
  END la_data_out_core[102]
  PIN la_data_out_core[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 156.000 1768.150 162.000 ;
    END
  END la_data_out_core[103]
  PIN la_data_out_core[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.290 156.000 1780.570 162.000 ;
    END
  END la_data_out_core[104]
  PIN la_data_out_core[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.710 156.000 1792.990 162.000 ;
    END
  END la_data_out_core[105]
  PIN la_data_out_core[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.130 156.000 1805.410 162.000 ;
    END
  END la_data_out_core[106]
  PIN la_data_out_core[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.550 156.000 1817.830 162.000 ;
    END
  END la_data_out_core[107]
  PIN la_data_out_core[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.970 156.000 1830.250 162.000 ;
    END
  END la_data_out_core[108]
  PIN la_data_out_core[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.390 156.000 1842.670 162.000 ;
    END
  END la_data_out_core[109]
  PIN la_data_out_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 156.000 613.090 162.000 ;
    END
  END la_data_out_core[10]
  PIN la_data_out_core[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 156.000 1855.090 162.000 ;
    END
  END la_data_out_core[110]
  PIN la_data_out_core[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.230 156.000 1867.510 162.000 ;
    END
  END la_data_out_core[111]
  PIN la_data_out_core[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.650 156.000 1879.930 162.000 ;
    END
  END la_data_out_core[112]
  PIN la_data_out_core[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.070 156.000 1892.350 162.000 ;
    END
  END la_data_out_core[113]
  PIN la_data_out_core[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.490 156.000 1904.770 162.000 ;
    END
  END la_data_out_core[114]
  PIN la_data_out_core[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.910 156.000 1917.190 162.000 ;
    END
  END la_data_out_core[115]
  PIN la_data_out_core[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.330 156.000 1929.610 162.000 ;
    END
  END la_data_out_core[116]
  PIN la_data_out_core[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 156.000 1942.030 162.000 ;
    END
  END la_data_out_core[117]
  PIN la_data_out_core[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.170 156.000 1954.450 162.000 ;
    END
  END la_data_out_core[118]
  PIN la_data_out_core[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.590 156.000 1966.870 162.000 ;
    END
  END la_data_out_core[119]
  PIN la_data_out_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 156.000 625.510 162.000 ;
    END
  END la_data_out_core[11]
  PIN la_data_out_core[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.010 156.000 1979.290 162.000 ;
    END
  END la_data_out_core[120]
  PIN la_data_out_core[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.430 156.000 1991.710 162.000 ;
    END
  END la_data_out_core[121]
  PIN la_data_out_core[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.850 156.000 2004.130 162.000 ;
    END
  END la_data_out_core[122]
  PIN la_data_out_core[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2016.270 156.000 2016.550 162.000 ;
    END
  END la_data_out_core[123]
  PIN la_data_out_core[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.690 156.000 2028.970 162.000 ;
    END
  END la_data_out_core[124]
  PIN la_data_out_core[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.110 156.000 2041.390 162.000 ;
    END
  END la_data_out_core[125]
  PIN la_data_out_core[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.530 156.000 2053.810 162.000 ;
    END
  END la_data_out_core[126]
  PIN la_data_out_core[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.950 156.000 2066.230 162.000 ;
    END
  END la_data_out_core[127]
  PIN la_data_out_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 156.000 637.930 162.000 ;
    END
  END la_data_out_core[12]
  PIN la_data_out_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 156.000 650.350 162.000 ;
    END
  END la_data_out_core[13]
  PIN la_data_out_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 156.000 662.770 162.000 ;
    END
  END la_data_out_core[14]
  PIN la_data_out_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 156.000 675.190 162.000 ;
    END
  END la_data_out_core[15]
  PIN la_data_out_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 156.000 687.610 162.000 ;
    END
  END la_data_out_core[16]
  PIN la_data_out_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 156.000 700.030 162.000 ;
    END
  END la_data_out_core[17]
  PIN la_data_out_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 156.000 712.450 162.000 ;
    END
  END la_data_out_core[18]
  PIN la_data_out_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 156.000 724.870 162.000 ;
    END
  END la_data_out_core[19]
  PIN la_data_out_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 156.000 501.310 162.000 ;
    END
  END la_data_out_core[1]
  PIN la_data_out_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 156.000 737.290 162.000 ;
    END
  END la_data_out_core[20]
  PIN la_data_out_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 156.000 749.710 162.000 ;
    END
  END la_data_out_core[21]
  PIN la_data_out_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 156.000 762.130 162.000 ;
    END
  END la_data_out_core[22]
  PIN la_data_out_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 156.000 774.550 162.000 ;
    END
  END la_data_out_core[23]
  PIN la_data_out_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 156.000 786.970 162.000 ;
    END
  END la_data_out_core[24]
  PIN la_data_out_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 156.000 799.390 162.000 ;
    END
  END la_data_out_core[25]
  PIN la_data_out_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 156.000 811.810 162.000 ;
    END
  END la_data_out_core[26]
  PIN la_data_out_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 156.000 824.230 162.000 ;
    END
  END la_data_out_core[27]
  PIN la_data_out_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 156.000 836.650 162.000 ;
    END
  END la_data_out_core[28]
  PIN la_data_out_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 156.000 849.070 162.000 ;
    END
  END la_data_out_core[29]
  PIN la_data_out_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 156.000 513.730 162.000 ;
    END
  END la_data_out_core[2]
  PIN la_data_out_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 156.000 861.490 162.000 ;
    END
  END la_data_out_core[30]
  PIN la_data_out_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 156.000 873.910 162.000 ;
    END
  END la_data_out_core[31]
  PIN la_data_out_core[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 156.000 886.330 162.000 ;
    END
  END la_data_out_core[32]
  PIN la_data_out_core[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 156.000 898.750 162.000 ;
    END
  END la_data_out_core[33]
  PIN la_data_out_core[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 156.000 911.170 162.000 ;
    END
  END la_data_out_core[34]
  PIN la_data_out_core[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.310 156.000 923.590 162.000 ;
    END
  END la_data_out_core[35]
  PIN la_data_out_core[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 156.000 936.010 162.000 ;
    END
  END la_data_out_core[36]
  PIN la_data_out_core[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 156.000 948.430 162.000 ;
    END
  END la_data_out_core[37]
  PIN la_data_out_core[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.570 156.000 960.850 162.000 ;
    END
  END la_data_out_core[38]
  PIN la_data_out_core[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 156.000 973.270 162.000 ;
    END
  END la_data_out_core[39]
  PIN la_data_out_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 156.000 526.150 162.000 ;
    END
  END la_data_out_core[3]
  PIN la_data_out_core[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 156.000 985.690 162.000 ;
    END
  END la_data_out_core[40]
  PIN la_data_out_core[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 156.000 998.110 162.000 ;
    END
  END la_data_out_core[41]
  PIN la_data_out_core[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 156.000 1010.530 162.000 ;
    END
  END la_data_out_core[42]
  PIN la_data_out_core[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.670 156.000 1022.950 162.000 ;
    END
  END la_data_out_core[43]
  PIN la_data_out_core[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 156.000 1035.370 162.000 ;
    END
  END la_data_out_core[44]
  PIN la_data_out_core[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 156.000 1047.790 162.000 ;
    END
  END la_data_out_core[45]
  PIN la_data_out_core[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 156.000 1060.210 162.000 ;
    END
  END la_data_out_core[46]
  PIN la_data_out_core[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 156.000 1072.630 162.000 ;
    END
  END la_data_out_core[47]
  PIN la_data_out_core[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 156.000 1085.050 162.000 ;
    END
  END la_data_out_core[48]
  PIN la_data_out_core[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 156.000 1097.470 162.000 ;
    END
  END la_data_out_core[49]
  PIN la_data_out_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 156.000 538.570 162.000 ;
    END
  END la_data_out_core[4]
  PIN la_data_out_core[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 156.000 1109.890 162.000 ;
    END
  END la_data_out_core[50]
  PIN la_data_out_core[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 156.000 1122.310 162.000 ;
    END
  END la_data_out_core[51]
  PIN la_data_out_core[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 156.000 1134.730 162.000 ;
    END
  END la_data_out_core[52]
  PIN la_data_out_core[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 156.000 1147.150 162.000 ;
    END
  END la_data_out_core[53]
  PIN la_data_out_core[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 156.000 1159.570 162.000 ;
    END
  END la_data_out_core[54]
  PIN la_data_out_core[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 156.000 1171.990 162.000 ;
    END
  END la_data_out_core[55]
  PIN la_data_out_core[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 156.000 1184.410 162.000 ;
    END
  END la_data_out_core[56]
  PIN la_data_out_core[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 156.000 1196.830 162.000 ;
    END
  END la_data_out_core[57]
  PIN la_data_out_core[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 156.000 1209.250 162.000 ;
    END
  END la_data_out_core[58]
  PIN la_data_out_core[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 156.000 1221.670 162.000 ;
    END
  END la_data_out_core[59]
  PIN la_data_out_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 156.000 550.990 162.000 ;
    END
  END la_data_out_core[5]
  PIN la_data_out_core[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 156.000 1234.090 162.000 ;
    END
  END la_data_out_core[60]
  PIN la_data_out_core[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 156.000 1246.510 162.000 ;
    END
  END la_data_out_core[61]
  PIN la_data_out_core[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 156.000 1258.930 162.000 ;
    END
  END la_data_out_core[62]
  PIN la_data_out_core[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.070 156.000 1271.350 162.000 ;
    END
  END la_data_out_core[63]
  PIN la_data_out_core[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.490 156.000 1283.770 162.000 ;
    END
  END la_data_out_core[64]
  PIN la_data_out_core[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.910 156.000 1296.190 162.000 ;
    END
  END la_data_out_core[65]
  PIN la_data_out_core[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 156.000 1308.610 162.000 ;
    END
  END la_data_out_core[66]
  PIN la_data_out_core[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 156.000 1321.030 162.000 ;
    END
  END la_data_out_core[67]
  PIN la_data_out_core[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 156.000 1333.450 162.000 ;
    END
  END la_data_out_core[68]
  PIN la_data_out_core[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.590 156.000 1345.870 162.000 ;
    END
  END la_data_out_core[69]
  PIN la_data_out_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 156.000 563.410 162.000 ;
    END
  END la_data_out_core[6]
  PIN la_data_out_core[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 156.000 1358.290 162.000 ;
    END
  END la_data_out_core[70]
  PIN la_data_out_core[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 156.000 1370.710 162.000 ;
    END
  END la_data_out_core[71]
  PIN la_data_out_core[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.850 156.000 1383.130 162.000 ;
    END
  END la_data_out_core[72]
  PIN la_data_out_core[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.270 156.000 1395.550 162.000 ;
    END
  END la_data_out_core[73]
  PIN la_data_out_core[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 156.000 1407.970 162.000 ;
    END
  END la_data_out_core[74]
  PIN la_data_out_core[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 156.000 1420.390 162.000 ;
    END
  END la_data_out_core[75]
  PIN la_data_out_core[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.530 156.000 1432.810 162.000 ;
    END
  END la_data_out_core[76]
  PIN la_data_out_core[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.950 156.000 1445.230 162.000 ;
    END
  END la_data_out_core[77]
  PIN la_data_out_core[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 156.000 1457.650 162.000 ;
    END
  END la_data_out_core[78]
  PIN la_data_out_core[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.790 156.000 1470.070 162.000 ;
    END
  END la_data_out_core[79]
  PIN la_data_out_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 156.000 575.830 162.000 ;
    END
  END la_data_out_core[7]
  PIN la_data_out_core[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.210 156.000 1482.490 162.000 ;
    END
  END la_data_out_core[80]
  PIN la_data_out_core[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.630 156.000 1494.910 162.000 ;
    END
  END la_data_out_core[81]
  PIN la_data_out_core[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 156.000 1507.330 162.000 ;
    END
  END la_data_out_core[82]
  PIN la_data_out_core[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.470 156.000 1519.750 162.000 ;
    END
  END la_data_out_core[83]
  PIN la_data_out_core[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.890 156.000 1532.170 162.000 ;
    END
  END la_data_out_core[84]
  PIN la_data_out_core[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.310 156.000 1544.590 162.000 ;
    END
  END la_data_out_core[85]
  PIN la_data_out_core[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.730 156.000 1557.010 162.000 ;
    END
  END la_data_out_core[86]
  PIN la_data_out_core[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.150 156.000 1569.430 162.000 ;
    END
  END la_data_out_core[87]
  PIN la_data_out_core[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.570 156.000 1581.850 162.000 ;
    END
  END la_data_out_core[88]
  PIN la_data_out_core[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990 156.000 1594.270 162.000 ;
    END
  END la_data_out_core[89]
  PIN la_data_out_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 156.000 588.250 162.000 ;
    END
  END la_data_out_core[8]
  PIN la_data_out_core[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.410 156.000 1606.690 162.000 ;
    END
  END la_data_out_core[90]
  PIN la_data_out_core[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.830 156.000 1619.110 162.000 ;
    END
  END la_data_out_core[91]
  PIN la_data_out_core[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.250 156.000 1631.530 162.000 ;
    END
  END la_data_out_core[92]
  PIN la_data_out_core[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 156.000 1643.950 162.000 ;
    END
  END la_data_out_core[93]
  PIN la_data_out_core[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.090 156.000 1656.370 162.000 ;
    END
  END la_data_out_core[94]
  PIN la_data_out_core[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.510 156.000 1668.790 162.000 ;
    END
  END la_data_out_core[95]
  PIN la_data_out_core[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 156.000 1681.210 162.000 ;
    END
  END la_data_out_core[96]
  PIN la_data_out_core[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.350 156.000 1693.630 162.000 ;
    END
  END la_data_out_core[97]
  PIN la_data_out_core[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 156.000 1706.050 162.000 ;
    END
  END la_data_out_core[98]
  PIN la_data_out_core[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 156.000 1718.470 162.000 ;
    END
  END la_data_out_core[99]
  PIN la_data_out_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 156.000 600.670 162.000 ;
    END
  END la_data_out_core[9]
  PIN la_data_out_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 -2.000 68.450 4.000 ;
    END
  END la_data_out_mprj[0]
  PIN la_data_out_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 -2.000 1362.890 4.000 ;
    END
  END la_data_out_mprj[100]
  PIN la_data_out_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.490 -2.000 1375.770 4.000 ;
    END
  END la_data_out_mprj[101]
  PIN la_data_out_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.370 -2.000 1388.650 4.000 ;
    END
  END la_data_out_mprj[102]
  PIN la_data_out_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 -2.000 1401.530 4.000 ;
    END
  END la_data_out_mprj[103]
  PIN la_data_out_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.130 -2.000 1414.410 4.000 ;
    END
  END la_data_out_mprj[104]
  PIN la_data_out_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 -2.000 1427.290 4.000 ;
    END
  END la_data_out_mprj[105]
  PIN la_data_out_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 -2.000 1440.170 4.000 ;
    END
  END la_data_out_mprj[106]
  PIN la_data_out_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.770 -2.000 1453.050 4.000 ;
    END
  END la_data_out_mprj[107]
  PIN la_data_out_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.650 -2.000 1465.930 4.000 ;
    END
  END la_data_out_mprj[108]
  PIN la_data_out_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.530 -2.000 1478.810 4.000 ;
    END
  END la_data_out_mprj[109]
  PIN la_data_out_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 -2.000 197.250 4.000 ;
    END
  END la_data_out_mprj[10]
  PIN la_data_out_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 -2.000 1491.690 4.000 ;
    END
  END la_data_out_mprj[110]
  PIN la_data_out_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 -2.000 1504.570 4.000 ;
    END
  END la_data_out_mprj[111]
  PIN la_data_out_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.170 -2.000 1517.450 4.000 ;
    END
  END la_data_out_mprj[112]
  PIN la_data_out_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.050 -2.000 1530.330 4.000 ;
    END
  END la_data_out_mprj[113]
  PIN la_data_out_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 -2.000 1543.210 4.000 ;
    END
  END la_data_out_mprj[114]
  PIN la_data_out_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.810 -2.000 1556.090 4.000 ;
    END
  END la_data_out_mprj[115]
  PIN la_data_out_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.690 -2.000 1568.970 4.000 ;
    END
  END la_data_out_mprj[116]
  PIN la_data_out_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.570 -2.000 1581.850 4.000 ;
    END
  END la_data_out_mprj[117]
  PIN la_data_out_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.450 -2.000 1594.730 4.000 ;
    END
  END la_data_out_mprj[118]
  PIN la_data_out_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.330 -2.000 1607.610 4.000 ;
    END
  END la_data_out_mprj[119]
  PIN la_data_out_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 -2.000 210.130 4.000 ;
    END
  END la_data_out_mprj[11]
  PIN la_data_out_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.210 -2.000 1620.490 4.000 ;
    END
  END la_data_out_mprj[120]
  PIN la_data_out_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.090 -2.000 1633.370 4.000 ;
    END
  END la_data_out_mprj[121]
  PIN la_data_out_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.970 -2.000 1646.250 4.000 ;
    END
  END la_data_out_mprj[122]
  PIN la_data_out_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 -2.000 1659.130 4.000 ;
    END
  END la_data_out_mprj[123]
  PIN la_data_out_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.730 -2.000 1672.010 4.000 ;
    END
  END la_data_out_mprj[124]
  PIN la_data_out_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.610 -2.000 1684.890 4.000 ;
    END
  END la_data_out_mprj[125]
  PIN la_data_out_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 -2.000 1697.770 4.000 ;
    END
  END la_data_out_mprj[126]
  PIN la_data_out_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.370 -2.000 1710.650 4.000 ;
    END
  END la_data_out_mprj[127]
  PIN la_data_out_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 -2.000 223.010 4.000 ;
    END
  END la_data_out_mprj[12]
  PIN la_data_out_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 -2.000 235.890 4.000 ;
    END
  END la_data_out_mprj[13]
  PIN la_data_out_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 -2.000 248.770 4.000 ;
    END
  END la_data_out_mprj[14]
  PIN la_data_out_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 -2.000 261.650 4.000 ;
    END
  END la_data_out_mprj[15]
  PIN la_data_out_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 -2.000 274.530 4.000 ;
    END
  END la_data_out_mprj[16]
  PIN la_data_out_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 -2.000 287.410 4.000 ;
    END
  END la_data_out_mprj[17]
  PIN la_data_out_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 -2.000 300.290 4.000 ;
    END
  END la_data_out_mprj[18]
  PIN la_data_out_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 -2.000 313.170 4.000 ;
    END
  END la_data_out_mprj[19]
  PIN la_data_out_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 -2.000 81.330 4.000 ;
    END
  END la_data_out_mprj[1]
  PIN la_data_out_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 -2.000 326.050 4.000 ;
    END
  END la_data_out_mprj[20]
  PIN la_data_out_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 -2.000 338.930 4.000 ;
    END
  END la_data_out_mprj[21]
  PIN la_data_out_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 -2.000 351.810 4.000 ;
    END
  END la_data_out_mprj[22]
  PIN la_data_out_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 -2.000 364.690 4.000 ;
    END
  END la_data_out_mprj[23]
  PIN la_data_out_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 -2.000 377.570 4.000 ;
    END
  END la_data_out_mprj[24]
  PIN la_data_out_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 -2.000 390.450 4.000 ;
    END
  END la_data_out_mprj[25]
  PIN la_data_out_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 -2.000 403.330 4.000 ;
    END
  END la_data_out_mprj[26]
  PIN la_data_out_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 -2.000 416.210 4.000 ;
    END
  END la_data_out_mprj[27]
  PIN la_data_out_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 -2.000 429.090 4.000 ;
    END
  END la_data_out_mprj[28]
  PIN la_data_out_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 -2.000 441.970 4.000 ;
    END
  END la_data_out_mprj[29]
  PIN la_data_out_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 -2.000 94.210 4.000 ;
    END
  END la_data_out_mprj[2]
  PIN la_data_out_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 -2.000 454.850 4.000 ;
    END
  END la_data_out_mprj[30]
  PIN la_data_out_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 -2.000 467.730 4.000 ;
    END
  END la_data_out_mprj[31]
  PIN la_data_out_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 -2.000 480.610 4.000 ;
    END
  END la_data_out_mprj[32]
  PIN la_data_out_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 -2.000 493.490 4.000 ;
    END
  END la_data_out_mprj[33]
  PIN la_data_out_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 -2.000 506.370 4.000 ;
    END
  END la_data_out_mprj[34]
  PIN la_data_out_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 -2.000 519.250 4.000 ;
    END
  END la_data_out_mprj[35]
  PIN la_data_out_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 -2.000 532.130 4.000 ;
    END
  END la_data_out_mprj[36]
  PIN la_data_out_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 -2.000 545.010 4.000 ;
    END
  END la_data_out_mprj[37]
  PIN la_data_out_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 -2.000 557.890 4.000 ;
    END
  END la_data_out_mprj[38]
  PIN la_data_out_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 -2.000 570.770 4.000 ;
    END
  END la_data_out_mprj[39]
  PIN la_data_out_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 -2.000 107.090 4.000 ;
    END
  END la_data_out_mprj[3]
  PIN la_data_out_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 -2.000 583.650 4.000 ;
    END
  END la_data_out_mprj[40]
  PIN la_data_out_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 -2.000 596.530 4.000 ;
    END
  END la_data_out_mprj[41]
  PIN la_data_out_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 -2.000 609.410 4.000 ;
    END
  END la_data_out_mprj[42]
  PIN la_data_out_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 -2.000 622.290 4.000 ;
    END
  END la_data_out_mprj[43]
  PIN la_data_out_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 -2.000 635.170 4.000 ;
    END
  END la_data_out_mprj[44]
  PIN la_data_out_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 -2.000 648.050 4.000 ;
    END
  END la_data_out_mprj[45]
  PIN la_data_out_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 -2.000 660.930 4.000 ;
    END
  END la_data_out_mprj[46]
  PIN la_data_out_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 -2.000 673.810 4.000 ;
    END
  END la_data_out_mprj[47]
  PIN la_data_out_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 -2.000 686.690 4.000 ;
    END
  END la_data_out_mprj[48]
  PIN la_data_out_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 -2.000 699.570 4.000 ;
    END
  END la_data_out_mprj[49]
  PIN la_data_out_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 -2.000 119.970 4.000 ;
    END
  END la_data_out_mprj[4]
  PIN la_data_out_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 -2.000 712.450 4.000 ;
    END
  END la_data_out_mprj[50]
  PIN la_data_out_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 -2.000 725.330 4.000 ;
    END
  END la_data_out_mprj[51]
  PIN la_data_out_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 -2.000 738.210 4.000 ;
    END
  END la_data_out_mprj[52]
  PIN la_data_out_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 -2.000 751.090 4.000 ;
    END
  END la_data_out_mprj[53]
  PIN la_data_out_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 -2.000 763.970 4.000 ;
    END
  END la_data_out_mprj[54]
  PIN la_data_out_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 -2.000 776.850 4.000 ;
    END
  END la_data_out_mprj[55]
  PIN la_data_out_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 -2.000 789.730 4.000 ;
    END
  END la_data_out_mprj[56]
  PIN la_data_out_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 -2.000 802.610 4.000 ;
    END
  END la_data_out_mprj[57]
  PIN la_data_out_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 -2.000 815.490 4.000 ;
    END
  END la_data_out_mprj[58]
  PIN la_data_out_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 -2.000 828.370 4.000 ;
    END
  END la_data_out_mprj[59]
  PIN la_data_out_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 -2.000 132.850 4.000 ;
    END
  END la_data_out_mprj[5]
  PIN la_data_out_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 -2.000 841.250 4.000 ;
    END
  END la_data_out_mprj[60]
  PIN la_data_out_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 -2.000 854.130 4.000 ;
    END
  END la_data_out_mprj[61]
  PIN la_data_out_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 -2.000 867.010 4.000 ;
    END
  END la_data_out_mprj[62]
  PIN la_data_out_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 -2.000 879.890 4.000 ;
    END
  END la_data_out_mprj[63]
  PIN la_data_out_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 -2.000 892.770 4.000 ;
    END
  END la_data_out_mprj[64]
  PIN la_data_out_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 -2.000 905.650 4.000 ;
    END
  END la_data_out_mprj[65]
  PIN la_data_out_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 -2.000 918.530 4.000 ;
    END
  END la_data_out_mprj[66]
  PIN la_data_out_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 -2.000 931.410 4.000 ;
    END
  END la_data_out_mprj[67]
  PIN la_data_out_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 -2.000 944.290 4.000 ;
    END
  END la_data_out_mprj[68]
  PIN la_data_out_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 -2.000 957.170 4.000 ;
    END
  END la_data_out_mprj[69]
  PIN la_data_out_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 -2.000 145.730 4.000 ;
    END
  END la_data_out_mprj[6]
  PIN la_data_out_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 -2.000 970.050 4.000 ;
    END
  END la_data_out_mprj[70]
  PIN la_data_out_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 -2.000 989.370 4.000 ;
    END
  END la_data_out_mprj[71]
  PIN la_data_out_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 -2.000 1002.250 4.000 ;
    END
  END la_data_out_mprj[72]
  PIN la_data_out_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 -2.000 1015.130 4.000 ;
    END
  END la_data_out_mprj[73]
  PIN la_data_out_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.730 -2.000 1028.010 4.000 ;
    END
  END la_data_out_mprj[74]
  PIN la_data_out_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 -2.000 1040.890 4.000 ;
    END
  END la_data_out_mprj[75]
  PIN la_data_out_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.490 -2.000 1053.770 4.000 ;
    END
  END la_data_out_mprj[76]
  PIN la_data_out_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 -2.000 1066.650 4.000 ;
    END
  END la_data_out_mprj[77]
  PIN la_data_out_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 -2.000 1079.530 4.000 ;
    END
  END la_data_out_mprj[78]
  PIN la_data_out_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 -2.000 1092.410 4.000 ;
    END
  END la_data_out_mprj[79]
  PIN la_data_out_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 -2.000 158.610 4.000 ;
    END
  END la_data_out_mprj[7]
  PIN la_data_out_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.010 -2.000 1105.290 4.000 ;
    END
  END la_data_out_mprj[80]
  PIN la_data_out_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 -2.000 1118.170 4.000 ;
    END
  END la_data_out_mprj[81]
  PIN la_data_out_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.770 -2.000 1131.050 4.000 ;
    END
  END la_data_out_mprj[82]
  PIN la_data_out_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 -2.000 1143.930 4.000 ;
    END
  END la_data_out_mprj[83]
  PIN la_data_out_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.530 -2.000 1156.810 4.000 ;
    END
  END la_data_out_mprj[84]
  PIN la_data_out_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 -2.000 1169.690 4.000 ;
    END
  END la_data_out_mprj[85]
  PIN la_data_out_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 -2.000 1182.570 4.000 ;
    END
  END la_data_out_mprj[86]
  PIN la_data_out_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 -2.000 1195.450 4.000 ;
    END
  END la_data_out_mprj[87]
  PIN la_data_out_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.050 -2.000 1208.330 4.000 ;
    END
  END la_data_out_mprj[88]
  PIN la_data_out_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.930 -2.000 1221.210 4.000 ;
    END
  END la_data_out_mprj[89]
  PIN la_data_out_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 -2.000 171.490 4.000 ;
    END
  END la_data_out_mprj[8]
  PIN la_data_out_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 -2.000 1234.090 4.000 ;
    END
  END la_data_out_mprj[90]
  PIN la_data_out_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 -2.000 1246.970 4.000 ;
    END
  END la_data_out_mprj[91]
  PIN la_data_out_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.570 -2.000 1259.850 4.000 ;
    END
  END la_data_out_mprj[92]
  PIN la_data_out_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 -2.000 1272.730 4.000 ;
    END
  END la_data_out_mprj[93]
  PIN la_data_out_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 -2.000 1285.610 4.000 ;
    END
  END la_data_out_mprj[94]
  PIN la_data_out_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 -2.000 1298.490 4.000 ;
    END
  END la_data_out_mprj[95]
  PIN la_data_out_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.090 -2.000 1311.370 4.000 ;
    END
  END la_data_out_mprj[96]
  PIN la_data_out_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.970 -2.000 1324.250 4.000 ;
    END
  END la_data_out_mprj[97]
  PIN la_data_out_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 -2.000 1337.130 4.000 ;
    END
  END la_data_out_mprj[98]
  PIN la_data_out_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 -2.000 1350.010 4.000 ;
    END
  END la_data_out_mprj[99]
  PIN la_data_out_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 -2.000 184.370 4.000 ;
    END
  END la_data_out_mprj[9]
  PIN la_iena_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 -2.000 71.670 4.000 ;
    END
  END la_iena_mprj[0]
  PIN la_iena_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.830 -2.000 1366.110 4.000 ;
    END
  END la_iena_mprj[100]
  PIN la_iena_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 -2.000 1378.990 4.000 ;
    END
  END la_iena_mprj[101]
  PIN la_iena_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.590 -2.000 1391.870 4.000 ;
    END
  END la_iena_mprj[102]
  PIN la_iena_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.470 -2.000 1404.750 4.000 ;
    END
  END la_iena_mprj[103]
  PIN la_iena_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 -2.000 1417.630 4.000 ;
    END
  END la_iena_mprj[104]
  PIN la_iena_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.230 -2.000 1430.510 4.000 ;
    END
  END la_iena_mprj[105]
  PIN la_iena_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 -2.000 1443.390 4.000 ;
    END
  END la_iena_mprj[106]
  PIN la_iena_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 -2.000 1456.270 4.000 ;
    END
  END la_iena_mprj[107]
  PIN la_iena_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.870 -2.000 1469.150 4.000 ;
    END
  END la_iena_mprj[108]
  PIN la_iena_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.750 -2.000 1482.030 4.000 ;
    END
  END la_iena_mprj[109]
  PIN la_iena_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 -2.000 200.470 4.000 ;
    END
  END la_iena_mprj[10]
  PIN la_iena_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.630 -2.000 1494.910 4.000 ;
    END
  END la_iena_mprj[110]
  PIN la_iena_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 -2.000 1507.790 4.000 ;
    END
  END la_iena_mprj[111]
  PIN la_iena_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.390 -2.000 1520.670 4.000 ;
    END
  END la_iena_mprj[112]
  PIN la_iena_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 -2.000 1533.550 4.000 ;
    END
  END la_iena_mprj[113]
  PIN la_iena_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 -2.000 1546.430 4.000 ;
    END
  END la_iena_mprj[114]
  PIN la_iena_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.030 -2.000 1559.310 4.000 ;
    END
  END la_iena_mprj[115]
  PIN la_iena_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 -2.000 1572.190 4.000 ;
    END
  END la_iena_mprj[116]
  PIN la_iena_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 -2.000 1585.070 4.000 ;
    END
  END la_iena_mprj[117]
  PIN la_iena_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 -2.000 1597.950 4.000 ;
    END
  END la_iena_mprj[118]
  PIN la_iena_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.550 -2.000 1610.830 4.000 ;
    END
  END la_iena_mprj[119]
  PIN la_iena_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 -2.000 213.350 4.000 ;
    END
  END la_iena_mprj[11]
  PIN la_iena_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.430 -2.000 1623.710 4.000 ;
    END
  END la_iena_mprj[120]
  PIN la_iena_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.310 -2.000 1636.590 4.000 ;
    END
  END la_iena_mprj[121]
  PIN la_iena_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.190 -2.000 1649.470 4.000 ;
    END
  END la_iena_mprj[122]
  PIN la_iena_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.070 -2.000 1662.350 4.000 ;
    END
  END la_iena_mprj[123]
  PIN la_iena_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.950 -2.000 1675.230 4.000 ;
    END
  END la_iena_mprj[124]
  PIN la_iena_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 -2.000 1688.110 4.000 ;
    END
  END la_iena_mprj[125]
  PIN la_iena_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.710 -2.000 1700.990 4.000 ;
    END
  END la_iena_mprj[126]
  PIN la_iena_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.590 -2.000 1713.870 4.000 ;
    END
  END la_iena_mprj[127]
  PIN la_iena_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 -2.000 226.230 4.000 ;
    END
  END la_iena_mprj[12]
  PIN la_iena_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 -2.000 239.110 4.000 ;
    END
  END la_iena_mprj[13]
  PIN la_iena_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 -2.000 251.990 4.000 ;
    END
  END la_iena_mprj[14]
  PIN la_iena_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 -2.000 264.870 4.000 ;
    END
  END la_iena_mprj[15]
  PIN la_iena_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 -2.000 277.750 4.000 ;
    END
  END la_iena_mprj[16]
  PIN la_iena_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 -2.000 290.630 4.000 ;
    END
  END la_iena_mprj[17]
  PIN la_iena_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 -2.000 303.510 4.000 ;
    END
  END la_iena_mprj[18]
  PIN la_iena_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 -2.000 316.390 4.000 ;
    END
  END la_iena_mprj[19]
  PIN la_iena_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 -2.000 84.550 4.000 ;
    END
  END la_iena_mprj[1]
  PIN la_iena_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 -2.000 329.270 4.000 ;
    END
  END la_iena_mprj[20]
  PIN la_iena_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 -2.000 342.150 4.000 ;
    END
  END la_iena_mprj[21]
  PIN la_iena_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 -2.000 355.030 4.000 ;
    END
  END la_iena_mprj[22]
  PIN la_iena_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 -2.000 367.910 4.000 ;
    END
  END la_iena_mprj[23]
  PIN la_iena_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 -2.000 380.790 4.000 ;
    END
  END la_iena_mprj[24]
  PIN la_iena_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 -2.000 393.670 4.000 ;
    END
  END la_iena_mprj[25]
  PIN la_iena_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 -2.000 406.550 4.000 ;
    END
  END la_iena_mprj[26]
  PIN la_iena_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 -2.000 419.430 4.000 ;
    END
  END la_iena_mprj[27]
  PIN la_iena_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 -2.000 432.310 4.000 ;
    END
  END la_iena_mprj[28]
  PIN la_iena_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 -2.000 445.190 4.000 ;
    END
  END la_iena_mprj[29]
  PIN la_iena_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 -2.000 97.430 4.000 ;
    END
  END la_iena_mprj[2]
  PIN la_iena_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 -2.000 458.070 4.000 ;
    END
  END la_iena_mprj[30]
  PIN la_iena_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 -2.000 470.950 4.000 ;
    END
  END la_iena_mprj[31]
  PIN la_iena_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 -2.000 483.830 4.000 ;
    END
  END la_iena_mprj[32]
  PIN la_iena_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 -2.000 496.710 4.000 ;
    END
  END la_iena_mprj[33]
  PIN la_iena_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 -2.000 509.590 4.000 ;
    END
  END la_iena_mprj[34]
  PIN la_iena_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 -2.000 522.470 4.000 ;
    END
  END la_iena_mprj[35]
  PIN la_iena_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 -2.000 535.350 4.000 ;
    END
  END la_iena_mprj[36]
  PIN la_iena_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 -2.000 548.230 4.000 ;
    END
  END la_iena_mprj[37]
  PIN la_iena_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 -2.000 561.110 4.000 ;
    END
  END la_iena_mprj[38]
  PIN la_iena_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 -2.000 573.990 4.000 ;
    END
  END la_iena_mprj[39]
  PIN la_iena_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 -2.000 110.310 4.000 ;
    END
  END la_iena_mprj[3]
  PIN la_iena_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 -2.000 586.870 4.000 ;
    END
  END la_iena_mprj[40]
  PIN la_iena_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 -2.000 599.750 4.000 ;
    END
  END la_iena_mprj[41]
  PIN la_iena_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 -2.000 612.630 4.000 ;
    END
  END la_iena_mprj[42]
  PIN la_iena_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 -2.000 625.510 4.000 ;
    END
  END la_iena_mprj[43]
  PIN la_iena_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 -2.000 638.390 4.000 ;
    END
  END la_iena_mprj[44]
  PIN la_iena_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 -2.000 651.270 4.000 ;
    END
  END la_iena_mprj[45]
  PIN la_iena_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 -2.000 664.150 4.000 ;
    END
  END la_iena_mprj[46]
  PIN la_iena_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 -2.000 677.030 4.000 ;
    END
  END la_iena_mprj[47]
  PIN la_iena_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 -2.000 689.910 4.000 ;
    END
  END la_iena_mprj[48]
  PIN la_iena_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 -2.000 702.790 4.000 ;
    END
  END la_iena_mprj[49]
  PIN la_iena_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 -2.000 123.190 4.000 ;
    END
  END la_iena_mprj[4]
  PIN la_iena_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 -2.000 715.670 4.000 ;
    END
  END la_iena_mprj[50]
  PIN la_iena_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 -2.000 728.550 4.000 ;
    END
  END la_iena_mprj[51]
  PIN la_iena_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 -2.000 741.430 4.000 ;
    END
  END la_iena_mprj[52]
  PIN la_iena_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 -2.000 754.310 4.000 ;
    END
  END la_iena_mprj[53]
  PIN la_iena_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 -2.000 767.190 4.000 ;
    END
  END la_iena_mprj[54]
  PIN la_iena_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 -2.000 780.070 4.000 ;
    END
  END la_iena_mprj[55]
  PIN la_iena_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 -2.000 792.950 4.000 ;
    END
  END la_iena_mprj[56]
  PIN la_iena_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 -2.000 805.830 4.000 ;
    END
  END la_iena_mprj[57]
  PIN la_iena_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 -2.000 818.710 4.000 ;
    END
  END la_iena_mprj[58]
  PIN la_iena_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 -2.000 831.590 4.000 ;
    END
  END la_iena_mprj[59]
  PIN la_iena_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 -2.000 136.070 4.000 ;
    END
  END la_iena_mprj[5]
  PIN la_iena_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 -2.000 844.470 4.000 ;
    END
  END la_iena_mprj[60]
  PIN la_iena_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 -2.000 857.350 4.000 ;
    END
  END la_iena_mprj[61]
  PIN la_iena_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 -2.000 870.230 4.000 ;
    END
  END la_iena_mprj[62]
  PIN la_iena_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 -2.000 883.110 4.000 ;
    END
  END la_iena_mprj[63]
  PIN la_iena_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 -2.000 895.990 4.000 ;
    END
  END la_iena_mprj[64]
  PIN la_iena_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 -2.000 908.870 4.000 ;
    END
  END la_iena_mprj[65]
  PIN la_iena_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 -2.000 921.750 4.000 ;
    END
  END la_iena_mprj[66]
  PIN la_iena_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 -2.000 934.630 4.000 ;
    END
  END la_iena_mprj[67]
  PIN la_iena_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 -2.000 947.510 4.000 ;
    END
  END la_iena_mprj[68]
  PIN la_iena_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 -2.000 960.390 4.000 ;
    END
  END la_iena_mprj[69]
  PIN la_iena_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 -2.000 148.950 4.000 ;
    END
  END la_iena_mprj[6]
  PIN la_iena_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 -2.000 973.270 4.000 ;
    END
  END la_iena_mprj[70]
  PIN la_iena_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 -2.000 992.590 4.000 ;
    END
  END la_iena_mprj[71]
  PIN la_iena_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 -2.000 1005.470 4.000 ;
    END
  END la_iena_mprj[72]
  PIN la_iena_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 -2.000 1018.350 4.000 ;
    END
  END la_iena_mprj[73]
  PIN la_iena_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 -2.000 1031.230 4.000 ;
    END
  END la_iena_mprj[74]
  PIN la_iena_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.830 -2.000 1044.110 4.000 ;
    END
  END la_iena_mprj[75]
  PIN la_iena_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 -2.000 1056.990 4.000 ;
    END
  END la_iena_mprj[76]
  PIN la_iena_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 -2.000 1069.870 4.000 ;
    END
  END la_iena_mprj[77]
  PIN la_iena_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.470 -2.000 1082.750 4.000 ;
    END
  END la_iena_mprj[78]
  PIN la_iena_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 -2.000 1095.630 4.000 ;
    END
  END la_iena_mprj[79]
  PIN la_iena_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 -2.000 161.830 4.000 ;
    END
  END la_iena_mprj[7]
  PIN la_iena_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 -2.000 1108.510 4.000 ;
    END
  END la_iena_mprj[80]
  PIN la_iena_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 -2.000 1121.390 4.000 ;
    END
  END la_iena_mprj[81]
  PIN la_iena_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 -2.000 1134.270 4.000 ;
    END
  END la_iena_mprj[82]
  PIN la_iena_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 -2.000 1147.150 4.000 ;
    END
  END la_iena_mprj[83]
  PIN la_iena_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.750 -2.000 1160.030 4.000 ;
    END
  END la_iena_mprj[84]
  PIN la_iena_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 -2.000 1172.910 4.000 ;
    END
  END la_iena_mprj[85]
  PIN la_iena_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 -2.000 1185.790 4.000 ;
    END
  END la_iena_mprj[86]
  PIN la_iena_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 -2.000 1198.670 4.000 ;
    END
  END la_iena_mprj[87]
  PIN la_iena_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.270 -2.000 1211.550 4.000 ;
    END
  END la_iena_mprj[88]
  PIN la_iena_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 -2.000 1224.430 4.000 ;
    END
  END la_iena_mprj[89]
  PIN la_iena_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 -2.000 174.710 4.000 ;
    END
  END la_iena_mprj[8]
  PIN la_iena_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 -2.000 1237.310 4.000 ;
    END
  END la_iena_mprj[90]
  PIN la_iena_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 -2.000 1250.190 4.000 ;
    END
  END la_iena_mprj[91]
  PIN la_iena_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 -2.000 1263.070 4.000 ;
    END
  END la_iena_mprj[92]
  PIN la_iena_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 -2.000 1275.950 4.000 ;
    END
  END la_iena_mprj[93]
  PIN la_iena_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.550 -2.000 1288.830 4.000 ;
    END
  END la_iena_mprj[94]
  PIN la_iena_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 -2.000 1301.710 4.000 ;
    END
  END la_iena_mprj[95]
  PIN la_iena_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 -2.000 1314.590 4.000 ;
    END
  END la_iena_mprj[96]
  PIN la_iena_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 -2.000 1327.470 4.000 ;
    END
  END la_iena_mprj[97]
  PIN la_iena_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 -2.000 1340.350 4.000 ;
    END
  END la_iena_mprj[98]
  PIN la_iena_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 -2.000 1353.230 4.000 ;
    END
  END la_iena_mprj[99]
  PIN la_iena_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 -2.000 187.590 4.000 ;
    END
  END la_iena_mprj[9]
  PIN la_oenb_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 156.000 493.030 162.000 ;
    END
  END la_oenb_core[0]
  PIN la_oenb_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.750 156.000 1735.030 162.000 ;
    END
  END la_oenb_core[100]
  PIN la_oenb_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 156.000 1747.450 162.000 ;
    END
  END la_oenb_core[101]
  PIN la_oenb_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1759.590 156.000 1759.870 162.000 ;
    END
  END la_oenb_core[102]
  PIN la_oenb_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.010 156.000 1772.290 162.000 ;
    END
  END la_oenb_core[103]
  PIN la_oenb_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.430 156.000 1784.710 162.000 ;
    END
  END la_oenb_core[104]
  PIN la_oenb_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 156.000 1797.130 162.000 ;
    END
  END la_oenb_core[105]
  PIN la_oenb_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.270 156.000 1809.550 162.000 ;
    END
  END la_oenb_core[106]
  PIN la_oenb_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.690 156.000 1821.970 162.000 ;
    END
  END la_oenb_core[107]
  PIN la_oenb_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.110 156.000 1834.390 162.000 ;
    END
  END la_oenb_core[108]
  PIN la_oenb_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.530 156.000 1846.810 162.000 ;
    END
  END la_oenb_core[109]
  PIN la_oenb_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 156.000 617.230 162.000 ;
    END
  END la_oenb_core[10]
  PIN la_oenb_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.950 156.000 1859.230 162.000 ;
    END
  END la_oenb_core[110]
  PIN la_oenb_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.370 156.000 1871.650 162.000 ;
    END
  END la_oenb_core[111]
  PIN la_oenb_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.790 156.000 1884.070 162.000 ;
    END
  END la_oenb_core[112]
  PIN la_oenb_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.210 156.000 1896.490 162.000 ;
    END
  END la_oenb_core[113]
  PIN la_oenb_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.630 156.000 1908.910 162.000 ;
    END
  END la_oenb_core[114]
  PIN la_oenb_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.050 156.000 1921.330 162.000 ;
    END
  END la_oenb_core[115]
  PIN la_oenb_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.470 156.000 1933.750 162.000 ;
    END
  END la_oenb_core[116]
  PIN la_oenb_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.890 156.000 1946.170 162.000 ;
    END
  END la_oenb_core[117]
  PIN la_oenb_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.310 156.000 1958.590 162.000 ;
    END
  END la_oenb_core[118]
  PIN la_oenb_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.730 156.000 1971.010 162.000 ;
    END
  END la_oenb_core[119]
  PIN la_oenb_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 156.000 629.650 162.000 ;
    END
  END la_oenb_core[11]
  PIN la_oenb_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.150 156.000 1983.430 162.000 ;
    END
  END la_oenb_core[120]
  PIN la_oenb_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.570 156.000 1995.850 162.000 ;
    END
  END la_oenb_core[121]
  PIN la_oenb_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2007.990 156.000 2008.270 162.000 ;
    END
  END la_oenb_core[122]
  PIN la_oenb_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2020.410 156.000 2020.690 162.000 ;
    END
  END la_oenb_core[123]
  PIN la_oenb_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2032.830 156.000 2033.110 162.000 ;
    END
  END la_oenb_core[124]
  PIN la_oenb_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.250 156.000 2045.530 162.000 ;
    END
  END la_oenb_core[125]
  PIN la_oenb_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.670 156.000 2057.950 162.000 ;
    END
  END la_oenb_core[126]
  PIN la_oenb_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.090 156.000 2070.370 162.000 ;
    END
  END la_oenb_core[127]
  PIN la_oenb_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 156.000 642.070 162.000 ;
    END
  END la_oenb_core[12]
  PIN la_oenb_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 156.000 654.490 162.000 ;
    END
  END la_oenb_core[13]
  PIN la_oenb_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 156.000 666.910 162.000 ;
    END
  END la_oenb_core[14]
  PIN la_oenb_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 156.000 679.330 162.000 ;
    END
  END la_oenb_core[15]
  PIN la_oenb_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 156.000 691.750 162.000 ;
    END
  END la_oenb_core[16]
  PIN la_oenb_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 156.000 704.170 162.000 ;
    END
  END la_oenb_core[17]
  PIN la_oenb_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 156.000 716.590 162.000 ;
    END
  END la_oenb_core[18]
  PIN la_oenb_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 156.000 729.010 162.000 ;
    END
  END la_oenb_core[19]
  PIN la_oenb_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 156.000 505.450 162.000 ;
    END
  END la_oenb_core[1]
  PIN la_oenb_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 156.000 741.430 162.000 ;
    END
  END la_oenb_core[20]
  PIN la_oenb_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 156.000 753.850 162.000 ;
    END
  END la_oenb_core[21]
  PIN la_oenb_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 156.000 766.270 162.000 ;
    END
  END la_oenb_core[22]
  PIN la_oenb_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 156.000 778.690 162.000 ;
    END
  END la_oenb_core[23]
  PIN la_oenb_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 156.000 791.110 162.000 ;
    END
  END la_oenb_core[24]
  PIN la_oenb_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 156.000 803.530 162.000 ;
    END
  END la_oenb_core[25]
  PIN la_oenb_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 156.000 815.950 162.000 ;
    END
  END la_oenb_core[26]
  PIN la_oenb_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 156.000 828.370 162.000 ;
    END
  END la_oenb_core[27]
  PIN la_oenb_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 156.000 840.790 162.000 ;
    END
  END la_oenb_core[28]
  PIN la_oenb_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 156.000 853.210 162.000 ;
    END
  END la_oenb_core[29]
  PIN la_oenb_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 156.000 517.870 162.000 ;
    END
  END la_oenb_core[2]
  PIN la_oenb_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 156.000 865.630 162.000 ;
    END
  END la_oenb_core[30]
  PIN la_oenb_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 156.000 878.050 162.000 ;
    END
  END la_oenb_core[31]
  PIN la_oenb_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 156.000 890.470 162.000 ;
    END
  END la_oenb_core[32]
  PIN la_oenb_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 156.000 902.890 162.000 ;
    END
  END la_oenb_core[33]
  PIN la_oenb_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 156.000 915.310 162.000 ;
    END
  END la_oenb_core[34]
  PIN la_oenb_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 156.000 927.730 162.000 ;
    END
  END la_oenb_core[35]
  PIN la_oenb_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 156.000 940.150 162.000 ;
    END
  END la_oenb_core[36]
  PIN la_oenb_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 156.000 952.570 162.000 ;
    END
  END la_oenb_core[37]
  PIN la_oenb_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 156.000 964.990 162.000 ;
    END
  END la_oenb_core[38]
  PIN la_oenb_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 156.000 977.410 162.000 ;
    END
  END la_oenb_core[39]
  PIN la_oenb_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 156.000 530.290 162.000 ;
    END
  END la_oenb_core[3]
  PIN la_oenb_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 156.000 989.830 162.000 ;
    END
  END la_oenb_core[40]
  PIN la_oenb_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 156.000 1002.250 162.000 ;
    END
  END la_oenb_core[41]
  PIN la_oenb_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 156.000 1014.670 162.000 ;
    END
  END la_oenb_core[42]
  PIN la_oenb_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.810 156.000 1027.090 162.000 ;
    END
  END la_oenb_core[43]
  PIN la_oenb_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.230 156.000 1039.510 162.000 ;
    END
  END la_oenb_core[44]
  PIN la_oenb_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 156.000 1051.930 162.000 ;
    END
  END la_oenb_core[45]
  PIN la_oenb_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.070 156.000 1064.350 162.000 ;
    END
  END la_oenb_core[46]
  PIN la_oenb_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 156.000 1076.770 162.000 ;
    END
  END la_oenb_core[47]
  PIN la_oenb_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 156.000 1089.190 162.000 ;
    END
  END la_oenb_core[48]
  PIN la_oenb_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 156.000 1101.610 162.000 ;
    END
  END la_oenb_core[49]
  PIN la_oenb_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 156.000 542.710 162.000 ;
    END
  END la_oenb_core[4]
  PIN la_oenb_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.750 156.000 1114.030 162.000 ;
    END
  END la_oenb_core[50]
  PIN la_oenb_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.170 156.000 1126.450 162.000 ;
    END
  END la_oenb_core[51]
  PIN la_oenb_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.590 156.000 1138.870 162.000 ;
    END
  END la_oenb_core[52]
  PIN la_oenb_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.010 156.000 1151.290 162.000 ;
    END
  END la_oenb_core[53]
  PIN la_oenb_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.430 156.000 1163.710 162.000 ;
    END
  END la_oenb_core[54]
  PIN la_oenb_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 156.000 1176.130 162.000 ;
    END
  END la_oenb_core[55]
  PIN la_oenb_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 156.000 1188.550 162.000 ;
    END
  END la_oenb_core[56]
  PIN la_oenb_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.690 156.000 1200.970 162.000 ;
    END
  END la_oenb_core[57]
  PIN la_oenb_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 156.000 1213.390 162.000 ;
    END
  END la_oenb_core[58]
  PIN la_oenb_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.530 156.000 1225.810 162.000 ;
    END
  END la_oenb_core[59]
  PIN la_oenb_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 156.000 555.130 162.000 ;
    END
  END la_oenb_core[5]
  PIN la_oenb_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.950 156.000 1238.230 162.000 ;
    END
  END la_oenb_core[60]
  PIN la_oenb_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.370 156.000 1250.650 162.000 ;
    END
  END la_oenb_core[61]
  PIN la_oenb_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 156.000 1263.070 162.000 ;
    END
  END la_oenb_core[62]
  PIN la_oenb_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 156.000 1275.490 162.000 ;
    END
  END la_oenb_core[63]
  PIN la_oenb_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.630 156.000 1287.910 162.000 ;
    END
  END la_oenb_core[64]
  PIN la_oenb_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.050 156.000 1300.330 162.000 ;
    END
  END la_oenb_core[65]
  PIN la_oenb_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.470 156.000 1312.750 162.000 ;
    END
  END la_oenb_core[66]
  PIN la_oenb_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.890 156.000 1325.170 162.000 ;
    END
  END la_oenb_core[67]
  PIN la_oenb_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.310 156.000 1337.590 162.000 ;
    END
  END la_oenb_core[68]
  PIN la_oenb_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 156.000 1350.010 162.000 ;
    END
  END la_oenb_core[69]
  PIN la_oenb_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 156.000 567.550 162.000 ;
    END
  END la_oenb_core[6]
  PIN la_oenb_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 156.000 1362.430 162.000 ;
    END
  END la_oenb_core[70]
  PIN la_oenb_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.570 156.000 1374.850 162.000 ;
    END
  END la_oenb_core[71]
  PIN la_oenb_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 156.000 1387.270 162.000 ;
    END
  END la_oenb_core[72]
  PIN la_oenb_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.410 156.000 1399.690 162.000 ;
    END
  END la_oenb_core[73]
  PIN la_oenb_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 156.000 1412.110 162.000 ;
    END
  END la_oenb_core[74]
  PIN la_oenb_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.250 156.000 1424.530 162.000 ;
    END
  END la_oenb_core[75]
  PIN la_oenb_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.670 156.000 1436.950 162.000 ;
    END
  END la_oenb_core[76]
  PIN la_oenb_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 156.000 1449.370 162.000 ;
    END
  END la_oenb_core[77]
  PIN la_oenb_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.510 156.000 1461.790 162.000 ;
    END
  END la_oenb_core[78]
  PIN la_oenb_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 156.000 1474.210 162.000 ;
    END
  END la_oenb_core[79]
  PIN la_oenb_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 156.000 579.970 162.000 ;
    END
  END la_oenb_core[7]
  PIN la_oenb_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.350 156.000 1486.630 162.000 ;
    END
  END la_oenb_core[80]
  PIN la_oenb_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.770 156.000 1499.050 162.000 ;
    END
  END la_oenb_core[81]
  PIN la_oenb_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.190 156.000 1511.470 162.000 ;
    END
  END la_oenb_core[82]
  PIN la_oenb_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.610 156.000 1523.890 162.000 ;
    END
  END la_oenb_core[83]
  PIN la_oenb_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 156.000 1536.310 162.000 ;
    END
  END la_oenb_core[84]
  PIN la_oenb_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 156.000 1548.730 162.000 ;
    END
  END la_oenb_core[85]
  PIN la_oenb_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.870 156.000 1561.150 162.000 ;
    END
  END la_oenb_core[86]
  PIN la_oenb_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 156.000 1573.570 162.000 ;
    END
  END la_oenb_core[87]
  PIN la_oenb_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.710 156.000 1585.990 162.000 ;
    END
  END la_oenb_core[88]
  PIN la_oenb_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.130 156.000 1598.410 162.000 ;
    END
  END la_oenb_core[89]
  PIN la_oenb_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 156.000 592.390 162.000 ;
    END
  END la_oenb_core[8]
  PIN la_oenb_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.550 156.000 1610.830 162.000 ;
    END
  END la_oenb_core[90]
  PIN la_oenb_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 156.000 1623.250 162.000 ;
    END
  END la_oenb_core[91]
  PIN la_oenb_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.390 156.000 1635.670 162.000 ;
    END
  END la_oenb_core[92]
  PIN la_oenb_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.810 156.000 1648.090 162.000 ;
    END
  END la_oenb_core[93]
  PIN la_oenb_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.230 156.000 1660.510 162.000 ;
    END
  END la_oenb_core[94]
  PIN la_oenb_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.650 156.000 1672.930 162.000 ;
    END
  END la_oenb_core[95]
  PIN la_oenb_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.070 156.000 1685.350 162.000 ;
    END
  END la_oenb_core[96]
  PIN la_oenb_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 156.000 1697.770 162.000 ;
    END
  END la_oenb_core[97]
  PIN la_oenb_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.910 156.000 1710.190 162.000 ;
    END
  END la_oenb_core[98]
  PIN la_oenb_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 156.000 1722.610 162.000 ;
    END
  END la_oenb_core[99]
  PIN la_oenb_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 156.000 604.810 162.000 ;
    END
  END la_oenb_core[9]
  PIN la_oenb_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 -2.000 74.890 4.000 ;
    END
  END la_oenb_mprj[0]
  PIN la_oenb_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 -2.000 1369.330 4.000 ;
    END
  END la_oenb_mprj[100]
  PIN la_oenb_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 -2.000 1382.210 4.000 ;
    END
  END la_oenb_mprj[101]
  PIN la_oenb_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 -2.000 1395.090 4.000 ;
    END
  END la_oenb_mprj[102]
  PIN la_oenb_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 -2.000 1407.970 4.000 ;
    END
  END la_oenb_mprj[103]
  PIN la_oenb_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.570 -2.000 1420.850 4.000 ;
    END
  END la_oenb_mprj[104]
  PIN la_oenb_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 -2.000 1433.730 4.000 ;
    END
  END la_oenb_mprj[105]
  PIN la_oenb_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 -2.000 1446.610 4.000 ;
    END
  END la_oenb_mprj[106]
  PIN la_oenb_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.210 -2.000 1459.490 4.000 ;
    END
  END la_oenb_mprj[107]
  PIN la_oenb_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.090 -2.000 1472.370 4.000 ;
    END
  END la_oenb_mprj[108]
  PIN la_oenb_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 -2.000 1485.250 4.000 ;
    END
  END la_oenb_mprj[109]
  PIN la_oenb_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 -2.000 203.690 4.000 ;
    END
  END la_oenb_mprj[10]
  PIN la_oenb_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.850 -2.000 1498.130 4.000 ;
    END
  END la_oenb_mprj[110]
  PIN la_oenb_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 -2.000 1511.010 4.000 ;
    END
  END la_oenb_mprj[111]
  PIN la_oenb_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.610 -2.000 1523.890 4.000 ;
    END
  END la_oenb_mprj[112]
  PIN la_oenb_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.490 -2.000 1536.770 4.000 ;
    END
  END la_oenb_mprj[113]
  PIN la_oenb_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.370 -2.000 1549.650 4.000 ;
    END
  END la_oenb_mprj[114]
  PIN la_oenb_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.250 -2.000 1562.530 4.000 ;
    END
  END la_oenb_mprj[115]
  PIN la_oenb_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 -2.000 1575.410 4.000 ;
    END
  END la_oenb_mprj[116]
  PIN la_oenb_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.010 -2.000 1588.290 4.000 ;
    END
  END la_oenb_mprj[117]
  PIN la_oenb_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 -2.000 1601.170 4.000 ;
    END
  END la_oenb_mprj[118]
  PIN la_oenb_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.770 -2.000 1614.050 4.000 ;
    END
  END la_oenb_mprj[119]
  PIN la_oenb_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 -2.000 216.570 4.000 ;
    END
  END la_oenb_mprj[11]
  PIN la_oenb_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.650 -2.000 1626.930 4.000 ;
    END
  END la_oenb_mprj[120]
  PIN la_oenb_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 -2.000 1639.810 4.000 ;
    END
  END la_oenb_mprj[121]
  PIN la_oenb_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.410 -2.000 1652.690 4.000 ;
    END
  END la_oenb_mprj[122]
  PIN la_oenb_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.290 -2.000 1665.570 4.000 ;
    END
  END la_oenb_mprj[123]
  PIN la_oenb_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.170 -2.000 1678.450 4.000 ;
    END
  END la_oenb_mprj[124]
  PIN la_oenb_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.050 -2.000 1691.330 4.000 ;
    END
  END la_oenb_mprj[125]
  PIN la_oenb_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.930 -2.000 1704.210 4.000 ;
    END
  END la_oenb_mprj[126]
  PIN la_oenb_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 -2.000 1717.090 4.000 ;
    END
  END la_oenb_mprj[127]
  PIN la_oenb_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 -2.000 229.450 4.000 ;
    END
  END la_oenb_mprj[12]
  PIN la_oenb_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 -2.000 242.330 4.000 ;
    END
  END la_oenb_mprj[13]
  PIN la_oenb_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 -2.000 255.210 4.000 ;
    END
  END la_oenb_mprj[14]
  PIN la_oenb_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 -2.000 268.090 4.000 ;
    END
  END la_oenb_mprj[15]
  PIN la_oenb_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 -2.000 280.970 4.000 ;
    END
  END la_oenb_mprj[16]
  PIN la_oenb_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 -2.000 293.850 4.000 ;
    END
  END la_oenb_mprj[17]
  PIN la_oenb_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 -2.000 306.730 4.000 ;
    END
  END la_oenb_mprj[18]
  PIN la_oenb_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 -2.000 319.610 4.000 ;
    END
  END la_oenb_mprj[19]
  PIN la_oenb_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 -2.000 87.770 4.000 ;
    END
  END la_oenb_mprj[1]
  PIN la_oenb_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 -2.000 332.490 4.000 ;
    END
  END la_oenb_mprj[20]
  PIN la_oenb_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 -2.000 345.370 4.000 ;
    END
  END la_oenb_mprj[21]
  PIN la_oenb_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 -2.000 358.250 4.000 ;
    END
  END la_oenb_mprj[22]
  PIN la_oenb_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 -2.000 371.130 4.000 ;
    END
  END la_oenb_mprj[23]
  PIN la_oenb_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 -2.000 384.010 4.000 ;
    END
  END la_oenb_mprj[24]
  PIN la_oenb_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 -2.000 396.890 4.000 ;
    END
  END la_oenb_mprj[25]
  PIN la_oenb_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 -2.000 409.770 4.000 ;
    END
  END la_oenb_mprj[26]
  PIN la_oenb_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 -2.000 422.650 4.000 ;
    END
  END la_oenb_mprj[27]
  PIN la_oenb_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 -2.000 435.530 4.000 ;
    END
  END la_oenb_mprj[28]
  PIN la_oenb_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 -2.000 448.410 4.000 ;
    END
  END la_oenb_mprj[29]
  PIN la_oenb_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 -2.000 100.650 4.000 ;
    END
  END la_oenb_mprj[2]
  PIN la_oenb_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 -2.000 461.290 4.000 ;
    END
  END la_oenb_mprj[30]
  PIN la_oenb_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 -2.000 474.170 4.000 ;
    END
  END la_oenb_mprj[31]
  PIN la_oenb_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 -2.000 487.050 4.000 ;
    END
  END la_oenb_mprj[32]
  PIN la_oenb_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 -2.000 499.930 4.000 ;
    END
  END la_oenb_mprj[33]
  PIN la_oenb_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 -2.000 512.810 4.000 ;
    END
  END la_oenb_mprj[34]
  PIN la_oenb_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 -2.000 525.690 4.000 ;
    END
  END la_oenb_mprj[35]
  PIN la_oenb_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 -2.000 538.570 4.000 ;
    END
  END la_oenb_mprj[36]
  PIN la_oenb_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 -2.000 551.450 4.000 ;
    END
  END la_oenb_mprj[37]
  PIN la_oenb_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 -2.000 564.330 4.000 ;
    END
  END la_oenb_mprj[38]
  PIN la_oenb_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 -2.000 577.210 4.000 ;
    END
  END la_oenb_mprj[39]
  PIN la_oenb_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 -2.000 113.530 4.000 ;
    END
  END la_oenb_mprj[3]
  PIN la_oenb_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 -2.000 590.090 4.000 ;
    END
  END la_oenb_mprj[40]
  PIN la_oenb_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 -2.000 602.970 4.000 ;
    END
  END la_oenb_mprj[41]
  PIN la_oenb_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 -2.000 615.850 4.000 ;
    END
  END la_oenb_mprj[42]
  PIN la_oenb_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 -2.000 628.730 4.000 ;
    END
  END la_oenb_mprj[43]
  PIN la_oenb_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 -2.000 641.610 4.000 ;
    END
  END la_oenb_mprj[44]
  PIN la_oenb_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 -2.000 654.490 4.000 ;
    END
  END la_oenb_mprj[45]
  PIN la_oenb_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 -2.000 667.370 4.000 ;
    END
  END la_oenb_mprj[46]
  PIN la_oenb_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 -2.000 680.250 4.000 ;
    END
  END la_oenb_mprj[47]
  PIN la_oenb_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 -2.000 693.130 4.000 ;
    END
  END la_oenb_mprj[48]
  PIN la_oenb_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 -2.000 706.010 4.000 ;
    END
  END la_oenb_mprj[49]
  PIN la_oenb_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 -2.000 126.410 4.000 ;
    END
  END la_oenb_mprj[4]
  PIN la_oenb_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 -2.000 718.890 4.000 ;
    END
  END la_oenb_mprj[50]
  PIN la_oenb_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 -2.000 731.770 4.000 ;
    END
  END la_oenb_mprj[51]
  PIN la_oenb_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 -2.000 744.650 4.000 ;
    END
  END la_oenb_mprj[52]
  PIN la_oenb_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 -2.000 757.530 4.000 ;
    END
  END la_oenb_mprj[53]
  PIN la_oenb_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 -2.000 770.410 4.000 ;
    END
  END la_oenb_mprj[54]
  PIN la_oenb_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 -2.000 783.290 4.000 ;
    END
  END la_oenb_mprj[55]
  PIN la_oenb_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 -2.000 796.170 4.000 ;
    END
  END la_oenb_mprj[56]
  PIN la_oenb_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 -2.000 809.050 4.000 ;
    END
  END la_oenb_mprj[57]
  PIN la_oenb_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 -2.000 821.930 4.000 ;
    END
  END la_oenb_mprj[58]
  PIN la_oenb_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 -2.000 834.810 4.000 ;
    END
  END la_oenb_mprj[59]
  PIN la_oenb_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 -2.000 139.290 4.000 ;
    END
  END la_oenb_mprj[5]
  PIN la_oenb_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 -2.000 847.690 4.000 ;
    END
  END la_oenb_mprj[60]
  PIN la_oenb_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 -2.000 860.570 4.000 ;
    END
  END la_oenb_mprj[61]
  PIN la_oenb_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 -2.000 873.450 4.000 ;
    END
  END la_oenb_mprj[62]
  PIN la_oenb_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 -2.000 886.330 4.000 ;
    END
  END la_oenb_mprj[63]
  PIN la_oenb_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 -2.000 899.210 4.000 ;
    END
  END la_oenb_mprj[64]
  PIN la_oenb_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 -2.000 912.090 4.000 ;
    END
  END la_oenb_mprj[65]
  PIN la_oenb_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 -2.000 924.970 4.000 ;
    END
  END la_oenb_mprj[66]
  PIN la_oenb_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 -2.000 937.850 4.000 ;
    END
  END la_oenb_mprj[67]
  PIN la_oenb_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 -2.000 950.730 4.000 ;
    END
  END la_oenb_mprj[68]
  PIN la_oenb_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 -2.000 963.610 4.000 ;
    END
  END la_oenb_mprj[69]
  PIN la_oenb_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 -2.000 152.170 4.000 ;
    END
  END la_oenb_mprj[6]
  PIN la_oenb_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 -2.000 976.490 4.000 ;
    END
  END la_oenb_mprj[70]
  PIN la_oenb_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.530 -2.000 995.810 4.000 ;
    END
  END la_oenb_mprj[71]
  PIN la_oenb_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 -2.000 1008.690 4.000 ;
    END
  END la_oenb_mprj[72]
  PIN la_oenb_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 -2.000 1021.570 4.000 ;
    END
  END la_oenb_mprj[73]
  PIN la_oenb_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 -2.000 1034.450 4.000 ;
    END
  END la_oenb_mprj[74]
  PIN la_oenb_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 -2.000 1047.330 4.000 ;
    END
  END la_oenb_mprj[75]
  PIN la_oenb_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 -2.000 1060.210 4.000 ;
    END
  END la_oenb_mprj[76]
  PIN la_oenb_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.810 -2.000 1073.090 4.000 ;
    END
  END la_oenb_mprj[77]
  PIN la_oenb_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 -2.000 1085.970 4.000 ;
    END
  END la_oenb_mprj[78]
  PIN la_oenb_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 -2.000 1098.850 4.000 ;
    END
  END la_oenb_mprj[79]
  PIN la_oenb_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 -2.000 165.050 4.000 ;
    END
  END la_oenb_mprj[7]
  PIN la_oenb_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.450 -2.000 1111.730 4.000 ;
    END
  END la_oenb_mprj[80]
  PIN la_oenb_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 -2.000 1124.610 4.000 ;
    END
  END la_oenb_mprj[81]
  PIN la_oenb_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 -2.000 1137.490 4.000 ;
    END
  END la_oenb_mprj[82]
  PIN la_oenb_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 -2.000 1150.370 4.000 ;
    END
  END la_oenb_mprj[83]
  PIN la_oenb_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.970 -2.000 1163.250 4.000 ;
    END
  END la_oenb_mprj[84]
  PIN la_oenb_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 -2.000 1176.130 4.000 ;
    END
  END la_oenb_mprj[85]
  PIN la_oenb_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.730 -2.000 1189.010 4.000 ;
    END
  END la_oenb_mprj[86]
  PIN la_oenb_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.610 -2.000 1201.890 4.000 ;
    END
  END la_oenb_mprj[87]
  PIN la_oenb_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 -2.000 1214.770 4.000 ;
    END
  END la_oenb_mprj[88]
  PIN la_oenb_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 -2.000 1227.650 4.000 ;
    END
  END la_oenb_mprj[89]
  PIN la_oenb_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 -2.000 177.930 4.000 ;
    END
  END la_oenb_mprj[8]
  PIN la_oenb_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.250 -2.000 1240.530 4.000 ;
    END
  END la_oenb_mprj[90]
  PIN la_oenb_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 -2.000 1253.410 4.000 ;
    END
  END la_oenb_mprj[91]
  PIN la_oenb_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 -2.000 1266.290 4.000 ;
    END
  END la_oenb_mprj[92]
  PIN la_oenb_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 -2.000 1279.170 4.000 ;
    END
  END la_oenb_mprj[93]
  PIN la_oenb_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 -2.000 1292.050 4.000 ;
    END
  END la_oenb_mprj[94]
  PIN la_oenb_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.650 -2.000 1304.930 4.000 ;
    END
  END la_oenb_mprj[95]
  PIN la_oenb_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.530 -2.000 1317.810 4.000 ;
    END
  END la_oenb_mprj[96]
  PIN la_oenb_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 -2.000 1330.690 4.000 ;
    END
  END la_oenb_mprj[97]
  PIN la_oenb_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.290 -2.000 1343.570 4.000 ;
    END
  END la_oenb_mprj[98]
  PIN la_oenb_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 -2.000 1356.450 4.000 ;
    END
  END la_oenb_mprj[99]
  PIN la_oenb_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 -2.000 190.810 4.000 ;
    END
  END la_oenb_mprj[9]
  PIN mprj_ack_i_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.030 -2.000 1720.310 4.000 ;
    END
  END mprj_ack_i_core
  PIN mprj_ack_i_user
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 156.000 54.190 162.000 ;
    END
  END mprj_ack_i_user
  PIN mprj_adr_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 -2.000 1733.190 4.000 ;
    END
  END mprj_adr_o_core[0]
  PIN mprj_adr_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.390 -2.000 1842.670 4.000 ;
    END
  END mprj_adr_o_core[10]
  PIN mprj_adr_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.050 -2.000 1852.330 4.000 ;
    END
  END mprj_adr_o_core[11]
  PIN mprj_adr_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 -2.000 1861.990 4.000 ;
    END
  END mprj_adr_o_core[12]
  PIN mprj_adr_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.370 -2.000 1871.650 4.000 ;
    END
  END mprj_adr_o_core[13]
  PIN mprj_adr_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.030 -2.000 1881.310 4.000 ;
    END
  END mprj_adr_o_core[14]
  PIN mprj_adr_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.690 -2.000 1890.970 4.000 ;
    END
  END mprj_adr_o_core[15]
  PIN mprj_adr_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.350 -2.000 1900.630 4.000 ;
    END
  END mprj_adr_o_core[16]
  PIN mprj_adr_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.010 -2.000 1910.290 4.000 ;
    END
  END mprj_adr_o_core[17]
  PIN mprj_adr_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.670 -2.000 1919.950 4.000 ;
    END
  END mprj_adr_o_core[18]
  PIN mprj_adr_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.330 -2.000 1929.610 4.000 ;
    END
  END mprj_adr_o_core[19]
  PIN mprj_adr_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.790 -2.000 1746.070 4.000 ;
    END
  END mprj_adr_o_core[1]
  PIN mprj_adr_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.990 -2.000 1939.270 4.000 ;
    END
  END mprj_adr_o_core[20]
  PIN mprj_adr_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.650 -2.000 1948.930 4.000 ;
    END
  END mprj_adr_o_core[21]
  PIN mprj_adr_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.310 -2.000 1958.590 4.000 ;
    END
  END mprj_adr_o_core[22]
  PIN mprj_adr_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.970 -2.000 1968.250 4.000 ;
    END
  END mprj_adr_o_core[23]
  PIN mprj_adr_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.630 -2.000 1977.910 4.000 ;
    END
  END mprj_adr_o_core[24]
  PIN mprj_adr_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.290 -2.000 1987.570 4.000 ;
    END
  END mprj_adr_o_core[25]
  PIN mprj_adr_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.950 -2.000 1997.230 4.000 ;
    END
  END mprj_adr_o_core[26]
  PIN mprj_adr_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.610 -2.000 2006.890 4.000 ;
    END
  END mprj_adr_o_core[27]
  PIN mprj_adr_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2016.270 -2.000 2016.550 4.000 ;
    END
  END mprj_adr_o_core[28]
  PIN mprj_adr_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.930 -2.000 2026.210 4.000 ;
    END
  END mprj_adr_o_core[29]
  PIN mprj_adr_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.670 -2.000 1758.950 4.000 ;
    END
  END mprj_adr_o_core[2]
  PIN mprj_adr_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.590 -2.000 2035.870 4.000 ;
    END
  END mprj_adr_o_core[30]
  PIN mprj_adr_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.250 -2.000 2045.530 4.000 ;
    END
  END mprj_adr_o_core[31]
  PIN mprj_adr_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.550 -2.000 1771.830 4.000 ;
    END
  END mprj_adr_o_core[3]
  PIN mprj_adr_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.430 -2.000 1784.710 4.000 ;
    END
  END mprj_adr_o_core[4]
  PIN mprj_adr_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.090 -2.000 1794.370 4.000 ;
    END
  END mprj_adr_o_core[5]
  PIN mprj_adr_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.750 -2.000 1804.030 4.000 ;
    END
  END mprj_adr_o_core[6]
  PIN mprj_adr_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.410 -2.000 1813.690 4.000 ;
    END
  END mprj_adr_o_core[7]
  PIN mprj_adr_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.070 -2.000 1823.350 4.000 ;
    END
  END mprj_adr_o_core[8]
  PIN mprj_adr_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.730 -2.000 1833.010 4.000 ;
    END
  END mprj_adr_o_core[9]
  PIN mprj_adr_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 156.000 70.750 162.000 ;
    END
  END mprj_adr_o_user[0]
  PIN mprj_adr_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 156.000 211.510 162.000 ;
    END
  END mprj_adr_o_user[10]
  PIN mprj_adr_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 156.000 223.930 162.000 ;
    END
  END mprj_adr_o_user[11]
  PIN mprj_adr_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 156.000 236.350 162.000 ;
    END
  END mprj_adr_o_user[12]
  PIN mprj_adr_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 156.000 248.770 162.000 ;
    END
  END mprj_adr_o_user[13]
  PIN mprj_adr_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 156.000 261.190 162.000 ;
    END
  END mprj_adr_o_user[14]
  PIN mprj_adr_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 156.000 273.610 162.000 ;
    END
  END mprj_adr_o_user[15]
  PIN mprj_adr_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 156.000 286.030 162.000 ;
    END
  END mprj_adr_o_user[16]
  PIN mprj_adr_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 156.000 298.450 162.000 ;
    END
  END mprj_adr_o_user[17]
  PIN mprj_adr_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 156.000 310.870 162.000 ;
    END
  END mprj_adr_o_user[18]
  PIN mprj_adr_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 156.000 323.290 162.000 ;
    END
  END mprj_adr_o_user[19]
  PIN mprj_adr_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 156.000 87.310 162.000 ;
    END
  END mprj_adr_o_user[1]
  PIN mprj_adr_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 156.000 335.710 162.000 ;
    END
  END mprj_adr_o_user[20]
  PIN mprj_adr_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 156.000 348.130 162.000 ;
    END
  END mprj_adr_o_user[21]
  PIN mprj_adr_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 156.000 360.550 162.000 ;
    END
  END mprj_adr_o_user[22]
  PIN mprj_adr_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 156.000 372.970 162.000 ;
    END
  END mprj_adr_o_user[23]
  PIN mprj_adr_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 156.000 385.390 162.000 ;
    END
  END mprj_adr_o_user[24]
  PIN mprj_adr_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 156.000 397.810 162.000 ;
    END
  END mprj_adr_o_user[25]
  PIN mprj_adr_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 156.000 410.230 162.000 ;
    END
  END mprj_adr_o_user[26]
  PIN mprj_adr_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 156.000 422.650 162.000 ;
    END
  END mprj_adr_o_user[27]
  PIN mprj_adr_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 156.000 435.070 162.000 ;
    END
  END mprj_adr_o_user[28]
  PIN mprj_adr_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 156.000 447.490 162.000 ;
    END
  END mprj_adr_o_user[29]
  PIN mprj_adr_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 156.000 103.870 162.000 ;
    END
  END mprj_adr_o_user[2]
  PIN mprj_adr_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 156.000 459.910 162.000 ;
    END
  END mprj_adr_o_user[30]
  PIN mprj_adr_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 156.000 472.330 162.000 ;
    END
  END mprj_adr_o_user[31]
  PIN mprj_adr_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 156.000 120.430 162.000 ;
    END
  END mprj_adr_o_user[3]
  PIN mprj_adr_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 156.000 136.990 162.000 ;
    END
  END mprj_adr_o_user[4]
  PIN mprj_adr_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 156.000 149.410 162.000 ;
    END
  END mprj_adr_o_user[5]
  PIN mprj_adr_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 156.000 161.830 162.000 ;
    END
  END mprj_adr_o_user[6]
  PIN mprj_adr_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 156.000 174.250 162.000 ;
    END
  END mprj_adr_o_user[7]
  PIN mprj_adr_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 156.000 186.670 162.000 ;
    END
  END mprj_adr_o_user[8]
  PIN mprj_adr_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 156.000 199.090 162.000 ;
    END
  END mprj_adr_o_user[9]
  PIN mprj_cyc_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.250 -2.000 1723.530 4.000 ;
    END
  END mprj_cyc_o_core
  PIN mprj_cyc_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 156.000 58.330 162.000 ;
    END
  END mprj_cyc_o_user
  PIN mprj_dat_i_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 -2.000 1736.410 4.000 ;
    END
  END mprj_dat_i_core[0]
  PIN mprj_dat_i_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.610 -2.000 1845.890 4.000 ;
    END
  END mprj_dat_i_core[10]
  PIN mprj_dat_i_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.270 -2.000 1855.550 4.000 ;
    END
  END mprj_dat_i_core[11]
  PIN mprj_dat_i_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.930 -2.000 1865.210 4.000 ;
    END
  END mprj_dat_i_core[12]
  PIN mprj_dat_i_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.590 -2.000 1874.870 4.000 ;
    END
  END mprj_dat_i_core[13]
  PIN mprj_dat_i_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1884.250 -2.000 1884.530 4.000 ;
    END
  END mprj_dat_i_core[14]
  PIN mprj_dat_i_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.910 -2.000 1894.190 4.000 ;
    END
  END mprj_dat_i_core[15]
  PIN mprj_dat_i_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.570 -2.000 1903.850 4.000 ;
    END
  END mprj_dat_i_core[16]
  PIN mprj_dat_i_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.230 -2.000 1913.510 4.000 ;
    END
  END mprj_dat_i_core[17]
  PIN mprj_dat_i_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.890 -2.000 1923.170 4.000 ;
    END
  END mprj_dat_i_core[18]
  PIN mprj_dat_i_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.550 -2.000 1932.830 4.000 ;
    END
  END mprj_dat_i_core[19]
  PIN mprj_dat_i_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.010 -2.000 1749.290 4.000 ;
    END
  END mprj_dat_i_core[1]
  PIN mprj_dat_i_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.210 -2.000 1942.490 4.000 ;
    END
  END mprj_dat_i_core[20]
  PIN mprj_dat_i_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.870 -2.000 1952.150 4.000 ;
    END
  END mprj_dat_i_core[21]
  PIN mprj_dat_i_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.530 -2.000 1961.810 4.000 ;
    END
  END mprj_dat_i_core[22]
  PIN mprj_dat_i_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.190 -2.000 1971.470 4.000 ;
    END
  END mprj_dat_i_core[23]
  PIN mprj_dat_i_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.850 -2.000 1981.130 4.000 ;
    END
  END mprj_dat_i_core[24]
  PIN mprj_dat_i_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.510 -2.000 1990.790 4.000 ;
    END
  END mprj_dat_i_core[25]
  PIN mprj_dat_i_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.170 -2.000 2000.450 4.000 ;
    END
  END mprj_dat_i_core[26]
  PIN mprj_dat_i_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.830 -2.000 2010.110 4.000 ;
    END
  END mprj_dat_i_core[27]
  PIN mprj_dat_i_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.490 -2.000 2019.770 4.000 ;
    END
  END mprj_dat_i_core[28]
  PIN mprj_dat_i_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.150 -2.000 2029.430 4.000 ;
    END
  END mprj_dat_i_core[29]
  PIN mprj_dat_i_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.890 -2.000 1762.170 4.000 ;
    END
  END mprj_dat_i_core[2]
  PIN mprj_dat_i_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.810 -2.000 2039.090 4.000 ;
    END
  END mprj_dat_i_core[30]
  PIN mprj_dat_i_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.470 -2.000 2048.750 4.000 ;
    END
  END mprj_dat_i_core[31]
  PIN mprj_dat_i_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.770 -2.000 1775.050 4.000 ;
    END
  END mprj_dat_i_core[3]
  PIN mprj_dat_i_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.650 -2.000 1787.930 4.000 ;
    END
  END mprj_dat_i_core[4]
  PIN mprj_dat_i_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1797.310 -2.000 1797.590 4.000 ;
    END
  END mprj_dat_i_core[5]
  PIN mprj_dat_i_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.970 -2.000 1807.250 4.000 ;
    END
  END mprj_dat_i_core[6]
  PIN mprj_dat_i_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.630 -2.000 1816.910 4.000 ;
    END
  END mprj_dat_i_core[7]
  PIN mprj_dat_i_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.290 -2.000 1826.570 4.000 ;
    END
  END mprj_dat_i_core[8]
  PIN mprj_dat_i_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.950 -2.000 1836.230 4.000 ;
    END
  END mprj_dat_i_core[9]
  PIN mprj_dat_i_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 156.000 74.890 162.000 ;
    END
  END mprj_dat_i_user[0]
  PIN mprj_dat_i_user[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 156.000 215.650 162.000 ;
    END
  END mprj_dat_i_user[10]
  PIN mprj_dat_i_user[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 156.000 228.070 162.000 ;
    END
  END mprj_dat_i_user[11]
  PIN mprj_dat_i_user[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 156.000 240.490 162.000 ;
    END
  END mprj_dat_i_user[12]
  PIN mprj_dat_i_user[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 156.000 252.910 162.000 ;
    END
  END mprj_dat_i_user[13]
  PIN mprj_dat_i_user[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 156.000 265.330 162.000 ;
    END
  END mprj_dat_i_user[14]
  PIN mprj_dat_i_user[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 156.000 277.750 162.000 ;
    END
  END mprj_dat_i_user[15]
  PIN mprj_dat_i_user[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 156.000 290.170 162.000 ;
    END
  END mprj_dat_i_user[16]
  PIN mprj_dat_i_user[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 156.000 302.590 162.000 ;
    END
  END mprj_dat_i_user[17]
  PIN mprj_dat_i_user[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 156.000 315.010 162.000 ;
    END
  END mprj_dat_i_user[18]
  PIN mprj_dat_i_user[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 156.000 327.430 162.000 ;
    END
  END mprj_dat_i_user[19]
  PIN mprj_dat_i_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 156.000 91.450 162.000 ;
    END
  END mprj_dat_i_user[1]
  PIN mprj_dat_i_user[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 156.000 339.850 162.000 ;
    END
  END mprj_dat_i_user[20]
  PIN mprj_dat_i_user[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 156.000 352.270 162.000 ;
    END
  END mprj_dat_i_user[21]
  PIN mprj_dat_i_user[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 156.000 364.690 162.000 ;
    END
  END mprj_dat_i_user[22]
  PIN mprj_dat_i_user[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 156.000 377.110 162.000 ;
    END
  END mprj_dat_i_user[23]
  PIN mprj_dat_i_user[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 156.000 389.530 162.000 ;
    END
  END mprj_dat_i_user[24]
  PIN mprj_dat_i_user[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 156.000 401.950 162.000 ;
    END
  END mprj_dat_i_user[25]
  PIN mprj_dat_i_user[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 156.000 414.370 162.000 ;
    END
  END mprj_dat_i_user[26]
  PIN mprj_dat_i_user[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 156.000 426.790 162.000 ;
    END
  END mprj_dat_i_user[27]
  PIN mprj_dat_i_user[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 156.000 439.210 162.000 ;
    END
  END mprj_dat_i_user[28]
  PIN mprj_dat_i_user[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 156.000 451.630 162.000 ;
    END
  END mprj_dat_i_user[29]
  PIN mprj_dat_i_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 156.000 108.010 162.000 ;
    END
  END mprj_dat_i_user[2]
  PIN mprj_dat_i_user[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 156.000 464.050 162.000 ;
    END
  END mprj_dat_i_user[30]
  PIN mprj_dat_i_user[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 156.000 476.470 162.000 ;
    END
  END mprj_dat_i_user[31]
  PIN mprj_dat_i_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 156.000 124.570 162.000 ;
    END
  END mprj_dat_i_user[3]
  PIN mprj_dat_i_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 156.000 141.130 162.000 ;
    END
  END mprj_dat_i_user[4]
  PIN mprj_dat_i_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 156.000 153.550 162.000 ;
    END
  END mprj_dat_i_user[5]
  PIN mprj_dat_i_user[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 156.000 165.970 162.000 ;
    END
  END mprj_dat_i_user[6]
  PIN mprj_dat_i_user[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 156.000 178.390 162.000 ;
    END
  END mprj_dat_i_user[7]
  PIN mprj_dat_i_user[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 156.000 190.810 162.000 ;
    END
  END mprj_dat_i_user[8]
  PIN mprj_dat_i_user[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 156.000 203.230 162.000 ;
    END
  END mprj_dat_i_user[9]
  PIN mprj_dat_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.350 -2.000 1739.630 4.000 ;
    END
  END mprj_dat_o_core[0]
  PIN mprj_dat_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.830 -2.000 1849.110 4.000 ;
    END
  END mprj_dat_o_core[10]
  PIN mprj_dat_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.490 -2.000 1858.770 4.000 ;
    END
  END mprj_dat_o_core[11]
  PIN mprj_dat_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 -2.000 1868.430 4.000 ;
    END
  END mprj_dat_o_core[12]
  PIN mprj_dat_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.810 -2.000 1878.090 4.000 ;
    END
  END mprj_dat_o_core[13]
  PIN mprj_dat_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 -2.000 1887.750 4.000 ;
    END
  END mprj_dat_o_core[14]
  PIN mprj_dat_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.130 -2.000 1897.410 4.000 ;
    END
  END mprj_dat_o_core[15]
  PIN mprj_dat_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.790 -2.000 1907.070 4.000 ;
    END
  END mprj_dat_o_core[16]
  PIN mprj_dat_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.450 -2.000 1916.730 4.000 ;
    END
  END mprj_dat_o_core[17]
  PIN mprj_dat_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.110 -2.000 1926.390 4.000 ;
    END
  END mprj_dat_o_core[18]
  PIN mprj_dat_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.770 -2.000 1936.050 4.000 ;
    END
  END mprj_dat_o_core[19]
  PIN mprj_dat_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.230 -2.000 1752.510 4.000 ;
    END
  END mprj_dat_o_core[1]
  PIN mprj_dat_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.430 -2.000 1945.710 4.000 ;
    END
  END mprj_dat_o_core[20]
  PIN mprj_dat_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.090 -2.000 1955.370 4.000 ;
    END
  END mprj_dat_o_core[21]
  PIN mprj_dat_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.750 -2.000 1965.030 4.000 ;
    END
  END mprj_dat_o_core[22]
  PIN mprj_dat_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.410 -2.000 1974.690 4.000 ;
    END
  END mprj_dat_o_core[23]
  PIN mprj_dat_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.070 -2.000 1984.350 4.000 ;
    END
  END mprj_dat_o_core[24]
  PIN mprj_dat_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.730 -2.000 1994.010 4.000 ;
    END
  END mprj_dat_o_core[25]
  PIN mprj_dat_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.390 -2.000 2003.670 4.000 ;
    END
  END mprj_dat_o_core[26]
  PIN mprj_dat_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.050 -2.000 2013.330 4.000 ;
    END
  END mprj_dat_o_core[27]
  PIN mprj_dat_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.710 -2.000 2022.990 4.000 ;
    END
  END mprj_dat_o_core[28]
  PIN mprj_dat_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2032.370 -2.000 2032.650 4.000 ;
    END
  END mprj_dat_o_core[29]
  PIN mprj_dat_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.110 -2.000 1765.390 4.000 ;
    END
  END mprj_dat_o_core[2]
  PIN mprj_dat_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.030 -2.000 2042.310 4.000 ;
    END
  END mprj_dat_o_core[30]
  PIN mprj_dat_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.690 -2.000 2051.970 4.000 ;
    END
  END mprj_dat_o_core[31]
  PIN mprj_dat_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.990 -2.000 1778.270 4.000 ;
    END
  END mprj_dat_o_core[3]
  PIN mprj_dat_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.870 -2.000 1791.150 4.000 ;
    END
  END mprj_dat_o_core[4]
  PIN mprj_dat_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.530 -2.000 1800.810 4.000 ;
    END
  END mprj_dat_o_core[5]
  PIN mprj_dat_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.190 -2.000 1810.470 4.000 ;
    END
  END mprj_dat_o_core[6]
  PIN mprj_dat_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.850 -2.000 1820.130 4.000 ;
    END
  END mprj_dat_o_core[7]
  PIN mprj_dat_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.510 -2.000 1829.790 4.000 ;
    END
  END mprj_dat_o_core[8]
  PIN mprj_dat_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.170 -2.000 1839.450 4.000 ;
    END
  END mprj_dat_o_core[9]
  PIN mprj_dat_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 156.000 79.030 162.000 ;
    END
  END mprj_dat_o_user[0]
  PIN mprj_dat_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 156.000 219.790 162.000 ;
    END
  END mprj_dat_o_user[10]
  PIN mprj_dat_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 156.000 232.210 162.000 ;
    END
  END mprj_dat_o_user[11]
  PIN mprj_dat_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 156.000 244.630 162.000 ;
    END
  END mprj_dat_o_user[12]
  PIN mprj_dat_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 156.000 257.050 162.000 ;
    END
  END mprj_dat_o_user[13]
  PIN mprj_dat_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 156.000 269.470 162.000 ;
    END
  END mprj_dat_o_user[14]
  PIN mprj_dat_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 156.000 281.890 162.000 ;
    END
  END mprj_dat_o_user[15]
  PIN mprj_dat_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 156.000 294.310 162.000 ;
    END
  END mprj_dat_o_user[16]
  PIN mprj_dat_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 156.000 306.730 162.000 ;
    END
  END mprj_dat_o_user[17]
  PIN mprj_dat_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 156.000 319.150 162.000 ;
    END
  END mprj_dat_o_user[18]
  PIN mprj_dat_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 156.000 331.570 162.000 ;
    END
  END mprj_dat_o_user[19]
  PIN mprj_dat_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 156.000 95.590 162.000 ;
    END
  END mprj_dat_o_user[1]
  PIN mprj_dat_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 156.000 343.990 162.000 ;
    END
  END mprj_dat_o_user[20]
  PIN mprj_dat_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 156.000 356.410 162.000 ;
    END
  END mprj_dat_o_user[21]
  PIN mprj_dat_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 156.000 368.830 162.000 ;
    END
  END mprj_dat_o_user[22]
  PIN mprj_dat_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 156.000 381.250 162.000 ;
    END
  END mprj_dat_o_user[23]
  PIN mprj_dat_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 156.000 393.670 162.000 ;
    END
  END mprj_dat_o_user[24]
  PIN mprj_dat_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 156.000 406.090 162.000 ;
    END
  END mprj_dat_o_user[25]
  PIN mprj_dat_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 156.000 418.510 162.000 ;
    END
  END mprj_dat_o_user[26]
  PIN mprj_dat_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 156.000 430.930 162.000 ;
    END
  END mprj_dat_o_user[27]
  PIN mprj_dat_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 156.000 443.350 162.000 ;
    END
  END mprj_dat_o_user[28]
  PIN mprj_dat_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 156.000 455.770 162.000 ;
    END
  END mprj_dat_o_user[29]
  PIN mprj_dat_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 156.000 112.150 162.000 ;
    END
  END mprj_dat_o_user[2]
  PIN mprj_dat_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 156.000 468.190 162.000 ;
    END
  END mprj_dat_o_user[30]
  PIN mprj_dat_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 156.000 480.610 162.000 ;
    END
  END mprj_dat_o_user[31]
  PIN mprj_dat_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 156.000 128.710 162.000 ;
    END
  END mprj_dat_o_user[3]
  PIN mprj_dat_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 156.000 145.270 162.000 ;
    END
  END mprj_dat_o_user[4]
  PIN mprj_dat_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 156.000 157.690 162.000 ;
    END
  END mprj_dat_o_user[5]
  PIN mprj_dat_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 156.000 170.110 162.000 ;
    END
  END mprj_dat_o_user[6]
  PIN mprj_dat_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 156.000 182.530 162.000 ;
    END
  END mprj_dat_o_user[7]
  PIN mprj_dat_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 156.000 194.950 162.000 ;
    END
  END mprj_dat_o_user[8]
  PIN mprj_dat_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 156.000 207.370 162.000 ;
    END
  END mprj_dat_o_user[9]
  PIN mprj_iena_wb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.910 -2.000 2055.190 4.000 ;
    END
  END mprj_iena_wb
  PIN mprj_sel_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.570 -2.000 1742.850 4.000 ;
    END
  END mprj_sel_o_core[0]
  PIN mprj_sel_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.450 -2.000 1755.730 4.000 ;
    END
  END mprj_sel_o_core[1]
  PIN mprj_sel_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.330 -2.000 1768.610 4.000 ;
    END
  END mprj_sel_o_core[2]
  PIN mprj_sel_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.210 -2.000 1781.490 4.000 ;
    END
  END mprj_sel_o_core[3]
  PIN mprj_sel_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 156.000 83.170 162.000 ;
    END
  END mprj_sel_o_user[0]
  PIN mprj_sel_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 156.000 99.730 162.000 ;
    END
  END mprj_sel_o_user[1]
  PIN mprj_sel_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 156.000 116.290 162.000 ;
    END
  END mprj_sel_o_user[2]
  PIN mprj_sel_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 156.000 132.850 162.000 ;
    END
  END mprj_sel_o_user[3]
  PIN mprj_stb_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.470 -2.000 1726.750 4.000 ;
    END
  END mprj_stb_o_core
  PIN mprj_stb_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 156.000 62.470 162.000 ;
    END
  END mprj_stb_o_user
  PIN mprj_we_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.690 -2.000 1729.970 4.000 ;
    END
  END mprj_we_o_core
  PIN mprj_we_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 156.000 66.610 162.000 ;
    END
  END mprj_we_o_user
  PIN user1_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 52.400 2122.000 53.000 ;
    END
  END user1_vcc_powergood
  PIN user1_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 63.280 2122.000 63.880 ;
    END
  END user1_vdd_powergood
  PIN user2_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 74.160 2122.000 74.760 ;
    END
  END user2_vcc_powergood
  PIN user2_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 85.040 2122.000 85.640 ;
    END
  END user2_vdd_powergood
  PIN user_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 156.000 45.910 162.000 ;
    END
  END user_clock
  PIN user_clock2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2074.230 156.000 2074.510 162.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 95.920 2122.000 96.520 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 106.800 2122.000 107.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 117.680 2122.000 118.280 ;
    END
  END user_irq[2]
  PIN user_irq_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 8.880 2122.000 9.480 ;
    END
  END user_irq_core[0]
  PIN user_irq_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 19.760 2122.000 20.360 ;
    END
  END user_irq_core[1]
  PIN user_irq_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 30.640 2122.000 31.240 ;
    END
  END user_irq_core[2]
  PIN user_irq_ena[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 128.560 2122.000 129.160 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 139.440 2122.000 140.040 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2116.000 150.320 2122.000 150.920 ;
    END
  END user_irq_ena[2]
  PIN user_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 156.000 50.050 162.000 ;
    END
  END user_reset
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.070 5.200 25.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.320 5.200 101.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.570 5.200 176.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.820 5.200 251.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.070 5.200 326.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 401.320 5.200 402.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 476.570 5.200 477.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 551.820 5.200 552.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.070 5.200 627.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 702.320 5.200 703.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 5.200 778.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 852.820 5.200 853.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 928.070 5.200 928.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1003.320 5.200 1004.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1078.570 5.200 1079.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1153.820 5.200 1154.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1229.070 5.200 1229.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.320 5.200 1305.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1379.570 5.200 1380.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.820 5.200 1455.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1530.070 5.200 1530.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1605.320 5.200 1606.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1680.570 5.200 1681.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.820 5.200 1756.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.070 5.200 1831.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1906.320 5.200 1907.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1981.570 5.200 1982.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.820 5.200 2057.720 152.560 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 706.420 5.200 707.320 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 781.670 5.200 782.570 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.920 5.200 857.820 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.170 5.200 933.070 152.560 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.270 5.200 335.170 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.270 5.200 385.170 152.560 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1279.070 5.200 1279.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1354.320 5.200 1355.220 152.560 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1283.070 5.200 1283.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.320 5.200 1359.220 152.560 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1315.970 5.200 1316.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1391.220 5.200 1392.120 152.560 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1319.970 5.200 1320.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.220 5.200 1396.120 152.560 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 61.970 5.200 62.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 137.220 5.200 138.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.470 5.200 213.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 287.720 5.200 288.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 362.970 5.200 363.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 438.220 5.200 439.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.470 5.200 514.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 588.720 5.200 589.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 663.970 5.200 664.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 739.220 5.200 740.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.470 5.200 815.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 889.720 5.200 890.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.970 5.200 965.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1040.220 5.200 1041.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.470 5.200 1116.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1190.720 5.200 1191.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1265.970 5.200 1266.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1341.220 5.200 1342.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1416.470 5.200 1417.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.720 5.200 1492.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1566.970 5.200 1567.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1642.220 5.200 1643.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1717.470 5.200 1718.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1792.720 5.200 1793.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1867.970 5.200 1868.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.220 5.200 1944.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2018.470 5.200 2019.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2093.720 5.200 2094.620 152.560 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 743.320 5.200 744.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.570 5.200 819.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 893.820 5.200 894.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 969.070 5.200 969.970 152.560 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 355.170 5.200 356.070 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.170 5.200 406.070 152.560 ;
    END
  END vssd2
  OBS
      LAYER nwell ;
        RECT 5.330 148.185 2114.350 151.015 ;
        RECT 5.330 142.745 2114.350 145.575 ;
        RECT 5.330 137.305 2114.350 140.135 ;
        RECT 5.330 131.865 2114.350 134.695 ;
        RECT 5.330 126.425 2114.350 129.255 ;
        RECT 5.330 120.985 2114.350 123.815 ;
        RECT 5.330 115.545 2114.350 118.375 ;
        RECT 5.330 110.105 2114.350 112.935 ;
        RECT 5.330 104.665 2114.350 107.495 ;
        RECT 5.330 99.225 2114.350 102.055 ;
        RECT 5.330 93.785 2114.350 96.615 ;
        RECT 5.330 88.345 2114.350 91.175 ;
        RECT 5.330 82.905 2114.350 85.735 ;
        RECT 5.330 77.465 668.570 80.295 ;
        RECT 5.330 72.025 668.570 74.855 ;
        RECT 5.330 66.585 668.570 69.415 ;
        RECT 5.330 61.145 668.570 63.975 ;
        RECT 5.330 56.930 668.570 58.535 ;
        RECT 5.330 55.705 320.350 56.930 ;
        RECT 5.330 50.265 320.350 53.095 ;
        RECT 5.330 44.825 320.350 47.655 ;
        RECT 5.330 39.385 320.350 42.215 ;
        RECT 5.330 33.945 320.350 36.775 ;
        RECT 5.330 28.505 320.350 31.335 ;
        RECT 5.330 23.065 2114.350 25.895 ;
        RECT 5.330 17.625 2114.350 20.455 ;
        RECT 5.330 12.185 2114.350 15.015 ;
        RECT 5.330 6.745 2114.350 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 2114.160 152.405 ;
      LAYER met1 ;
        RECT 5.520 0.040 2114.160 155.680 ;
      LAYER met2 ;
        RECT 25.180 155.720 45.350 156.810 ;
        RECT 46.190 155.720 49.490 156.810 ;
        RECT 50.330 155.720 53.630 156.810 ;
        RECT 54.470 155.720 57.770 156.810 ;
        RECT 58.610 155.720 61.910 156.810 ;
        RECT 62.750 155.720 66.050 156.810 ;
        RECT 66.890 155.720 70.190 156.810 ;
        RECT 71.030 155.720 74.330 156.810 ;
        RECT 75.170 155.720 78.470 156.810 ;
        RECT 79.310 155.720 82.610 156.810 ;
        RECT 83.450 155.720 86.750 156.810 ;
        RECT 87.590 155.720 90.890 156.810 ;
        RECT 91.730 155.720 95.030 156.810 ;
        RECT 95.870 155.720 99.170 156.810 ;
        RECT 100.010 155.720 103.310 156.810 ;
        RECT 104.150 155.720 107.450 156.810 ;
        RECT 108.290 155.720 111.590 156.810 ;
        RECT 112.430 155.720 115.730 156.810 ;
        RECT 116.570 155.720 119.870 156.810 ;
        RECT 120.710 155.720 124.010 156.810 ;
        RECT 124.850 155.720 128.150 156.810 ;
        RECT 128.990 155.720 132.290 156.810 ;
        RECT 133.130 155.720 136.430 156.810 ;
        RECT 137.270 155.720 140.570 156.810 ;
        RECT 141.410 155.720 144.710 156.810 ;
        RECT 145.550 155.720 148.850 156.810 ;
        RECT 149.690 155.720 152.990 156.810 ;
        RECT 153.830 155.720 157.130 156.810 ;
        RECT 157.970 155.720 161.270 156.810 ;
        RECT 162.110 155.720 165.410 156.810 ;
        RECT 166.250 155.720 169.550 156.810 ;
        RECT 170.390 155.720 173.690 156.810 ;
        RECT 174.530 155.720 177.830 156.810 ;
        RECT 178.670 155.720 181.970 156.810 ;
        RECT 182.810 155.720 186.110 156.810 ;
        RECT 186.950 155.720 190.250 156.810 ;
        RECT 191.090 155.720 194.390 156.810 ;
        RECT 195.230 155.720 198.530 156.810 ;
        RECT 199.370 155.720 202.670 156.810 ;
        RECT 203.510 155.720 206.810 156.810 ;
        RECT 207.650 155.720 210.950 156.810 ;
        RECT 211.790 155.720 215.090 156.810 ;
        RECT 215.930 155.720 219.230 156.810 ;
        RECT 220.070 155.720 223.370 156.810 ;
        RECT 224.210 155.720 227.510 156.810 ;
        RECT 228.350 155.720 231.650 156.810 ;
        RECT 232.490 155.720 235.790 156.810 ;
        RECT 236.630 155.720 239.930 156.810 ;
        RECT 240.770 155.720 244.070 156.810 ;
        RECT 244.910 155.720 248.210 156.810 ;
        RECT 249.050 155.720 252.350 156.810 ;
        RECT 253.190 155.720 256.490 156.810 ;
        RECT 257.330 155.720 260.630 156.810 ;
        RECT 261.470 155.720 264.770 156.810 ;
        RECT 265.610 155.720 268.910 156.810 ;
        RECT 269.750 155.720 273.050 156.810 ;
        RECT 273.890 155.720 277.190 156.810 ;
        RECT 278.030 155.720 281.330 156.810 ;
        RECT 282.170 155.720 285.470 156.810 ;
        RECT 286.310 155.720 289.610 156.810 ;
        RECT 290.450 155.720 293.750 156.810 ;
        RECT 294.590 155.720 297.890 156.810 ;
        RECT 298.730 155.720 302.030 156.810 ;
        RECT 302.870 155.720 306.170 156.810 ;
        RECT 307.010 155.720 310.310 156.810 ;
        RECT 311.150 155.720 314.450 156.810 ;
        RECT 315.290 155.720 318.590 156.810 ;
        RECT 319.430 155.720 322.730 156.810 ;
        RECT 323.570 155.720 326.870 156.810 ;
        RECT 327.710 155.720 331.010 156.810 ;
        RECT 331.850 155.720 335.150 156.810 ;
        RECT 335.990 155.720 339.290 156.810 ;
        RECT 340.130 155.720 343.430 156.810 ;
        RECT 344.270 155.720 347.570 156.810 ;
        RECT 348.410 155.720 351.710 156.810 ;
        RECT 352.550 155.720 355.850 156.810 ;
        RECT 356.690 155.720 359.990 156.810 ;
        RECT 360.830 155.720 364.130 156.810 ;
        RECT 364.970 155.720 368.270 156.810 ;
        RECT 369.110 155.720 372.410 156.810 ;
        RECT 373.250 155.720 376.550 156.810 ;
        RECT 377.390 155.720 380.690 156.810 ;
        RECT 381.530 155.720 384.830 156.810 ;
        RECT 385.670 155.720 388.970 156.810 ;
        RECT 389.810 155.720 393.110 156.810 ;
        RECT 393.950 155.720 397.250 156.810 ;
        RECT 398.090 155.720 401.390 156.810 ;
        RECT 402.230 155.720 405.530 156.810 ;
        RECT 406.370 155.720 409.670 156.810 ;
        RECT 410.510 155.720 413.810 156.810 ;
        RECT 414.650 155.720 417.950 156.810 ;
        RECT 418.790 155.720 422.090 156.810 ;
        RECT 422.930 155.720 426.230 156.810 ;
        RECT 427.070 155.720 430.370 156.810 ;
        RECT 431.210 155.720 434.510 156.810 ;
        RECT 435.350 155.720 438.650 156.810 ;
        RECT 439.490 155.720 442.790 156.810 ;
        RECT 443.630 155.720 446.930 156.810 ;
        RECT 447.770 155.720 451.070 156.810 ;
        RECT 451.910 155.720 455.210 156.810 ;
        RECT 456.050 155.720 459.350 156.810 ;
        RECT 460.190 155.720 463.490 156.810 ;
        RECT 464.330 155.720 467.630 156.810 ;
        RECT 468.470 155.720 471.770 156.810 ;
        RECT 472.610 155.720 475.910 156.810 ;
        RECT 476.750 155.720 480.050 156.810 ;
        RECT 480.890 155.720 484.190 156.810 ;
        RECT 485.030 155.720 488.330 156.810 ;
        RECT 489.170 155.720 492.470 156.810 ;
        RECT 493.310 155.720 496.610 156.810 ;
        RECT 497.450 155.720 500.750 156.810 ;
        RECT 501.590 155.720 504.890 156.810 ;
        RECT 505.730 155.720 509.030 156.810 ;
        RECT 509.870 155.720 513.170 156.810 ;
        RECT 514.010 155.720 517.310 156.810 ;
        RECT 518.150 155.720 521.450 156.810 ;
        RECT 522.290 155.720 525.590 156.810 ;
        RECT 526.430 155.720 529.730 156.810 ;
        RECT 530.570 155.720 533.870 156.810 ;
        RECT 534.710 155.720 538.010 156.810 ;
        RECT 538.850 155.720 542.150 156.810 ;
        RECT 542.990 155.720 546.290 156.810 ;
        RECT 547.130 155.720 550.430 156.810 ;
        RECT 551.270 155.720 554.570 156.810 ;
        RECT 555.410 155.720 558.710 156.810 ;
        RECT 559.550 155.720 562.850 156.810 ;
        RECT 563.690 155.720 566.990 156.810 ;
        RECT 567.830 155.720 571.130 156.810 ;
        RECT 571.970 155.720 575.270 156.810 ;
        RECT 576.110 155.720 579.410 156.810 ;
        RECT 580.250 155.720 583.550 156.810 ;
        RECT 584.390 155.720 587.690 156.810 ;
        RECT 588.530 155.720 591.830 156.810 ;
        RECT 592.670 155.720 595.970 156.810 ;
        RECT 596.810 155.720 600.110 156.810 ;
        RECT 600.950 155.720 604.250 156.810 ;
        RECT 605.090 155.720 608.390 156.810 ;
        RECT 609.230 155.720 612.530 156.810 ;
        RECT 613.370 155.720 616.670 156.810 ;
        RECT 617.510 155.720 620.810 156.810 ;
        RECT 621.650 155.720 624.950 156.810 ;
        RECT 625.790 155.720 629.090 156.810 ;
        RECT 629.930 155.720 633.230 156.810 ;
        RECT 634.070 155.720 637.370 156.810 ;
        RECT 638.210 155.720 641.510 156.810 ;
        RECT 642.350 155.720 645.650 156.810 ;
        RECT 646.490 155.720 649.790 156.810 ;
        RECT 650.630 155.720 653.930 156.810 ;
        RECT 654.770 155.720 658.070 156.810 ;
        RECT 658.910 155.720 662.210 156.810 ;
        RECT 663.050 155.720 666.350 156.810 ;
        RECT 667.190 155.720 670.490 156.810 ;
        RECT 671.330 155.720 674.630 156.810 ;
        RECT 675.470 155.720 678.770 156.810 ;
        RECT 679.610 155.720 682.910 156.810 ;
        RECT 683.750 155.720 687.050 156.810 ;
        RECT 687.890 155.720 691.190 156.810 ;
        RECT 692.030 155.720 695.330 156.810 ;
        RECT 696.170 155.720 699.470 156.810 ;
        RECT 700.310 155.720 703.610 156.810 ;
        RECT 704.450 155.720 707.750 156.810 ;
        RECT 708.590 155.720 711.890 156.810 ;
        RECT 712.730 155.720 716.030 156.810 ;
        RECT 716.870 155.720 720.170 156.810 ;
        RECT 721.010 155.720 724.310 156.810 ;
        RECT 725.150 155.720 728.450 156.810 ;
        RECT 729.290 155.720 732.590 156.810 ;
        RECT 733.430 155.720 736.730 156.810 ;
        RECT 737.570 155.720 740.870 156.810 ;
        RECT 741.710 155.720 745.010 156.810 ;
        RECT 745.850 155.720 749.150 156.810 ;
        RECT 749.990 155.720 753.290 156.810 ;
        RECT 754.130 155.720 757.430 156.810 ;
        RECT 758.270 155.720 761.570 156.810 ;
        RECT 762.410 155.720 765.710 156.810 ;
        RECT 766.550 155.720 769.850 156.810 ;
        RECT 770.690 155.720 773.990 156.810 ;
        RECT 774.830 155.720 778.130 156.810 ;
        RECT 778.970 155.720 782.270 156.810 ;
        RECT 783.110 155.720 786.410 156.810 ;
        RECT 787.250 155.720 790.550 156.810 ;
        RECT 791.390 155.720 794.690 156.810 ;
        RECT 795.530 155.720 798.830 156.810 ;
        RECT 799.670 155.720 802.970 156.810 ;
        RECT 803.810 155.720 807.110 156.810 ;
        RECT 807.950 155.720 811.250 156.810 ;
        RECT 812.090 155.720 815.390 156.810 ;
        RECT 816.230 155.720 819.530 156.810 ;
        RECT 820.370 155.720 823.670 156.810 ;
        RECT 824.510 155.720 827.810 156.810 ;
        RECT 828.650 155.720 831.950 156.810 ;
        RECT 832.790 155.720 836.090 156.810 ;
        RECT 836.930 155.720 840.230 156.810 ;
        RECT 841.070 155.720 844.370 156.810 ;
        RECT 845.210 155.720 848.510 156.810 ;
        RECT 849.350 155.720 852.650 156.810 ;
        RECT 853.490 155.720 856.790 156.810 ;
        RECT 857.630 155.720 860.930 156.810 ;
        RECT 861.770 155.720 865.070 156.810 ;
        RECT 865.910 155.720 869.210 156.810 ;
        RECT 870.050 155.720 873.350 156.810 ;
        RECT 874.190 155.720 877.490 156.810 ;
        RECT 878.330 155.720 881.630 156.810 ;
        RECT 882.470 155.720 885.770 156.810 ;
        RECT 886.610 155.720 889.910 156.810 ;
        RECT 890.750 155.720 894.050 156.810 ;
        RECT 894.890 155.720 898.190 156.810 ;
        RECT 899.030 155.720 902.330 156.810 ;
        RECT 903.170 155.720 906.470 156.810 ;
        RECT 907.310 155.720 910.610 156.810 ;
        RECT 911.450 155.720 914.750 156.810 ;
        RECT 915.590 155.720 918.890 156.810 ;
        RECT 919.730 155.720 923.030 156.810 ;
        RECT 923.870 155.720 927.170 156.810 ;
        RECT 928.010 155.720 931.310 156.810 ;
        RECT 932.150 155.720 935.450 156.810 ;
        RECT 936.290 155.720 939.590 156.810 ;
        RECT 940.430 155.720 943.730 156.810 ;
        RECT 944.570 155.720 947.870 156.810 ;
        RECT 948.710 155.720 952.010 156.810 ;
        RECT 952.850 155.720 956.150 156.810 ;
        RECT 956.990 155.720 960.290 156.810 ;
        RECT 961.130 155.720 964.430 156.810 ;
        RECT 965.270 155.720 968.570 156.810 ;
        RECT 969.410 155.720 972.710 156.810 ;
        RECT 973.550 155.720 976.850 156.810 ;
        RECT 977.690 155.720 980.990 156.810 ;
        RECT 981.830 155.720 985.130 156.810 ;
        RECT 985.970 155.720 989.270 156.810 ;
        RECT 990.110 155.720 993.410 156.810 ;
        RECT 994.250 155.720 997.550 156.810 ;
        RECT 998.390 155.720 1001.690 156.810 ;
        RECT 1002.530 155.720 1005.830 156.810 ;
        RECT 1006.670 155.720 1009.970 156.810 ;
        RECT 1010.810 155.720 1014.110 156.810 ;
        RECT 1014.950 155.720 1018.250 156.810 ;
        RECT 1019.090 155.720 1022.390 156.810 ;
        RECT 1023.230 155.720 1026.530 156.810 ;
        RECT 1027.370 155.720 1030.670 156.810 ;
        RECT 1031.510 155.720 1034.810 156.810 ;
        RECT 1035.650 155.720 1038.950 156.810 ;
        RECT 1039.790 155.720 1043.090 156.810 ;
        RECT 1043.930 155.720 1047.230 156.810 ;
        RECT 1048.070 155.720 1051.370 156.810 ;
        RECT 1052.210 155.720 1055.510 156.810 ;
        RECT 1056.350 155.720 1059.650 156.810 ;
        RECT 1060.490 155.720 1063.790 156.810 ;
        RECT 1064.630 155.720 1067.930 156.810 ;
        RECT 1068.770 155.720 1072.070 156.810 ;
        RECT 1072.910 155.720 1076.210 156.810 ;
        RECT 1077.050 155.720 1080.350 156.810 ;
        RECT 1081.190 155.720 1084.490 156.810 ;
        RECT 1085.330 155.720 1088.630 156.810 ;
        RECT 1089.470 155.720 1092.770 156.810 ;
        RECT 1093.610 155.720 1096.910 156.810 ;
        RECT 1097.750 155.720 1101.050 156.810 ;
        RECT 1101.890 155.720 1105.190 156.810 ;
        RECT 1106.030 155.720 1109.330 156.810 ;
        RECT 1110.170 155.720 1113.470 156.810 ;
        RECT 1114.310 155.720 1117.610 156.810 ;
        RECT 1118.450 155.720 1121.750 156.810 ;
        RECT 1122.590 155.720 1125.890 156.810 ;
        RECT 1126.730 155.720 1130.030 156.810 ;
        RECT 1130.870 155.720 1134.170 156.810 ;
        RECT 1135.010 155.720 1138.310 156.810 ;
        RECT 1139.150 155.720 1142.450 156.810 ;
        RECT 1143.290 155.720 1146.590 156.810 ;
        RECT 1147.430 155.720 1150.730 156.810 ;
        RECT 1151.570 155.720 1154.870 156.810 ;
        RECT 1155.710 155.720 1159.010 156.810 ;
        RECT 1159.850 155.720 1163.150 156.810 ;
        RECT 1163.990 155.720 1167.290 156.810 ;
        RECT 1168.130 155.720 1171.430 156.810 ;
        RECT 1172.270 155.720 1175.570 156.810 ;
        RECT 1176.410 155.720 1179.710 156.810 ;
        RECT 1180.550 155.720 1183.850 156.810 ;
        RECT 1184.690 155.720 1187.990 156.810 ;
        RECT 1188.830 155.720 1192.130 156.810 ;
        RECT 1192.970 155.720 1196.270 156.810 ;
        RECT 1197.110 155.720 1200.410 156.810 ;
        RECT 1201.250 155.720 1204.550 156.810 ;
        RECT 1205.390 155.720 1208.690 156.810 ;
        RECT 1209.530 155.720 1212.830 156.810 ;
        RECT 1213.670 155.720 1216.970 156.810 ;
        RECT 1217.810 155.720 1221.110 156.810 ;
        RECT 1221.950 155.720 1225.250 156.810 ;
        RECT 1226.090 155.720 1229.390 156.810 ;
        RECT 1230.230 155.720 1233.530 156.810 ;
        RECT 1234.370 155.720 1237.670 156.810 ;
        RECT 1238.510 155.720 1241.810 156.810 ;
        RECT 1242.650 155.720 1245.950 156.810 ;
        RECT 1246.790 155.720 1250.090 156.810 ;
        RECT 1250.930 155.720 1254.230 156.810 ;
        RECT 1255.070 155.720 1258.370 156.810 ;
        RECT 1259.210 155.720 1262.510 156.810 ;
        RECT 1263.350 155.720 1266.650 156.810 ;
        RECT 1267.490 155.720 1270.790 156.810 ;
        RECT 1271.630 155.720 1274.930 156.810 ;
        RECT 1275.770 155.720 1279.070 156.810 ;
        RECT 1279.910 155.720 1283.210 156.810 ;
        RECT 1284.050 155.720 1287.350 156.810 ;
        RECT 1288.190 155.720 1291.490 156.810 ;
        RECT 1292.330 155.720 1295.630 156.810 ;
        RECT 1296.470 155.720 1299.770 156.810 ;
        RECT 1300.610 155.720 1303.910 156.810 ;
        RECT 1304.750 155.720 1308.050 156.810 ;
        RECT 1308.890 155.720 1312.190 156.810 ;
        RECT 1313.030 155.720 1316.330 156.810 ;
        RECT 1317.170 155.720 1320.470 156.810 ;
        RECT 1321.310 155.720 1324.610 156.810 ;
        RECT 1325.450 155.720 1328.750 156.810 ;
        RECT 1329.590 155.720 1332.890 156.810 ;
        RECT 1333.730 155.720 1337.030 156.810 ;
        RECT 1337.870 155.720 1341.170 156.810 ;
        RECT 1342.010 155.720 1345.310 156.810 ;
        RECT 1346.150 155.720 1349.450 156.810 ;
        RECT 1350.290 155.720 1353.590 156.810 ;
        RECT 1354.430 155.720 1357.730 156.810 ;
        RECT 1358.570 155.720 1361.870 156.810 ;
        RECT 1362.710 155.720 1366.010 156.810 ;
        RECT 1366.850 155.720 1370.150 156.810 ;
        RECT 1370.990 155.720 1374.290 156.810 ;
        RECT 1375.130 155.720 1378.430 156.810 ;
        RECT 1379.270 155.720 1382.570 156.810 ;
        RECT 1383.410 155.720 1386.710 156.810 ;
        RECT 1387.550 155.720 1390.850 156.810 ;
        RECT 1391.690 155.720 1394.990 156.810 ;
        RECT 1395.830 155.720 1399.130 156.810 ;
        RECT 1399.970 155.720 1403.270 156.810 ;
        RECT 1404.110 155.720 1407.410 156.810 ;
        RECT 1408.250 155.720 1411.550 156.810 ;
        RECT 1412.390 155.720 1415.690 156.810 ;
        RECT 1416.530 155.720 1419.830 156.810 ;
        RECT 1420.670 155.720 1423.970 156.810 ;
        RECT 1424.810 155.720 1428.110 156.810 ;
        RECT 1428.950 155.720 1432.250 156.810 ;
        RECT 1433.090 155.720 1436.390 156.810 ;
        RECT 1437.230 155.720 1440.530 156.810 ;
        RECT 1441.370 155.720 1444.670 156.810 ;
        RECT 1445.510 155.720 1448.810 156.810 ;
        RECT 1449.650 155.720 1452.950 156.810 ;
        RECT 1453.790 155.720 1457.090 156.810 ;
        RECT 1457.930 155.720 1461.230 156.810 ;
        RECT 1462.070 155.720 1465.370 156.810 ;
        RECT 1466.210 155.720 1469.510 156.810 ;
        RECT 1470.350 155.720 1473.650 156.810 ;
        RECT 1474.490 155.720 1477.790 156.810 ;
        RECT 1478.630 155.720 1481.930 156.810 ;
        RECT 1482.770 155.720 1486.070 156.810 ;
        RECT 1486.910 155.720 1490.210 156.810 ;
        RECT 1491.050 155.720 1494.350 156.810 ;
        RECT 1495.190 155.720 1498.490 156.810 ;
        RECT 1499.330 155.720 1502.630 156.810 ;
        RECT 1503.470 155.720 1506.770 156.810 ;
        RECT 1507.610 155.720 1510.910 156.810 ;
        RECT 1511.750 155.720 1515.050 156.810 ;
        RECT 1515.890 155.720 1519.190 156.810 ;
        RECT 1520.030 155.720 1523.330 156.810 ;
        RECT 1524.170 155.720 1527.470 156.810 ;
        RECT 1528.310 155.720 1531.610 156.810 ;
        RECT 1532.450 155.720 1535.750 156.810 ;
        RECT 1536.590 155.720 1539.890 156.810 ;
        RECT 1540.730 155.720 1544.030 156.810 ;
        RECT 1544.870 155.720 1548.170 156.810 ;
        RECT 1549.010 155.720 1552.310 156.810 ;
        RECT 1553.150 155.720 1556.450 156.810 ;
        RECT 1557.290 155.720 1560.590 156.810 ;
        RECT 1561.430 155.720 1564.730 156.810 ;
        RECT 1565.570 155.720 1568.870 156.810 ;
        RECT 1569.710 155.720 1573.010 156.810 ;
        RECT 1573.850 155.720 1577.150 156.810 ;
        RECT 1577.990 155.720 1581.290 156.810 ;
        RECT 1582.130 155.720 1585.430 156.810 ;
        RECT 1586.270 155.720 1589.570 156.810 ;
        RECT 1590.410 155.720 1593.710 156.810 ;
        RECT 1594.550 155.720 1597.850 156.810 ;
        RECT 1598.690 155.720 1601.990 156.810 ;
        RECT 1602.830 155.720 1606.130 156.810 ;
        RECT 1606.970 155.720 1610.270 156.810 ;
        RECT 1611.110 155.720 1614.410 156.810 ;
        RECT 1615.250 155.720 1618.550 156.810 ;
        RECT 1619.390 155.720 1622.690 156.810 ;
        RECT 1623.530 155.720 1626.830 156.810 ;
        RECT 1627.670 155.720 1630.970 156.810 ;
        RECT 1631.810 155.720 1635.110 156.810 ;
        RECT 1635.950 155.720 1639.250 156.810 ;
        RECT 1640.090 155.720 1643.390 156.810 ;
        RECT 1644.230 155.720 1647.530 156.810 ;
        RECT 1648.370 155.720 1651.670 156.810 ;
        RECT 1652.510 155.720 1655.810 156.810 ;
        RECT 1656.650 155.720 1659.950 156.810 ;
        RECT 1660.790 155.720 1664.090 156.810 ;
        RECT 1664.930 155.720 1668.230 156.810 ;
        RECT 1669.070 155.720 1672.370 156.810 ;
        RECT 1673.210 155.720 1676.510 156.810 ;
        RECT 1677.350 155.720 1680.650 156.810 ;
        RECT 1681.490 155.720 1684.790 156.810 ;
        RECT 1685.630 155.720 1688.930 156.810 ;
        RECT 1689.770 155.720 1693.070 156.810 ;
        RECT 1693.910 155.720 1697.210 156.810 ;
        RECT 1698.050 155.720 1701.350 156.810 ;
        RECT 1702.190 155.720 1705.490 156.810 ;
        RECT 1706.330 155.720 1709.630 156.810 ;
        RECT 1710.470 155.720 1713.770 156.810 ;
        RECT 1714.610 155.720 1717.910 156.810 ;
        RECT 1718.750 155.720 1722.050 156.810 ;
        RECT 1722.890 155.720 1726.190 156.810 ;
        RECT 1727.030 155.720 1730.330 156.810 ;
        RECT 1731.170 155.720 1734.470 156.810 ;
        RECT 1735.310 155.720 1738.610 156.810 ;
        RECT 1739.450 155.720 1742.750 156.810 ;
        RECT 1743.590 155.720 1746.890 156.810 ;
        RECT 1747.730 155.720 1751.030 156.810 ;
        RECT 1751.870 155.720 1755.170 156.810 ;
        RECT 1756.010 155.720 1759.310 156.810 ;
        RECT 1760.150 155.720 1763.450 156.810 ;
        RECT 1764.290 155.720 1767.590 156.810 ;
        RECT 1768.430 155.720 1771.730 156.810 ;
        RECT 1772.570 155.720 1775.870 156.810 ;
        RECT 1776.710 155.720 1780.010 156.810 ;
        RECT 1780.850 155.720 1784.150 156.810 ;
        RECT 1784.990 155.720 1788.290 156.810 ;
        RECT 1789.130 155.720 1792.430 156.810 ;
        RECT 1793.270 155.720 1796.570 156.810 ;
        RECT 1797.410 155.720 1800.710 156.810 ;
        RECT 1801.550 155.720 1804.850 156.810 ;
        RECT 1805.690 155.720 1808.990 156.810 ;
        RECT 1809.830 155.720 1813.130 156.810 ;
        RECT 1813.970 155.720 1817.270 156.810 ;
        RECT 1818.110 155.720 1821.410 156.810 ;
        RECT 1822.250 155.720 1825.550 156.810 ;
        RECT 1826.390 155.720 1829.690 156.810 ;
        RECT 1830.530 155.720 1833.830 156.810 ;
        RECT 1834.670 155.720 1837.970 156.810 ;
        RECT 1838.810 155.720 1842.110 156.810 ;
        RECT 1842.950 155.720 1846.250 156.810 ;
        RECT 1847.090 155.720 1850.390 156.810 ;
        RECT 1851.230 155.720 1854.530 156.810 ;
        RECT 1855.370 155.720 1858.670 156.810 ;
        RECT 1859.510 155.720 1862.810 156.810 ;
        RECT 1863.650 155.720 1866.950 156.810 ;
        RECT 1867.790 155.720 1871.090 156.810 ;
        RECT 1871.930 155.720 1875.230 156.810 ;
        RECT 1876.070 155.720 1879.370 156.810 ;
        RECT 1880.210 155.720 1883.510 156.810 ;
        RECT 1884.350 155.720 1887.650 156.810 ;
        RECT 1888.490 155.720 1891.790 156.810 ;
        RECT 1892.630 155.720 1895.930 156.810 ;
        RECT 1896.770 155.720 1900.070 156.810 ;
        RECT 1900.910 155.720 1904.210 156.810 ;
        RECT 1905.050 155.720 1908.350 156.810 ;
        RECT 1909.190 155.720 1912.490 156.810 ;
        RECT 1913.330 155.720 1916.630 156.810 ;
        RECT 1917.470 155.720 1920.770 156.810 ;
        RECT 1921.610 155.720 1924.910 156.810 ;
        RECT 1925.750 155.720 1929.050 156.810 ;
        RECT 1929.890 155.720 1933.190 156.810 ;
        RECT 1934.030 155.720 1937.330 156.810 ;
        RECT 1938.170 155.720 1941.470 156.810 ;
        RECT 1942.310 155.720 1945.610 156.810 ;
        RECT 1946.450 155.720 1949.750 156.810 ;
        RECT 1950.590 155.720 1953.890 156.810 ;
        RECT 1954.730 155.720 1958.030 156.810 ;
        RECT 1958.870 155.720 1962.170 156.810 ;
        RECT 1963.010 155.720 1966.310 156.810 ;
        RECT 1967.150 155.720 1970.450 156.810 ;
        RECT 1971.290 155.720 1974.590 156.810 ;
        RECT 1975.430 155.720 1978.730 156.810 ;
        RECT 1979.570 155.720 1982.870 156.810 ;
        RECT 1983.710 155.720 1987.010 156.810 ;
        RECT 1987.850 155.720 1991.150 156.810 ;
        RECT 1991.990 155.720 1995.290 156.810 ;
        RECT 1996.130 155.720 1999.430 156.810 ;
        RECT 2000.270 155.720 2003.570 156.810 ;
        RECT 2004.410 155.720 2007.710 156.810 ;
        RECT 2008.550 155.720 2011.850 156.810 ;
        RECT 2012.690 155.720 2015.990 156.810 ;
        RECT 2016.830 155.720 2020.130 156.810 ;
        RECT 2020.970 155.720 2024.270 156.810 ;
        RECT 2025.110 155.720 2028.410 156.810 ;
        RECT 2029.250 155.720 2032.550 156.810 ;
        RECT 2033.390 155.720 2036.690 156.810 ;
        RECT 2037.530 155.720 2040.830 156.810 ;
        RECT 2041.670 155.720 2044.970 156.810 ;
        RECT 2045.810 155.720 2049.110 156.810 ;
        RECT 2049.950 155.720 2053.250 156.810 ;
        RECT 2054.090 155.720 2057.390 156.810 ;
        RECT 2058.230 155.720 2061.530 156.810 ;
        RECT 2062.370 155.720 2065.670 156.810 ;
        RECT 2066.510 155.720 2069.810 156.810 ;
        RECT 2070.650 155.720 2073.950 156.810 ;
        RECT 2074.790 155.720 2113.150 156.810 ;
        RECT 25.180 4.280 2113.150 155.720 ;
        RECT 25.180 0.010 64.670 4.280 ;
        RECT 65.510 0.010 67.890 4.280 ;
        RECT 68.730 0.010 71.110 4.280 ;
        RECT 71.950 0.010 74.330 4.280 ;
        RECT 75.170 0.010 77.550 4.280 ;
        RECT 78.390 0.010 80.770 4.280 ;
        RECT 81.610 0.010 83.990 4.280 ;
        RECT 84.830 0.010 87.210 4.280 ;
        RECT 88.050 0.010 90.430 4.280 ;
        RECT 91.270 0.010 93.650 4.280 ;
        RECT 94.490 0.010 96.870 4.280 ;
        RECT 97.710 0.010 100.090 4.280 ;
        RECT 100.930 0.010 103.310 4.280 ;
        RECT 104.150 0.010 106.530 4.280 ;
        RECT 107.370 0.010 109.750 4.280 ;
        RECT 110.590 0.010 112.970 4.280 ;
        RECT 113.810 0.010 116.190 4.280 ;
        RECT 117.030 0.010 119.410 4.280 ;
        RECT 120.250 0.010 122.630 4.280 ;
        RECT 123.470 0.010 125.850 4.280 ;
        RECT 126.690 0.010 129.070 4.280 ;
        RECT 129.910 0.010 132.290 4.280 ;
        RECT 133.130 0.010 135.510 4.280 ;
        RECT 136.350 0.010 138.730 4.280 ;
        RECT 139.570 0.010 141.950 4.280 ;
        RECT 142.790 0.010 145.170 4.280 ;
        RECT 146.010 0.010 148.390 4.280 ;
        RECT 149.230 0.010 151.610 4.280 ;
        RECT 152.450 0.010 154.830 4.280 ;
        RECT 155.670 0.010 158.050 4.280 ;
        RECT 158.890 0.010 161.270 4.280 ;
        RECT 162.110 0.010 164.490 4.280 ;
        RECT 165.330 0.010 167.710 4.280 ;
        RECT 168.550 0.010 170.930 4.280 ;
        RECT 171.770 0.010 174.150 4.280 ;
        RECT 174.990 0.010 177.370 4.280 ;
        RECT 178.210 0.010 180.590 4.280 ;
        RECT 181.430 0.010 183.810 4.280 ;
        RECT 184.650 0.010 187.030 4.280 ;
        RECT 187.870 0.010 190.250 4.280 ;
        RECT 191.090 0.010 193.470 4.280 ;
        RECT 194.310 0.010 196.690 4.280 ;
        RECT 197.530 0.010 199.910 4.280 ;
        RECT 200.750 0.010 203.130 4.280 ;
        RECT 203.970 0.010 206.350 4.280 ;
        RECT 207.190 0.010 209.570 4.280 ;
        RECT 210.410 0.010 212.790 4.280 ;
        RECT 213.630 0.010 216.010 4.280 ;
        RECT 216.850 0.010 219.230 4.280 ;
        RECT 220.070 0.010 222.450 4.280 ;
        RECT 223.290 0.010 225.670 4.280 ;
        RECT 226.510 0.010 228.890 4.280 ;
        RECT 229.730 0.010 232.110 4.280 ;
        RECT 232.950 0.010 235.330 4.280 ;
        RECT 236.170 0.010 238.550 4.280 ;
        RECT 239.390 0.010 241.770 4.280 ;
        RECT 242.610 0.010 244.990 4.280 ;
        RECT 245.830 0.010 248.210 4.280 ;
        RECT 249.050 0.010 251.430 4.280 ;
        RECT 252.270 0.010 254.650 4.280 ;
        RECT 255.490 0.010 257.870 4.280 ;
        RECT 258.710 0.010 261.090 4.280 ;
        RECT 261.930 0.010 264.310 4.280 ;
        RECT 265.150 0.010 267.530 4.280 ;
        RECT 268.370 0.010 270.750 4.280 ;
        RECT 271.590 0.010 273.970 4.280 ;
        RECT 274.810 0.010 277.190 4.280 ;
        RECT 278.030 0.010 280.410 4.280 ;
        RECT 281.250 0.010 283.630 4.280 ;
        RECT 284.470 0.010 286.850 4.280 ;
        RECT 287.690 0.010 290.070 4.280 ;
        RECT 290.910 0.010 293.290 4.280 ;
        RECT 294.130 0.010 296.510 4.280 ;
        RECT 297.350 0.010 299.730 4.280 ;
        RECT 300.570 0.010 302.950 4.280 ;
        RECT 303.790 0.010 306.170 4.280 ;
        RECT 307.010 0.010 309.390 4.280 ;
        RECT 310.230 0.010 312.610 4.280 ;
        RECT 313.450 0.010 315.830 4.280 ;
        RECT 316.670 0.010 319.050 4.280 ;
        RECT 319.890 0.010 322.270 4.280 ;
        RECT 323.110 0.010 325.490 4.280 ;
        RECT 326.330 0.010 328.710 4.280 ;
        RECT 329.550 0.010 331.930 4.280 ;
        RECT 332.770 0.010 335.150 4.280 ;
        RECT 335.990 0.010 338.370 4.280 ;
        RECT 339.210 0.010 341.590 4.280 ;
        RECT 342.430 0.010 344.810 4.280 ;
        RECT 345.650 0.010 348.030 4.280 ;
        RECT 348.870 0.010 351.250 4.280 ;
        RECT 352.090 0.010 354.470 4.280 ;
        RECT 355.310 0.010 357.690 4.280 ;
        RECT 358.530 0.010 360.910 4.280 ;
        RECT 361.750 0.010 364.130 4.280 ;
        RECT 364.970 0.010 367.350 4.280 ;
        RECT 368.190 0.010 370.570 4.280 ;
        RECT 371.410 0.010 373.790 4.280 ;
        RECT 374.630 0.010 377.010 4.280 ;
        RECT 377.850 0.010 380.230 4.280 ;
        RECT 381.070 0.010 383.450 4.280 ;
        RECT 384.290 0.010 386.670 4.280 ;
        RECT 387.510 0.010 389.890 4.280 ;
        RECT 390.730 0.010 393.110 4.280 ;
        RECT 393.950 0.010 396.330 4.280 ;
        RECT 397.170 0.010 399.550 4.280 ;
        RECT 400.390 0.010 402.770 4.280 ;
        RECT 403.610 0.010 405.990 4.280 ;
        RECT 406.830 0.010 409.210 4.280 ;
        RECT 410.050 0.010 412.430 4.280 ;
        RECT 413.270 0.010 415.650 4.280 ;
        RECT 416.490 0.010 418.870 4.280 ;
        RECT 419.710 0.010 422.090 4.280 ;
        RECT 422.930 0.010 425.310 4.280 ;
        RECT 426.150 0.010 428.530 4.280 ;
        RECT 429.370 0.010 431.750 4.280 ;
        RECT 432.590 0.010 434.970 4.280 ;
        RECT 435.810 0.010 438.190 4.280 ;
        RECT 439.030 0.010 441.410 4.280 ;
        RECT 442.250 0.010 444.630 4.280 ;
        RECT 445.470 0.010 447.850 4.280 ;
        RECT 448.690 0.010 451.070 4.280 ;
        RECT 451.910 0.010 454.290 4.280 ;
        RECT 455.130 0.010 457.510 4.280 ;
        RECT 458.350 0.010 460.730 4.280 ;
        RECT 461.570 0.010 463.950 4.280 ;
        RECT 464.790 0.010 467.170 4.280 ;
        RECT 468.010 0.010 470.390 4.280 ;
        RECT 471.230 0.010 473.610 4.280 ;
        RECT 474.450 0.010 476.830 4.280 ;
        RECT 477.670 0.010 480.050 4.280 ;
        RECT 480.890 0.010 483.270 4.280 ;
        RECT 484.110 0.010 486.490 4.280 ;
        RECT 487.330 0.010 489.710 4.280 ;
        RECT 490.550 0.010 492.930 4.280 ;
        RECT 493.770 0.010 496.150 4.280 ;
        RECT 496.990 0.010 499.370 4.280 ;
        RECT 500.210 0.010 502.590 4.280 ;
        RECT 503.430 0.010 505.810 4.280 ;
        RECT 506.650 0.010 509.030 4.280 ;
        RECT 509.870 0.010 512.250 4.280 ;
        RECT 513.090 0.010 515.470 4.280 ;
        RECT 516.310 0.010 518.690 4.280 ;
        RECT 519.530 0.010 521.910 4.280 ;
        RECT 522.750 0.010 525.130 4.280 ;
        RECT 525.970 0.010 528.350 4.280 ;
        RECT 529.190 0.010 531.570 4.280 ;
        RECT 532.410 0.010 534.790 4.280 ;
        RECT 535.630 0.010 538.010 4.280 ;
        RECT 538.850 0.010 541.230 4.280 ;
        RECT 542.070 0.010 544.450 4.280 ;
        RECT 545.290 0.010 547.670 4.280 ;
        RECT 548.510 0.010 550.890 4.280 ;
        RECT 551.730 0.010 554.110 4.280 ;
        RECT 554.950 0.010 557.330 4.280 ;
        RECT 558.170 0.010 560.550 4.280 ;
        RECT 561.390 0.010 563.770 4.280 ;
        RECT 564.610 0.010 566.990 4.280 ;
        RECT 567.830 0.010 570.210 4.280 ;
        RECT 571.050 0.010 573.430 4.280 ;
        RECT 574.270 0.010 576.650 4.280 ;
        RECT 577.490 0.010 579.870 4.280 ;
        RECT 580.710 0.010 583.090 4.280 ;
        RECT 583.930 0.010 586.310 4.280 ;
        RECT 587.150 0.010 589.530 4.280 ;
        RECT 590.370 0.010 592.750 4.280 ;
        RECT 593.590 0.010 595.970 4.280 ;
        RECT 596.810 0.010 599.190 4.280 ;
        RECT 600.030 0.010 602.410 4.280 ;
        RECT 603.250 0.010 605.630 4.280 ;
        RECT 606.470 0.010 608.850 4.280 ;
        RECT 609.690 0.010 612.070 4.280 ;
        RECT 612.910 0.010 615.290 4.280 ;
        RECT 616.130 0.010 618.510 4.280 ;
        RECT 619.350 0.010 621.730 4.280 ;
        RECT 622.570 0.010 624.950 4.280 ;
        RECT 625.790 0.010 628.170 4.280 ;
        RECT 629.010 0.010 631.390 4.280 ;
        RECT 632.230 0.010 634.610 4.280 ;
        RECT 635.450 0.010 637.830 4.280 ;
        RECT 638.670 0.010 641.050 4.280 ;
        RECT 641.890 0.010 644.270 4.280 ;
        RECT 645.110 0.010 647.490 4.280 ;
        RECT 648.330 0.010 650.710 4.280 ;
        RECT 651.550 0.010 653.930 4.280 ;
        RECT 654.770 0.010 657.150 4.280 ;
        RECT 657.990 0.010 660.370 4.280 ;
        RECT 661.210 0.010 663.590 4.280 ;
        RECT 664.430 0.010 666.810 4.280 ;
        RECT 667.650 0.010 670.030 4.280 ;
        RECT 670.870 0.010 673.250 4.280 ;
        RECT 674.090 0.010 676.470 4.280 ;
        RECT 677.310 0.010 679.690 4.280 ;
        RECT 680.530 0.010 682.910 4.280 ;
        RECT 683.750 0.010 686.130 4.280 ;
        RECT 686.970 0.010 689.350 4.280 ;
        RECT 690.190 0.010 692.570 4.280 ;
        RECT 693.410 0.010 695.790 4.280 ;
        RECT 696.630 0.010 699.010 4.280 ;
        RECT 699.850 0.010 702.230 4.280 ;
        RECT 703.070 0.010 705.450 4.280 ;
        RECT 706.290 0.010 708.670 4.280 ;
        RECT 709.510 0.010 711.890 4.280 ;
        RECT 712.730 0.010 715.110 4.280 ;
        RECT 715.950 0.010 718.330 4.280 ;
        RECT 719.170 0.010 721.550 4.280 ;
        RECT 722.390 0.010 724.770 4.280 ;
        RECT 725.610 0.010 727.990 4.280 ;
        RECT 728.830 0.010 731.210 4.280 ;
        RECT 732.050 0.010 734.430 4.280 ;
        RECT 735.270 0.010 737.650 4.280 ;
        RECT 738.490 0.010 740.870 4.280 ;
        RECT 741.710 0.010 744.090 4.280 ;
        RECT 744.930 0.010 747.310 4.280 ;
        RECT 748.150 0.010 750.530 4.280 ;
        RECT 751.370 0.010 753.750 4.280 ;
        RECT 754.590 0.010 756.970 4.280 ;
        RECT 757.810 0.010 760.190 4.280 ;
        RECT 761.030 0.010 763.410 4.280 ;
        RECT 764.250 0.010 766.630 4.280 ;
        RECT 767.470 0.010 769.850 4.280 ;
        RECT 770.690 0.010 773.070 4.280 ;
        RECT 773.910 0.010 776.290 4.280 ;
        RECT 777.130 0.010 779.510 4.280 ;
        RECT 780.350 0.010 782.730 4.280 ;
        RECT 783.570 0.010 785.950 4.280 ;
        RECT 786.790 0.010 789.170 4.280 ;
        RECT 790.010 0.010 792.390 4.280 ;
        RECT 793.230 0.010 795.610 4.280 ;
        RECT 796.450 0.010 798.830 4.280 ;
        RECT 799.670 0.010 802.050 4.280 ;
        RECT 802.890 0.010 805.270 4.280 ;
        RECT 806.110 0.010 808.490 4.280 ;
        RECT 809.330 0.010 811.710 4.280 ;
        RECT 812.550 0.010 814.930 4.280 ;
        RECT 815.770 0.010 818.150 4.280 ;
        RECT 818.990 0.010 821.370 4.280 ;
        RECT 822.210 0.010 824.590 4.280 ;
        RECT 825.430 0.010 827.810 4.280 ;
        RECT 828.650 0.010 831.030 4.280 ;
        RECT 831.870 0.010 834.250 4.280 ;
        RECT 835.090 0.010 837.470 4.280 ;
        RECT 838.310 0.010 840.690 4.280 ;
        RECT 841.530 0.010 843.910 4.280 ;
        RECT 844.750 0.010 847.130 4.280 ;
        RECT 847.970 0.010 850.350 4.280 ;
        RECT 851.190 0.010 853.570 4.280 ;
        RECT 854.410 0.010 856.790 4.280 ;
        RECT 857.630 0.010 860.010 4.280 ;
        RECT 860.850 0.010 863.230 4.280 ;
        RECT 864.070 0.010 866.450 4.280 ;
        RECT 867.290 0.010 869.670 4.280 ;
        RECT 870.510 0.010 872.890 4.280 ;
        RECT 873.730 0.010 876.110 4.280 ;
        RECT 876.950 0.010 879.330 4.280 ;
        RECT 880.170 0.010 882.550 4.280 ;
        RECT 883.390 0.010 885.770 4.280 ;
        RECT 886.610 0.010 888.990 4.280 ;
        RECT 889.830 0.010 892.210 4.280 ;
        RECT 893.050 0.010 895.430 4.280 ;
        RECT 896.270 0.010 898.650 4.280 ;
        RECT 899.490 0.010 901.870 4.280 ;
        RECT 902.710 0.010 905.090 4.280 ;
        RECT 905.930 0.010 908.310 4.280 ;
        RECT 909.150 0.010 911.530 4.280 ;
        RECT 912.370 0.010 914.750 4.280 ;
        RECT 915.590 0.010 917.970 4.280 ;
        RECT 918.810 0.010 921.190 4.280 ;
        RECT 922.030 0.010 924.410 4.280 ;
        RECT 925.250 0.010 927.630 4.280 ;
        RECT 928.470 0.010 930.850 4.280 ;
        RECT 931.690 0.010 934.070 4.280 ;
        RECT 934.910 0.010 937.290 4.280 ;
        RECT 938.130 0.010 940.510 4.280 ;
        RECT 941.350 0.010 943.730 4.280 ;
        RECT 944.570 0.010 946.950 4.280 ;
        RECT 947.790 0.010 950.170 4.280 ;
        RECT 951.010 0.010 953.390 4.280 ;
        RECT 954.230 0.010 956.610 4.280 ;
        RECT 957.450 0.010 959.830 4.280 ;
        RECT 960.670 0.010 963.050 4.280 ;
        RECT 963.890 0.010 966.270 4.280 ;
        RECT 967.110 0.010 969.490 4.280 ;
        RECT 970.330 0.010 972.710 4.280 ;
        RECT 973.550 0.010 975.930 4.280 ;
        RECT 976.770 0.010 979.150 4.280 ;
        RECT 979.990 0.010 982.370 4.280 ;
        RECT 983.210 0.010 985.590 4.280 ;
        RECT 986.430 0.010 988.810 4.280 ;
        RECT 989.650 0.010 992.030 4.280 ;
        RECT 992.870 0.010 995.250 4.280 ;
        RECT 996.090 0.010 998.470 4.280 ;
        RECT 999.310 0.010 1001.690 4.280 ;
        RECT 1002.530 0.010 1004.910 4.280 ;
        RECT 1005.750 0.010 1008.130 4.280 ;
        RECT 1008.970 0.010 1011.350 4.280 ;
        RECT 1012.190 0.010 1014.570 4.280 ;
        RECT 1015.410 0.010 1017.790 4.280 ;
        RECT 1018.630 0.010 1021.010 4.280 ;
        RECT 1021.850 0.010 1024.230 4.280 ;
        RECT 1025.070 0.010 1027.450 4.280 ;
        RECT 1028.290 0.010 1030.670 4.280 ;
        RECT 1031.510 0.010 1033.890 4.280 ;
        RECT 1034.730 0.010 1037.110 4.280 ;
        RECT 1037.950 0.010 1040.330 4.280 ;
        RECT 1041.170 0.010 1043.550 4.280 ;
        RECT 1044.390 0.010 1046.770 4.280 ;
        RECT 1047.610 0.010 1049.990 4.280 ;
        RECT 1050.830 0.010 1053.210 4.280 ;
        RECT 1054.050 0.010 1056.430 4.280 ;
        RECT 1057.270 0.010 1059.650 4.280 ;
        RECT 1060.490 0.010 1062.870 4.280 ;
        RECT 1063.710 0.010 1066.090 4.280 ;
        RECT 1066.930 0.010 1069.310 4.280 ;
        RECT 1070.150 0.010 1072.530 4.280 ;
        RECT 1073.370 0.010 1075.750 4.280 ;
        RECT 1076.590 0.010 1078.970 4.280 ;
        RECT 1079.810 0.010 1082.190 4.280 ;
        RECT 1083.030 0.010 1085.410 4.280 ;
        RECT 1086.250 0.010 1088.630 4.280 ;
        RECT 1089.470 0.010 1091.850 4.280 ;
        RECT 1092.690 0.010 1095.070 4.280 ;
        RECT 1095.910 0.010 1098.290 4.280 ;
        RECT 1099.130 0.010 1101.510 4.280 ;
        RECT 1102.350 0.010 1104.730 4.280 ;
        RECT 1105.570 0.010 1107.950 4.280 ;
        RECT 1108.790 0.010 1111.170 4.280 ;
        RECT 1112.010 0.010 1114.390 4.280 ;
        RECT 1115.230 0.010 1117.610 4.280 ;
        RECT 1118.450 0.010 1120.830 4.280 ;
        RECT 1121.670 0.010 1124.050 4.280 ;
        RECT 1124.890 0.010 1127.270 4.280 ;
        RECT 1128.110 0.010 1130.490 4.280 ;
        RECT 1131.330 0.010 1133.710 4.280 ;
        RECT 1134.550 0.010 1136.930 4.280 ;
        RECT 1137.770 0.010 1140.150 4.280 ;
        RECT 1140.990 0.010 1143.370 4.280 ;
        RECT 1144.210 0.010 1146.590 4.280 ;
        RECT 1147.430 0.010 1149.810 4.280 ;
        RECT 1150.650 0.010 1153.030 4.280 ;
        RECT 1153.870 0.010 1156.250 4.280 ;
        RECT 1157.090 0.010 1159.470 4.280 ;
        RECT 1160.310 0.010 1162.690 4.280 ;
        RECT 1163.530 0.010 1165.910 4.280 ;
        RECT 1166.750 0.010 1169.130 4.280 ;
        RECT 1169.970 0.010 1172.350 4.280 ;
        RECT 1173.190 0.010 1175.570 4.280 ;
        RECT 1176.410 0.010 1178.790 4.280 ;
        RECT 1179.630 0.010 1182.010 4.280 ;
        RECT 1182.850 0.010 1185.230 4.280 ;
        RECT 1186.070 0.010 1188.450 4.280 ;
        RECT 1189.290 0.010 1191.670 4.280 ;
        RECT 1192.510 0.010 1194.890 4.280 ;
        RECT 1195.730 0.010 1198.110 4.280 ;
        RECT 1198.950 0.010 1201.330 4.280 ;
        RECT 1202.170 0.010 1204.550 4.280 ;
        RECT 1205.390 0.010 1207.770 4.280 ;
        RECT 1208.610 0.010 1210.990 4.280 ;
        RECT 1211.830 0.010 1214.210 4.280 ;
        RECT 1215.050 0.010 1217.430 4.280 ;
        RECT 1218.270 0.010 1220.650 4.280 ;
        RECT 1221.490 0.010 1223.870 4.280 ;
        RECT 1224.710 0.010 1227.090 4.280 ;
        RECT 1227.930 0.010 1230.310 4.280 ;
        RECT 1231.150 0.010 1233.530 4.280 ;
        RECT 1234.370 0.010 1236.750 4.280 ;
        RECT 1237.590 0.010 1239.970 4.280 ;
        RECT 1240.810 0.010 1243.190 4.280 ;
        RECT 1244.030 0.010 1246.410 4.280 ;
        RECT 1247.250 0.010 1249.630 4.280 ;
        RECT 1250.470 0.010 1252.850 4.280 ;
        RECT 1253.690 0.010 1256.070 4.280 ;
        RECT 1256.910 0.010 1259.290 4.280 ;
        RECT 1260.130 0.010 1262.510 4.280 ;
        RECT 1263.350 0.010 1265.730 4.280 ;
        RECT 1266.570 0.010 1268.950 4.280 ;
        RECT 1269.790 0.010 1272.170 4.280 ;
        RECT 1273.010 0.010 1275.390 4.280 ;
        RECT 1276.230 0.010 1278.610 4.280 ;
        RECT 1279.450 0.010 1281.830 4.280 ;
        RECT 1282.670 0.010 1285.050 4.280 ;
        RECT 1285.890 0.010 1288.270 4.280 ;
        RECT 1289.110 0.010 1291.490 4.280 ;
        RECT 1292.330 0.010 1294.710 4.280 ;
        RECT 1295.550 0.010 1297.930 4.280 ;
        RECT 1298.770 0.010 1301.150 4.280 ;
        RECT 1301.990 0.010 1304.370 4.280 ;
        RECT 1305.210 0.010 1307.590 4.280 ;
        RECT 1308.430 0.010 1310.810 4.280 ;
        RECT 1311.650 0.010 1314.030 4.280 ;
        RECT 1314.870 0.010 1317.250 4.280 ;
        RECT 1318.090 0.010 1320.470 4.280 ;
        RECT 1321.310 0.010 1323.690 4.280 ;
        RECT 1324.530 0.010 1326.910 4.280 ;
        RECT 1327.750 0.010 1330.130 4.280 ;
        RECT 1330.970 0.010 1333.350 4.280 ;
        RECT 1334.190 0.010 1336.570 4.280 ;
        RECT 1337.410 0.010 1339.790 4.280 ;
        RECT 1340.630 0.010 1343.010 4.280 ;
        RECT 1343.850 0.010 1346.230 4.280 ;
        RECT 1347.070 0.010 1349.450 4.280 ;
        RECT 1350.290 0.010 1352.670 4.280 ;
        RECT 1353.510 0.010 1355.890 4.280 ;
        RECT 1356.730 0.010 1359.110 4.280 ;
        RECT 1359.950 0.010 1362.330 4.280 ;
        RECT 1363.170 0.010 1365.550 4.280 ;
        RECT 1366.390 0.010 1368.770 4.280 ;
        RECT 1369.610 0.010 1371.990 4.280 ;
        RECT 1372.830 0.010 1375.210 4.280 ;
        RECT 1376.050 0.010 1378.430 4.280 ;
        RECT 1379.270 0.010 1381.650 4.280 ;
        RECT 1382.490 0.010 1384.870 4.280 ;
        RECT 1385.710 0.010 1388.090 4.280 ;
        RECT 1388.930 0.010 1391.310 4.280 ;
        RECT 1392.150 0.010 1394.530 4.280 ;
        RECT 1395.370 0.010 1397.750 4.280 ;
        RECT 1398.590 0.010 1400.970 4.280 ;
        RECT 1401.810 0.010 1404.190 4.280 ;
        RECT 1405.030 0.010 1407.410 4.280 ;
        RECT 1408.250 0.010 1410.630 4.280 ;
        RECT 1411.470 0.010 1413.850 4.280 ;
        RECT 1414.690 0.010 1417.070 4.280 ;
        RECT 1417.910 0.010 1420.290 4.280 ;
        RECT 1421.130 0.010 1423.510 4.280 ;
        RECT 1424.350 0.010 1426.730 4.280 ;
        RECT 1427.570 0.010 1429.950 4.280 ;
        RECT 1430.790 0.010 1433.170 4.280 ;
        RECT 1434.010 0.010 1436.390 4.280 ;
        RECT 1437.230 0.010 1439.610 4.280 ;
        RECT 1440.450 0.010 1442.830 4.280 ;
        RECT 1443.670 0.010 1446.050 4.280 ;
        RECT 1446.890 0.010 1449.270 4.280 ;
        RECT 1450.110 0.010 1452.490 4.280 ;
        RECT 1453.330 0.010 1455.710 4.280 ;
        RECT 1456.550 0.010 1458.930 4.280 ;
        RECT 1459.770 0.010 1462.150 4.280 ;
        RECT 1462.990 0.010 1465.370 4.280 ;
        RECT 1466.210 0.010 1468.590 4.280 ;
        RECT 1469.430 0.010 1471.810 4.280 ;
        RECT 1472.650 0.010 1475.030 4.280 ;
        RECT 1475.870 0.010 1478.250 4.280 ;
        RECT 1479.090 0.010 1481.470 4.280 ;
        RECT 1482.310 0.010 1484.690 4.280 ;
        RECT 1485.530 0.010 1487.910 4.280 ;
        RECT 1488.750 0.010 1491.130 4.280 ;
        RECT 1491.970 0.010 1494.350 4.280 ;
        RECT 1495.190 0.010 1497.570 4.280 ;
        RECT 1498.410 0.010 1500.790 4.280 ;
        RECT 1501.630 0.010 1504.010 4.280 ;
        RECT 1504.850 0.010 1507.230 4.280 ;
        RECT 1508.070 0.010 1510.450 4.280 ;
        RECT 1511.290 0.010 1513.670 4.280 ;
        RECT 1514.510 0.010 1516.890 4.280 ;
        RECT 1517.730 0.010 1520.110 4.280 ;
        RECT 1520.950 0.010 1523.330 4.280 ;
        RECT 1524.170 0.010 1526.550 4.280 ;
        RECT 1527.390 0.010 1529.770 4.280 ;
        RECT 1530.610 0.010 1532.990 4.280 ;
        RECT 1533.830 0.010 1536.210 4.280 ;
        RECT 1537.050 0.010 1539.430 4.280 ;
        RECT 1540.270 0.010 1542.650 4.280 ;
        RECT 1543.490 0.010 1545.870 4.280 ;
        RECT 1546.710 0.010 1549.090 4.280 ;
        RECT 1549.930 0.010 1552.310 4.280 ;
        RECT 1553.150 0.010 1555.530 4.280 ;
        RECT 1556.370 0.010 1558.750 4.280 ;
        RECT 1559.590 0.010 1561.970 4.280 ;
        RECT 1562.810 0.010 1565.190 4.280 ;
        RECT 1566.030 0.010 1568.410 4.280 ;
        RECT 1569.250 0.010 1571.630 4.280 ;
        RECT 1572.470 0.010 1574.850 4.280 ;
        RECT 1575.690 0.010 1578.070 4.280 ;
        RECT 1578.910 0.010 1581.290 4.280 ;
        RECT 1582.130 0.010 1584.510 4.280 ;
        RECT 1585.350 0.010 1587.730 4.280 ;
        RECT 1588.570 0.010 1590.950 4.280 ;
        RECT 1591.790 0.010 1594.170 4.280 ;
        RECT 1595.010 0.010 1597.390 4.280 ;
        RECT 1598.230 0.010 1600.610 4.280 ;
        RECT 1601.450 0.010 1603.830 4.280 ;
        RECT 1604.670 0.010 1607.050 4.280 ;
        RECT 1607.890 0.010 1610.270 4.280 ;
        RECT 1611.110 0.010 1613.490 4.280 ;
        RECT 1614.330 0.010 1616.710 4.280 ;
        RECT 1617.550 0.010 1619.930 4.280 ;
        RECT 1620.770 0.010 1623.150 4.280 ;
        RECT 1623.990 0.010 1626.370 4.280 ;
        RECT 1627.210 0.010 1629.590 4.280 ;
        RECT 1630.430 0.010 1632.810 4.280 ;
        RECT 1633.650 0.010 1636.030 4.280 ;
        RECT 1636.870 0.010 1639.250 4.280 ;
        RECT 1640.090 0.010 1642.470 4.280 ;
        RECT 1643.310 0.010 1645.690 4.280 ;
        RECT 1646.530 0.010 1648.910 4.280 ;
        RECT 1649.750 0.010 1652.130 4.280 ;
        RECT 1652.970 0.010 1655.350 4.280 ;
        RECT 1656.190 0.010 1658.570 4.280 ;
        RECT 1659.410 0.010 1661.790 4.280 ;
        RECT 1662.630 0.010 1665.010 4.280 ;
        RECT 1665.850 0.010 1668.230 4.280 ;
        RECT 1669.070 0.010 1671.450 4.280 ;
        RECT 1672.290 0.010 1674.670 4.280 ;
        RECT 1675.510 0.010 1677.890 4.280 ;
        RECT 1678.730 0.010 1681.110 4.280 ;
        RECT 1681.950 0.010 1684.330 4.280 ;
        RECT 1685.170 0.010 1687.550 4.280 ;
        RECT 1688.390 0.010 1690.770 4.280 ;
        RECT 1691.610 0.010 1693.990 4.280 ;
        RECT 1694.830 0.010 1697.210 4.280 ;
        RECT 1698.050 0.010 1700.430 4.280 ;
        RECT 1701.270 0.010 1703.650 4.280 ;
        RECT 1704.490 0.010 1706.870 4.280 ;
        RECT 1707.710 0.010 1710.090 4.280 ;
        RECT 1710.930 0.010 1713.310 4.280 ;
        RECT 1714.150 0.010 1716.530 4.280 ;
        RECT 1717.370 0.010 1719.750 4.280 ;
        RECT 1720.590 0.010 1722.970 4.280 ;
        RECT 1723.810 0.010 1726.190 4.280 ;
        RECT 1727.030 0.010 1729.410 4.280 ;
        RECT 1730.250 0.010 1732.630 4.280 ;
        RECT 1733.470 0.010 1735.850 4.280 ;
        RECT 1736.690 0.010 1739.070 4.280 ;
        RECT 1739.910 0.010 1742.290 4.280 ;
        RECT 1743.130 0.010 1745.510 4.280 ;
        RECT 1746.350 0.010 1748.730 4.280 ;
        RECT 1749.570 0.010 1751.950 4.280 ;
        RECT 1752.790 0.010 1755.170 4.280 ;
        RECT 1756.010 0.010 1758.390 4.280 ;
        RECT 1759.230 0.010 1761.610 4.280 ;
        RECT 1762.450 0.010 1764.830 4.280 ;
        RECT 1765.670 0.010 1768.050 4.280 ;
        RECT 1768.890 0.010 1771.270 4.280 ;
        RECT 1772.110 0.010 1774.490 4.280 ;
        RECT 1775.330 0.010 1777.710 4.280 ;
        RECT 1778.550 0.010 1780.930 4.280 ;
        RECT 1781.770 0.010 1784.150 4.280 ;
        RECT 1784.990 0.010 1787.370 4.280 ;
        RECT 1788.210 0.010 1790.590 4.280 ;
        RECT 1791.430 0.010 1793.810 4.280 ;
        RECT 1794.650 0.010 1797.030 4.280 ;
        RECT 1797.870 0.010 1800.250 4.280 ;
        RECT 1801.090 0.010 1803.470 4.280 ;
        RECT 1804.310 0.010 1806.690 4.280 ;
        RECT 1807.530 0.010 1809.910 4.280 ;
        RECT 1810.750 0.010 1813.130 4.280 ;
        RECT 1813.970 0.010 1816.350 4.280 ;
        RECT 1817.190 0.010 1819.570 4.280 ;
        RECT 1820.410 0.010 1822.790 4.280 ;
        RECT 1823.630 0.010 1826.010 4.280 ;
        RECT 1826.850 0.010 1829.230 4.280 ;
        RECT 1830.070 0.010 1832.450 4.280 ;
        RECT 1833.290 0.010 1835.670 4.280 ;
        RECT 1836.510 0.010 1838.890 4.280 ;
        RECT 1839.730 0.010 1842.110 4.280 ;
        RECT 1842.950 0.010 1845.330 4.280 ;
        RECT 1846.170 0.010 1848.550 4.280 ;
        RECT 1849.390 0.010 1851.770 4.280 ;
        RECT 1852.610 0.010 1854.990 4.280 ;
        RECT 1855.830 0.010 1858.210 4.280 ;
        RECT 1859.050 0.010 1861.430 4.280 ;
        RECT 1862.270 0.010 1864.650 4.280 ;
        RECT 1865.490 0.010 1867.870 4.280 ;
        RECT 1868.710 0.010 1871.090 4.280 ;
        RECT 1871.930 0.010 1874.310 4.280 ;
        RECT 1875.150 0.010 1877.530 4.280 ;
        RECT 1878.370 0.010 1880.750 4.280 ;
        RECT 1881.590 0.010 1883.970 4.280 ;
        RECT 1884.810 0.010 1887.190 4.280 ;
        RECT 1888.030 0.010 1890.410 4.280 ;
        RECT 1891.250 0.010 1893.630 4.280 ;
        RECT 1894.470 0.010 1896.850 4.280 ;
        RECT 1897.690 0.010 1900.070 4.280 ;
        RECT 1900.910 0.010 1903.290 4.280 ;
        RECT 1904.130 0.010 1906.510 4.280 ;
        RECT 1907.350 0.010 1909.730 4.280 ;
        RECT 1910.570 0.010 1912.950 4.280 ;
        RECT 1913.790 0.010 1916.170 4.280 ;
        RECT 1917.010 0.010 1919.390 4.280 ;
        RECT 1920.230 0.010 1922.610 4.280 ;
        RECT 1923.450 0.010 1925.830 4.280 ;
        RECT 1926.670 0.010 1929.050 4.280 ;
        RECT 1929.890 0.010 1932.270 4.280 ;
        RECT 1933.110 0.010 1935.490 4.280 ;
        RECT 1936.330 0.010 1938.710 4.280 ;
        RECT 1939.550 0.010 1941.930 4.280 ;
        RECT 1942.770 0.010 1945.150 4.280 ;
        RECT 1945.990 0.010 1948.370 4.280 ;
        RECT 1949.210 0.010 1951.590 4.280 ;
        RECT 1952.430 0.010 1954.810 4.280 ;
        RECT 1955.650 0.010 1958.030 4.280 ;
        RECT 1958.870 0.010 1961.250 4.280 ;
        RECT 1962.090 0.010 1964.470 4.280 ;
        RECT 1965.310 0.010 1967.690 4.280 ;
        RECT 1968.530 0.010 1970.910 4.280 ;
        RECT 1971.750 0.010 1974.130 4.280 ;
        RECT 1974.970 0.010 1977.350 4.280 ;
        RECT 1978.190 0.010 1980.570 4.280 ;
        RECT 1981.410 0.010 1983.790 4.280 ;
        RECT 1984.630 0.010 1987.010 4.280 ;
        RECT 1987.850 0.010 1990.230 4.280 ;
        RECT 1991.070 0.010 1993.450 4.280 ;
        RECT 1994.290 0.010 1996.670 4.280 ;
        RECT 1997.510 0.010 1999.890 4.280 ;
        RECT 2000.730 0.010 2003.110 4.280 ;
        RECT 2003.950 0.010 2006.330 4.280 ;
        RECT 2007.170 0.010 2009.550 4.280 ;
        RECT 2010.390 0.010 2012.770 4.280 ;
        RECT 2013.610 0.010 2015.990 4.280 ;
        RECT 2016.830 0.010 2019.210 4.280 ;
        RECT 2020.050 0.010 2022.430 4.280 ;
        RECT 2023.270 0.010 2025.650 4.280 ;
        RECT 2026.490 0.010 2028.870 4.280 ;
        RECT 2029.710 0.010 2032.090 4.280 ;
        RECT 2032.930 0.010 2035.310 4.280 ;
        RECT 2036.150 0.010 2038.530 4.280 ;
        RECT 2039.370 0.010 2041.750 4.280 ;
        RECT 2042.590 0.010 2044.970 4.280 ;
        RECT 2045.810 0.010 2048.190 4.280 ;
        RECT 2049.030 0.010 2051.410 4.280 ;
        RECT 2052.250 0.010 2054.630 4.280 ;
        RECT 2055.470 0.010 2113.150 4.280 ;
      LAYER met3 ;
        RECT 25.130 151.320 2116.000 154.865 ;
        RECT 25.130 149.920 2115.600 151.320 ;
        RECT 25.130 140.440 2116.000 149.920 ;
        RECT 25.130 139.040 2115.600 140.440 ;
        RECT 25.130 129.560 2116.000 139.040 ;
        RECT 25.130 128.160 2115.600 129.560 ;
        RECT 25.130 118.680 2116.000 128.160 ;
        RECT 25.130 117.280 2115.600 118.680 ;
        RECT 25.130 107.800 2116.000 117.280 ;
        RECT 25.130 106.400 2115.600 107.800 ;
        RECT 25.130 96.920 2116.000 106.400 ;
        RECT 25.130 95.520 2115.600 96.920 ;
        RECT 25.130 86.040 2116.000 95.520 ;
        RECT 25.130 84.640 2115.600 86.040 ;
        RECT 25.130 75.160 2116.000 84.640 ;
        RECT 25.130 73.760 2115.600 75.160 ;
        RECT 25.130 64.280 2116.000 73.760 ;
        RECT 25.130 62.880 2115.600 64.280 ;
        RECT 25.130 53.400 2116.000 62.880 ;
        RECT 25.130 52.000 2115.600 53.400 ;
        RECT 25.130 42.520 2116.000 52.000 ;
        RECT 25.130 41.120 2115.600 42.520 ;
        RECT 25.130 31.640 2116.000 41.120 ;
        RECT 25.130 30.240 2115.600 31.640 ;
        RECT 25.130 20.760 2116.000 30.240 ;
        RECT 25.130 19.360 2115.600 20.760 ;
        RECT 25.130 9.880 2116.000 19.360 ;
        RECT 25.130 8.480 2115.600 9.880 ;
        RECT 25.130 0.175 2116.000 8.480 ;
      LAYER met4 ;
        RECT 290.095 4.800 325.670 152.825 ;
        RECT 327.370 4.800 333.870 152.825 ;
        RECT 335.570 4.800 354.770 152.825 ;
        RECT 356.470 4.800 362.570 152.825 ;
        RECT 364.270 4.800 383.870 152.825 ;
        RECT 385.570 4.800 400.920 152.825 ;
        RECT 402.620 4.800 404.770 152.825 ;
        RECT 406.470 4.800 437.820 152.825 ;
        RECT 439.520 4.800 476.170 152.825 ;
        RECT 477.870 4.800 513.070 152.825 ;
        RECT 514.770 4.800 551.420 152.825 ;
        RECT 553.120 4.800 588.320 152.825 ;
        RECT 590.020 4.800 626.670 152.825 ;
        RECT 628.370 4.800 663.570 152.825 ;
        RECT 665.270 4.800 701.920 152.825 ;
        RECT 703.620 4.800 706.020 152.825 ;
        RECT 707.720 4.800 738.820 152.825 ;
        RECT 740.520 4.800 742.920 152.825 ;
        RECT 744.620 4.800 777.170 152.825 ;
        RECT 778.870 4.800 781.270 152.825 ;
        RECT 782.970 4.800 814.070 152.825 ;
        RECT 815.770 4.800 818.170 152.825 ;
        RECT 819.870 4.800 852.420 152.825 ;
        RECT 854.120 4.800 856.520 152.825 ;
        RECT 858.220 4.800 889.320 152.825 ;
        RECT 891.020 4.800 893.420 152.825 ;
        RECT 895.120 4.800 927.670 152.825 ;
        RECT 929.370 4.800 931.770 152.825 ;
        RECT 933.470 4.800 964.570 152.825 ;
        RECT 966.270 4.800 968.670 152.825 ;
        RECT 970.370 4.800 1002.920 152.825 ;
        RECT 1004.620 4.800 1039.820 152.825 ;
        RECT 1041.520 4.800 1078.170 152.825 ;
        RECT 1079.870 4.800 1115.070 152.825 ;
        RECT 1116.770 4.800 1153.420 152.825 ;
        RECT 1155.120 4.800 1190.320 152.825 ;
        RECT 1192.020 4.800 1228.670 152.825 ;
        RECT 1230.370 4.800 1265.570 152.825 ;
        RECT 1267.270 4.800 1278.670 152.825 ;
        RECT 1280.370 4.800 1282.670 152.825 ;
        RECT 1284.370 4.800 1303.920 152.825 ;
        RECT 1305.620 4.800 1315.570 152.825 ;
        RECT 1317.270 4.800 1319.570 152.825 ;
        RECT 1321.270 4.800 1340.820 152.825 ;
        RECT 1342.520 4.800 1353.920 152.825 ;
        RECT 1355.620 4.800 1357.920 152.825 ;
        RECT 1359.620 4.800 1379.170 152.825 ;
        RECT 1380.870 4.800 1390.820 152.825 ;
        RECT 1392.520 4.800 1394.820 152.825 ;
        RECT 1396.520 4.800 1416.070 152.825 ;
        RECT 1417.770 4.800 1454.420 152.825 ;
        RECT 1456.120 4.800 1491.320 152.825 ;
        RECT 1493.020 4.800 1529.670 152.825 ;
        RECT 1531.370 4.800 1566.570 152.825 ;
        RECT 1568.270 4.800 1604.920 152.825 ;
        RECT 1606.620 4.800 1641.820 152.825 ;
        RECT 1643.520 4.800 1680.170 152.825 ;
        RECT 1681.870 4.800 1717.070 152.825 ;
        RECT 1718.770 4.800 1755.420 152.825 ;
        RECT 1757.120 4.800 1763.345 152.825 ;
        RECT 290.095 0.175 1763.345 4.800 ;
  END
END mgmt_protect
END LIBRARY

