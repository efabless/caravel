magic
tech sky130A
timestamp 1666994379
<< properties >>
string FIXED_BBOX 0 0 358800 518800
<< end >>
