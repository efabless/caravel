VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO manual_power_connections
  CLASS BLOCK ;
  FOREIGN manual_power_connections ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.100 BY 0.100 ;
  OBS
      LAYER met3 ;
        RECT 3048.235 4553.940 3140.235 4555.340 ;
        RECT 3053.000 4551.220 3134.300 4552.620 ;
        RECT 3081.800 4548.500 3128.300 4549.900 ;
        RECT 3077.000 4545.780 3122.300 4547.180 ;
        RECT 3072.250 4543.060 3116.300 4544.460 ;
        RECT 3067.300 4540.340 3110.300 4541.740 ;
        RECT 3062.500 4537.620 3104.300 4539.020 ;
        RECT 3057.800 4534.900 3098.300 4536.300 ;
        RECT 22.865 4529.460 114.865 4530.860 ;
        RECT 28.800 4526.740 110.100 4528.140 ;
        RECT 34.800 4524.020 81.300 4525.420 ;
        RECT 40.800 4521.300 86.100 4522.700 ;
        RECT 46.800 4518.580 90.850 4519.980 ;
        RECT 52.800 4515.860 95.800 4517.260 ;
        RECT 58.800 4513.140 100.600 4514.540 ;
        RECT 64.800 4510.420 105.300 4511.820 ;
        RECT 3048.235 4480.500 3140.235 4481.900 ;
        RECT 3053.000 4477.780 3134.300 4479.180 ;
        RECT 3081.800 4475.060 3128.300 4476.460 ;
        RECT 3077.000 4472.340 3122.300 4473.740 ;
        RECT 3072.250 4469.620 3116.300 4471.020 ;
        RECT 3067.300 4466.900 3110.300 4468.300 ;
        RECT 3062.500 4464.180 3104.300 4465.580 ;
        RECT 3057.800 4461.460 3098.300 4462.860 ;
        RECT 22.865 4456.020 114.865 4457.420 ;
        RECT 28.800 4453.300 110.100 4454.700 ;
        RECT 34.800 4450.580 81.300 4451.980 ;
        RECT 40.800 4447.860 86.100 4449.260 ;
        RECT 46.800 4445.140 90.850 4446.540 ;
        RECT 52.800 4442.420 95.800 4443.820 ;
        RECT 58.800 4439.700 100.600 4441.100 ;
        RECT 64.800 4436.980 105.300 4438.380 ;
        RECT 3048.235 4423.380 3140.235 4424.780 ;
        RECT 3053.000 4420.660 3134.300 4422.060 ;
        RECT 3081.800 4417.940 3128.300 4419.340 ;
        RECT 3077.000 4415.220 3122.300 4416.620 ;
        RECT 3072.250 4412.500 3116.300 4413.900 ;
        RECT 3067.300 4409.780 3110.300 4411.180 ;
        RECT 3062.500 4407.060 3104.300 4408.460 ;
        RECT 3057.800 4404.340 3098.300 4405.740 ;
        RECT 22.865 4390.740 114.865 4392.140 ;
        RECT 28.800 4388.020 110.100 4389.420 ;
        RECT 34.800 4385.300 81.300 4386.700 ;
        RECT 40.800 4382.580 86.100 4383.980 ;
        RECT 46.800 4379.860 90.850 4381.260 ;
        RECT 52.800 4377.140 95.800 4378.540 ;
        RECT 58.800 4374.420 100.600 4375.820 ;
        RECT 64.800 4371.700 105.300 4373.100 ;
        RECT 3048.235 4358.100 3140.235 4359.500 ;
        RECT 3053.000 4355.380 3134.300 4356.780 ;
        RECT 3081.800 4352.660 3128.300 4354.060 ;
        RECT 3077.000 4349.940 3122.300 4351.340 ;
        RECT 3072.250 4347.220 3116.300 4348.620 ;
        RECT 3067.300 4344.500 3110.300 4345.900 ;
        RECT 3062.500 4341.780 3104.300 4343.180 ;
        RECT 3057.800 4339.060 3098.300 4340.460 ;
        RECT 22.865 4325.460 114.865 4326.860 ;
        RECT 28.800 4322.740 110.100 4324.140 ;
        RECT 34.800 4320.020 81.300 4321.420 ;
        RECT 40.800 4317.300 86.100 4318.700 ;
        RECT 46.800 4314.580 90.850 4315.980 ;
        RECT 52.800 4311.860 95.800 4313.260 ;
        RECT 58.800 4309.140 100.600 4310.540 ;
        RECT 64.800 4306.420 105.300 4307.820 ;
        RECT 3048.235 4292.820 3140.235 4294.220 ;
        RECT 3053.000 4290.100 3134.300 4291.500 ;
        RECT 3081.800 4287.380 3128.300 4288.780 ;
        RECT 3077.000 4284.660 3122.300 4286.060 ;
        RECT 3072.250 4281.940 3116.300 4283.340 ;
        RECT 3067.300 4279.220 3110.300 4280.620 ;
        RECT 3062.500 4276.500 3104.300 4277.900 ;
        RECT 3057.800 4273.780 3098.300 4275.180 ;
        RECT 22.865 4260.180 114.865 4261.580 ;
        RECT 28.800 4257.460 110.100 4258.860 ;
        RECT 34.800 4254.740 81.300 4256.140 ;
        RECT 40.800 4252.020 86.100 4253.420 ;
        RECT 46.800 4249.300 90.850 4250.700 ;
        RECT 52.800 4246.580 95.800 4247.980 ;
        RECT 58.800 4243.860 100.600 4245.260 ;
        RECT 64.800 4241.140 105.300 4242.540 ;
        RECT 3048.235 4227.540 3140.235 4228.940 ;
        RECT 3053.000 4224.820 3134.300 4226.220 ;
        RECT 3081.800 4222.100 3128.300 4223.500 ;
        RECT 3077.000 4219.380 3122.300 4220.780 ;
        RECT 3072.250 4216.660 3116.300 4218.060 ;
        RECT 3067.300 4213.940 3110.300 4215.340 ;
        RECT 3062.500 4211.220 3104.300 4212.620 ;
        RECT 3057.800 4208.500 3098.300 4209.900 ;
        RECT 22.865 4194.900 114.865 4196.300 ;
        RECT 28.800 4192.180 110.100 4193.580 ;
        RECT 34.800 4189.460 81.300 4190.860 ;
        RECT 40.800 4186.740 86.100 4188.140 ;
        RECT 46.800 4184.020 90.850 4185.420 ;
        RECT 52.800 4181.300 95.800 4182.700 ;
        RECT 58.800 4178.580 100.600 4179.980 ;
        RECT 64.800 4175.860 105.300 4177.260 ;
        RECT 3048.235 4162.260 3140.235 4163.660 ;
        RECT 3053.000 4159.540 3134.300 4160.940 ;
        RECT 3081.800 4156.820 3128.300 4158.220 ;
        RECT 3077.000 4154.100 3122.300 4155.500 ;
        RECT 3072.250 4151.380 3116.300 4152.780 ;
        RECT 3067.300 4148.660 3110.300 4150.060 ;
        RECT 3062.500 4145.940 3104.300 4147.340 ;
        RECT 3057.800 4143.220 3098.300 4144.620 ;
        RECT 22.865 4129.620 114.865 4131.020 ;
        RECT 28.800 4126.900 110.100 4128.300 ;
        RECT 34.800 4124.180 81.300 4125.580 ;
        RECT 40.800 4121.460 86.100 4122.860 ;
        RECT 46.800 4118.740 90.850 4120.140 ;
        RECT 52.800 4116.020 95.800 4117.420 ;
        RECT 58.800 4113.300 100.600 4114.700 ;
        RECT 64.800 4110.580 105.300 4111.980 ;
        RECT 3048.235 4096.980 3140.235 4098.380 ;
        RECT 3053.000 4094.260 3134.300 4095.660 ;
        RECT 3081.800 4091.540 3128.300 4092.940 ;
        RECT 3077.000 4088.820 3122.300 4090.220 ;
        RECT 3072.250 4086.100 3116.300 4087.500 ;
        RECT 3067.300 4083.380 3110.300 4084.780 ;
        RECT 3062.500 4080.660 3104.300 4082.060 ;
        RECT 3057.800 4077.940 3098.300 4079.340 ;
        RECT 22.865 4064.340 114.865 4065.740 ;
        RECT 28.800 4061.620 110.100 4063.020 ;
        RECT 34.800 4058.900 81.300 4060.300 ;
        RECT 40.800 4056.180 86.100 4057.580 ;
        RECT 46.800 4053.460 90.850 4054.860 ;
        RECT 52.800 4050.740 95.800 4052.140 ;
        RECT 58.800 4048.020 100.600 4049.420 ;
        RECT 64.800 4045.300 105.300 4046.700 ;
        RECT 3048.235 4031.700 3140.235 4033.100 ;
        RECT 3053.000 4028.980 3134.300 4030.380 ;
        RECT 3081.800 4026.260 3128.300 4027.660 ;
        RECT 3077.000 4023.540 3122.300 4024.940 ;
        RECT 3072.250 4020.820 3116.300 4022.220 ;
        RECT 3067.300 4018.100 3110.300 4019.500 ;
        RECT 3062.500 4015.380 3104.300 4016.780 ;
        RECT 3057.800 4012.660 3098.300 4014.060 ;
        RECT 22.865 3999.060 114.865 4000.460 ;
        RECT 28.800 3996.340 110.100 3997.740 ;
        RECT 34.800 3993.620 81.300 3995.020 ;
        RECT 40.800 3990.900 86.100 3992.300 ;
        RECT 46.800 3988.180 90.850 3989.580 ;
        RECT 52.800 3985.460 95.800 3986.860 ;
        RECT 58.800 3982.740 100.600 3984.140 ;
        RECT 64.800 3980.020 105.300 3981.420 ;
        RECT 3048.235 3966.420 3140.235 3967.820 ;
        RECT 3053.000 3963.700 3134.300 3965.100 ;
        RECT 3081.800 3960.980 3128.300 3962.380 ;
        RECT 3077.000 3958.260 3122.300 3959.660 ;
        RECT 3072.250 3955.540 3116.300 3956.940 ;
        RECT 3067.300 3952.820 3110.300 3954.220 ;
        RECT 3062.500 3950.100 3104.300 3951.500 ;
        RECT 3057.800 3947.380 3098.300 3948.780 ;
        RECT 22.865 3933.780 114.865 3935.180 ;
        RECT 28.800 3931.060 110.100 3932.460 ;
        RECT 34.800 3928.340 81.300 3929.740 ;
        RECT 40.800 3925.620 86.100 3927.020 ;
        RECT 46.800 3922.900 90.850 3924.300 ;
        RECT 52.800 3920.180 95.800 3921.580 ;
        RECT 58.800 3917.460 100.600 3918.860 ;
        RECT 64.800 3914.740 105.300 3916.140 ;
        RECT 3048.235 3901.140 3140.235 3902.540 ;
        RECT 3053.000 3898.420 3134.300 3899.820 ;
        RECT 3081.800 3895.700 3128.300 3897.100 ;
        RECT 3077.000 3892.980 3122.300 3894.380 ;
        RECT 3072.250 3890.260 3116.300 3891.660 ;
        RECT 3067.300 3887.540 3110.300 3888.940 ;
        RECT 3062.500 3884.820 3104.300 3886.220 ;
        RECT 3057.800 3882.100 3098.300 3883.500 ;
        RECT 22.865 3868.500 114.865 3869.900 ;
        RECT 28.800 3865.780 110.100 3867.180 ;
        RECT 34.800 3863.060 81.300 3864.460 ;
        RECT 40.800 3860.340 86.100 3861.740 ;
        RECT 46.800 3857.620 90.850 3859.020 ;
        RECT 52.800 3854.900 95.800 3856.300 ;
        RECT 58.800 3852.180 100.600 3853.580 ;
        RECT 64.800 3849.460 105.300 3850.860 ;
        RECT 3048.235 3835.860 3140.235 3837.260 ;
        RECT 3053.000 3833.140 3134.300 3834.540 ;
        RECT 3081.800 3830.420 3128.300 3831.820 ;
        RECT 3077.000 3827.700 3122.300 3829.100 ;
        RECT 3072.250 3824.980 3116.300 3826.380 ;
        RECT 3067.300 3822.260 3110.300 3823.660 ;
        RECT 3062.500 3819.540 3104.300 3820.940 ;
        RECT 3057.800 3816.820 3098.300 3818.220 ;
        RECT 22.865 3803.220 114.865 3804.620 ;
        RECT 28.800 3800.500 110.100 3801.900 ;
        RECT 34.800 3797.780 81.300 3799.180 ;
        RECT 40.800 3795.060 86.100 3796.460 ;
        RECT 46.800 3792.340 90.850 3793.740 ;
        RECT 52.800 3789.620 95.800 3791.020 ;
        RECT 58.800 3786.900 100.600 3788.300 ;
        RECT 64.800 3784.180 105.300 3785.580 ;
        RECT 3048.235 3770.580 3140.235 3771.980 ;
        RECT 3053.000 3767.860 3134.300 3769.260 ;
        RECT 3081.800 3765.140 3128.300 3766.540 ;
        RECT 3077.000 3762.420 3122.300 3763.820 ;
        RECT 3072.250 3759.700 3116.300 3761.100 ;
        RECT 3067.300 3756.980 3110.300 3758.380 ;
        RECT 3062.500 3754.260 3104.300 3755.660 ;
        RECT 3057.800 3751.540 3098.300 3752.940 ;
        RECT 22.865 3737.940 114.865 3739.340 ;
        RECT 28.800 3735.220 110.100 3736.620 ;
        RECT 34.800 3732.500 81.300 3733.900 ;
        RECT 40.800 3729.780 86.100 3731.180 ;
        RECT 46.800 3727.060 90.850 3728.460 ;
        RECT 52.800 3724.340 95.800 3725.740 ;
        RECT 58.800 3721.620 100.600 3723.020 ;
        RECT 64.800 3718.900 105.300 3720.300 ;
        RECT 3048.235 3705.300 3140.235 3706.700 ;
        RECT 3053.000 3702.580 3134.300 3703.980 ;
        RECT 3081.800 3699.860 3128.300 3701.260 ;
        RECT 3077.000 3697.140 3122.300 3698.540 ;
        RECT 3072.250 3694.420 3116.300 3695.820 ;
        RECT 3067.300 3691.700 3110.300 3693.100 ;
        RECT 3062.500 3688.980 3104.300 3690.380 ;
        RECT 3057.800 3686.260 3098.300 3687.660 ;
        RECT 22.865 3680.820 114.865 3682.220 ;
        RECT 28.800 3678.100 110.100 3679.500 ;
        RECT 34.800 3675.380 81.300 3676.780 ;
        RECT 40.800 3672.660 86.100 3674.060 ;
        RECT 46.800 3669.940 90.850 3671.340 ;
        RECT 52.800 3667.220 95.800 3668.620 ;
        RECT 58.800 3664.500 100.600 3665.900 ;
        RECT 64.800 3661.780 105.300 3663.180 ;
        RECT 3048.235 3640.020 3140.235 3641.420 ;
        RECT 3053.000 3637.300 3134.300 3638.700 ;
        RECT 3081.800 3634.580 3128.300 3635.980 ;
        RECT 3077.000 3631.860 3122.300 3633.260 ;
        RECT 3072.250 3629.140 3116.300 3630.540 ;
        RECT 3067.300 3626.420 3110.300 3627.820 ;
        RECT 3062.500 3623.700 3104.300 3625.100 ;
        RECT 3057.800 3620.980 3098.300 3622.380 ;
        RECT 22.865 3607.380 114.865 3608.780 ;
        RECT 28.800 3604.660 110.100 3606.060 ;
        RECT 34.800 3601.940 81.300 3603.340 ;
        RECT 40.800 3599.220 86.100 3600.620 ;
        RECT 46.800 3596.500 90.850 3597.900 ;
        RECT 52.800 3593.780 95.800 3595.180 ;
        RECT 58.800 3591.060 100.600 3592.460 ;
        RECT 64.800 3588.340 105.300 3589.740 ;
        RECT 3048.235 3566.580 3140.235 3567.980 ;
        RECT 3053.000 3563.860 3134.300 3565.260 ;
        RECT 3081.800 3561.140 3128.300 3562.540 ;
        RECT 3077.000 3558.420 3122.300 3559.820 ;
        RECT 3072.250 3555.700 3116.300 3557.100 ;
        RECT 3067.300 3552.980 3110.300 3554.380 ;
        RECT 3062.500 3550.260 3104.300 3551.660 ;
        RECT 3057.800 3547.540 3098.300 3548.940 ;
        RECT 22.865 3542.100 114.865 3543.500 ;
        RECT 28.800 3539.380 110.100 3540.780 ;
        RECT 34.800 3536.660 81.300 3538.060 ;
        RECT 40.800 3533.940 86.100 3535.340 ;
        RECT 46.800 3531.220 90.850 3532.620 ;
        RECT 52.800 3528.500 95.800 3529.900 ;
        RECT 58.800 3525.780 100.600 3527.180 ;
        RECT 64.800 3523.060 105.300 3524.460 ;
        RECT 3048.235 3509.460 3140.235 3510.860 ;
        RECT 3053.000 3506.740 3134.300 3508.140 ;
        RECT 3081.800 3504.020 3128.300 3505.420 ;
        RECT 3077.000 3501.300 3122.300 3502.700 ;
        RECT 3072.250 3498.580 3116.300 3499.980 ;
        RECT 3067.300 3495.860 3110.300 3497.260 ;
        RECT 3062.500 3493.140 3104.300 3494.540 ;
        RECT 3057.800 3490.420 3098.300 3491.820 ;
        RECT 22.865 3460.500 114.865 3461.900 ;
        RECT 28.800 3457.780 110.100 3459.180 ;
        RECT 34.800 3455.060 81.300 3456.460 ;
        RECT 40.800 3452.340 86.100 3453.740 ;
        RECT 46.800 3449.620 90.850 3451.020 ;
        RECT 52.800 3446.900 95.800 3448.300 ;
        RECT 58.800 3444.180 100.600 3445.580 ;
        RECT 3048.235 3444.180 3140.235 3445.580 ;
        RECT 64.800 3441.460 105.300 3442.860 ;
        RECT 3053.000 3441.460 3134.300 3442.860 ;
        RECT 3081.800 3438.740 3128.300 3440.140 ;
        RECT 3077.000 3436.020 3122.300 3437.420 ;
        RECT 3072.250 3433.300 3116.300 3434.700 ;
        RECT 3067.300 3430.580 3110.300 3431.980 ;
        RECT 3062.500 3427.860 3104.300 3429.260 ;
        RECT 3057.800 3425.140 3098.300 3426.540 ;
        RECT 22.865 3411.540 114.865 3412.940 ;
        RECT 28.800 3408.820 110.100 3410.220 ;
        RECT 34.800 3406.100 81.300 3407.500 ;
        RECT 40.800 3403.380 86.100 3404.780 ;
        RECT 46.800 3400.660 90.850 3402.060 ;
        RECT 52.800 3397.940 95.800 3399.340 ;
        RECT 58.800 3395.220 100.600 3396.620 ;
        RECT 64.800 3392.500 105.300 3393.900 ;
        RECT 3048.235 3378.900 3140.235 3380.300 ;
        RECT 3053.000 3376.180 3134.300 3377.580 ;
        RECT 3081.800 3373.460 3128.300 3374.860 ;
        RECT 3077.000 3370.740 3122.300 3372.140 ;
        RECT 3072.250 3368.020 3116.300 3369.420 ;
        RECT 3067.300 3365.300 3110.300 3366.700 ;
        RECT 3062.500 3362.580 3104.300 3363.980 ;
        RECT 3057.800 3359.860 3098.300 3361.260 ;
        RECT 22.865 3346.260 114.865 3347.660 ;
        RECT 28.800 3343.540 110.100 3344.940 ;
        RECT 34.800 3340.820 81.300 3342.220 ;
        RECT 40.800 3338.100 86.100 3339.500 ;
        RECT 46.800 3335.380 90.850 3336.780 ;
        RECT 52.800 3332.660 95.800 3334.060 ;
        RECT 58.800 3329.940 100.600 3331.340 ;
        RECT 64.800 3327.220 105.300 3328.620 ;
        RECT 3048.235 3313.620 3140.235 3315.020 ;
        RECT 3053.000 3310.900 3134.300 3312.300 ;
        RECT 3081.800 3308.180 3128.300 3309.580 ;
        RECT 3077.000 3305.460 3122.300 3306.860 ;
        RECT 3072.250 3302.740 3116.300 3304.140 ;
        RECT 3067.300 3300.020 3110.300 3301.420 ;
        RECT 3062.500 3297.300 3104.300 3298.700 ;
        RECT 3057.800 3294.580 3098.300 3295.980 ;
        RECT 22.865 3280.980 114.865 3282.380 ;
        RECT 28.800 3278.260 110.100 3279.660 ;
        RECT 34.800 3275.540 81.300 3276.940 ;
        RECT 40.800 3272.820 86.100 3274.220 ;
        RECT 46.800 3270.100 90.850 3271.500 ;
        RECT 52.800 3267.380 95.800 3268.780 ;
        RECT 58.800 3264.660 100.600 3266.060 ;
        RECT 64.800 3261.940 105.300 3263.340 ;
        RECT 3048.235 3248.340 3140.235 3249.740 ;
        RECT 3053.000 3245.620 3134.300 3247.020 ;
        RECT 3081.800 3242.900 3128.300 3244.300 ;
        RECT 3077.000 3240.180 3122.300 3241.580 ;
        RECT 3072.250 3237.460 3116.300 3238.860 ;
        RECT 3067.300 3234.740 3110.300 3236.140 ;
        RECT 3062.500 3232.020 3104.300 3233.420 ;
        RECT 3057.800 3229.300 3098.300 3230.700 ;
        RECT 22.865 3207.540 114.865 3208.940 ;
        RECT 28.800 3204.820 110.100 3206.220 ;
        RECT 34.800 3202.100 81.300 3203.500 ;
        RECT 40.800 3199.380 86.100 3200.780 ;
        RECT 46.800 3196.660 90.850 3198.060 ;
        RECT 52.800 3193.940 95.800 3195.340 ;
        RECT 58.800 3191.220 100.600 3192.620 ;
        RECT 64.800 3188.500 105.300 3189.900 ;
        RECT 3048.235 3183.060 3140.235 3184.460 ;
        RECT 3053.000 3180.340 3134.300 3181.740 ;
        RECT 3081.800 3177.620 3128.300 3179.020 ;
        RECT 3077.000 3174.900 3122.300 3176.300 ;
        RECT 3072.250 3172.180 3116.300 3173.580 ;
        RECT 3067.300 3169.460 3110.300 3170.860 ;
        RECT 3062.500 3166.740 3104.300 3168.140 ;
        RECT 3057.800 3164.020 3098.300 3165.420 ;
        RECT 22.865 3150.420 114.865 3151.820 ;
        RECT 28.800 3147.700 110.100 3149.100 ;
        RECT 34.800 3144.980 81.300 3146.380 ;
        RECT 40.800 3142.260 86.100 3143.660 ;
        RECT 46.800 3139.540 90.850 3140.940 ;
        RECT 52.800 3136.820 95.800 3138.220 ;
        RECT 58.800 3134.100 100.600 3135.500 ;
        RECT 64.800 3131.380 105.300 3132.780 ;
        RECT 3048.235 3117.780 3140.235 3119.180 ;
        RECT 3053.000 3115.060 3134.300 3116.460 ;
        RECT 3081.800 3112.340 3128.300 3113.740 ;
        RECT 3077.000 3109.620 3122.300 3111.020 ;
        RECT 3072.250 3106.900 3116.300 3108.300 ;
        RECT 3067.300 3104.180 3110.300 3105.580 ;
        RECT 3062.500 3101.460 3104.300 3102.860 ;
        RECT 3057.800 3098.740 3098.300 3100.140 ;
        RECT 22.865 3085.140 114.865 3086.540 ;
        RECT 28.800 3082.420 110.100 3083.820 ;
        RECT 34.800 3079.700 81.300 3081.100 ;
        RECT 40.800 3076.980 86.100 3078.380 ;
        RECT 46.800 3074.260 90.850 3075.660 ;
        RECT 52.800 3071.540 95.800 3072.940 ;
        RECT 58.800 3068.820 100.600 3070.220 ;
        RECT 64.800 3066.100 105.300 3067.500 ;
        RECT 3048.235 3052.500 3140.235 3053.900 ;
        RECT 3053.000 3049.780 3134.300 3051.180 ;
        RECT 3081.800 3047.060 3128.300 3048.460 ;
        RECT 3077.000 3044.340 3122.300 3045.740 ;
        RECT 3072.250 3041.620 3116.300 3043.020 ;
        RECT 3067.300 3038.900 3110.300 3040.300 ;
        RECT 3062.500 3036.180 3104.300 3037.580 ;
        RECT 3057.800 3033.460 3098.300 3034.860 ;
        RECT 22.865 3030.740 114.865 3032.140 ;
        RECT 28.800 3028.020 110.100 3029.420 ;
        RECT 34.800 3025.300 81.300 3026.700 ;
        RECT 40.800 3022.580 86.100 3023.980 ;
        RECT 46.800 3019.860 90.850 3021.260 ;
        RECT 52.800 3017.140 95.800 3018.540 ;
        RECT 58.800 3014.420 100.600 3015.820 ;
        RECT 64.800 3011.700 105.300 3013.100 ;
        RECT 3048.235 2987.220 3140.235 2988.620 ;
        RECT 3053.000 2984.500 3134.300 2985.900 ;
        RECT 3081.800 2981.780 3128.300 2983.180 ;
        RECT 3077.000 2979.060 3122.300 2980.460 ;
        RECT 3072.250 2976.340 3116.300 2977.740 ;
        RECT 3067.300 2973.620 3110.300 2975.020 ;
        RECT 3062.500 2970.900 3104.300 2972.300 ;
        RECT 3057.800 2968.180 3098.300 2969.580 ;
        RECT 22.865 2954.580 114.865 2955.980 ;
        RECT 28.800 2951.860 110.100 2953.260 ;
        RECT 34.800 2949.140 81.300 2950.540 ;
        RECT 40.800 2946.420 86.100 2947.820 ;
        RECT 46.800 2943.700 90.850 2945.100 ;
        RECT 52.800 2940.980 95.800 2942.380 ;
        RECT 58.800 2938.260 100.600 2939.660 ;
        RECT 64.800 2935.540 105.300 2936.940 ;
        RECT 3048.235 2921.940 3140.235 2923.340 ;
        RECT 3053.000 2919.220 3134.300 2920.620 ;
        RECT 3081.800 2916.500 3128.300 2917.900 ;
        RECT 3077.000 2913.780 3122.300 2915.180 ;
        RECT 3072.250 2911.060 3116.300 2912.460 ;
        RECT 3067.300 2908.340 3110.300 2909.740 ;
        RECT 3062.500 2905.620 3104.300 2907.020 ;
        RECT 3057.800 2902.900 3098.300 2904.300 ;
        RECT 22.865 2889.300 114.865 2890.700 ;
        RECT 28.800 2886.580 110.100 2887.980 ;
        RECT 34.800 2883.860 81.300 2885.260 ;
        RECT 40.800 2881.140 86.100 2882.540 ;
        RECT 46.800 2878.420 90.850 2879.820 ;
        RECT 52.800 2875.700 95.800 2877.100 ;
        RECT 58.800 2872.980 100.600 2874.380 ;
        RECT 64.800 2870.260 105.300 2871.660 ;
        RECT 3048.235 2856.660 3140.235 2858.060 ;
        RECT 3053.000 2853.940 3134.300 2855.340 ;
        RECT 3081.800 2851.220 3128.300 2852.620 ;
        RECT 3077.000 2848.500 3122.300 2849.900 ;
        RECT 3072.250 2845.780 3116.300 2847.180 ;
        RECT 3067.300 2843.060 3110.300 2844.460 ;
        RECT 3062.500 2840.340 3104.300 2841.740 ;
        RECT 3057.800 2837.620 3098.300 2839.020 ;
        RECT 22.865 2834.900 114.865 2836.300 ;
        RECT 28.800 2832.180 110.100 2833.580 ;
        RECT 34.800 2829.460 81.300 2830.860 ;
        RECT 40.800 2826.740 86.100 2828.140 ;
        RECT 46.800 2824.020 90.850 2825.420 ;
        RECT 52.800 2821.300 95.800 2822.700 ;
        RECT 58.800 2818.580 100.600 2819.980 ;
        RECT 64.800 2815.860 105.300 2817.260 ;
        RECT 3048.235 2791.380 3140.235 2792.780 ;
        RECT 3053.000 2788.660 3134.300 2790.060 ;
        RECT 3081.800 2785.940 3128.300 2787.340 ;
        RECT 3077.000 2783.220 3122.300 2784.620 ;
        RECT 3072.250 2780.500 3116.300 2781.900 ;
        RECT 3067.300 2777.780 3110.300 2779.180 ;
        RECT 3062.500 2775.060 3104.300 2776.460 ;
        RECT 3057.800 2772.340 3098.300 2773.740 ;
        RECT 22.865 2758.740 114.865 2760.140 ;
        RECT 28.800 2756.020 110.100 2757.420 ;
        RECT 34.800 2753.300 81.300 2754.700 ;
        RECT 40.800 2750.580 86.100 2751.980 ;
        RECT 46.800 2747.860 90.850 2749.260 ;
        RECT 52.800 2745.140 95.800 2746.540 ;
        RECT 58.800 2742.420 100.600 2743.820 ;
        RECT 64.800 2739.700 105.300 2741.100 ;
        RECT 3072.250 2715.220 3116.300 2716.620 ;
        RECT 3067.300 2712.500 3110.300 2713.900 ;
        RECT 3062.500 2709.780 3104.300 2711.180 ;
        RECT 3057.800 2707.060 3098.300 2708.460 ;
        RECT 22.865 2693.460 114.865 2694.860 ;
        RECT 28.800 2690.740 110.100 2692.140 ;
        RECT 34.800 2688.020 81.300 2689.420 ;
        RECT 40.800 2685.300 86.100 2686.700 ;
        RECT 46.800 2682.580 90.850 2683.980 ;
        RECT 52.800 2679.860 95.800 2681.260 ;
        RECT 58.800 2677.140 100.600 2678.540 ;
        RECT 64.800 2674.420 105.300 2675.820 ;
        RECT 3048.235 2652.660 3140.235 2654.060 ;
        RECT 3053.000 2649.940 3134.300 2651.340 ;
        RECT 3081.800 2647.220 3128.300 2648.620 ;
        RECT 3077.000 2644.500 3122.300 2645.900 ;
        RECT 3072.250 2641.780 3116.300 2643.180 ;
        RECT 3067.300 2639.060 3110.300 2640.460 ;
        RECT 3062.500 2636.340 3104.300 2637.740 ;
        RECT 3057.800 2633.620 3098.300 2635.020 ;
        RECT 22.865 2628.180 114.865 2629.580 ;
        RECT 28.800 2625.460 110.100 2626.860 ;
        RECT 34.800 2622.740 81.300 2624.140 ;
        RECT 40.800 2620.020 86.100 2621.420 ;
        RECT 46.800 2617.300 90.850 2618.700 ;
        RECT 52.800 2614.580 95.800 2615.980 ;
        RECT 58.800 2611.860 100.600 2613.260 ;
        RECT 64.800 2609.140 105.300 2610.540 ;
        RECT 3048.235 2587.380 3140.235 2588.780 ;
        RECT 3053.000 2584.660 3134.300 2586.060 ;
        RECT 3081.800 2581.940 3128.300 2583.340 ;
        RECT 3077.000 2579.220 3122.300 2580.620 ;
        RECT 3072.250 2576.500 3116.300 2577.900 ;
        RECT 3067.300 2573.780 3110.300 2575.180 ;
        RECT 3062.500 2571.060 3104.300 2572.460 ;
        RECT 3057.800 2568.340 3098.300 2569.740 ;
        RECT 22.865 2562.900 114.865 2564.300 ;
        RECT 28.800 2560.180 110.100 2561.580 ;
        RECT 34.800 2557.460 81.300 2558.860 ;
        RECT 40.800 2554.740 86.100 2556.140 ;
        RECT 46.800 2552.020 90.850 2553.420 ;
        RECT 52.800 2549.300 95.800 2550.700 ;
        RECT 58.800 2546.580 100.600 2547.980 ;
        RECT 64.800 2543.860 105.300 2545.260 ;
        RECT 3048.235 2522.100 3140.235 2523.500 ;
        RECT 3053.000 2519.380 3134.300 2520.780 ;
        RECT 3081.800 2516.660 3128.300 2518.060 ;
        RECT 3077.000 2513.940 3122.300 2515.340 ;
        RECT 3072.250 2511.220 3116.300 2512.620 ;
        RECT 3067.300 2508.500 3110.300 2509.900 ;
        RECT 3062.500 2505.780 3104.300 2507.180 ;
        RECT 3057.800 2503.060 3098.300 2504.460 ;
        RECT 22.865 2497.620 114.865 2499.020 ;
        RECT 28.800 2494.900 110.100 2496.300 ;
        RECT 34.800 2492.180 81.300 2493.580 ;
        RECT 40.800 2489.460 86.100 2490.860 ;
        RECT 46.800 2486.740 90.850 2488.140 ;
        RECT 52.800 2484.020 95.800 2485.420 ;
        RECT 58.800 2481.300 100.600 2482.700 ;
        RECT 64.800 2478.580 105.300 2479.980 ;
        RECT 3048.235 2456.820 3140.235 2458.220 ;
        RECT 3053.000 2454.100 3134.300 2455.500 ;
        RECT 3081.800 2451.380 3128.300 2452.780 ;
        RECT 3077.000 2448.660 3122.300 2450.060 ;
        RECT 3072.250 2445.940 3116.300 2447.340 ;
        RECT 3067.300 2443.220 3110.300 2444.620 ;
        RECT 3062.500 2440.500 3104.300 2441.900 ;
        RECT 3057.800 2437.780 3098.300 2439.180 ;
        RECT 22.865 2432.340 114.865 2433.740 ;
        RECT 28.800 2429.620 110.100 2431.020 ;
        RECT 34.800 2426.900 81.300 2428.300 ;
        RECT 40.800 2424.180 86.100 2425.580 ;
        RECT 46.800 2421.460 90.850 2422.860 ;
        RECT 52.800 2418.740 95.800 2420.140 ;
        RECT 58.800 2416.020 100.600 2417.420 ;
        RECT 64.800 2413.300 105.300 2414.700 ;
        RECT 3048.235 2383.380 3140.235 2384.780 ;
        RECT 3053.000 2380.660 3134.300 2382.060 ;
        RECT 3081.800 2377.940 3128.300 2379.340 ;
        RECT 3077.000 2375.220 3122.300 2376.620 ;
        RECT 3072.250 2372.500 3116.300 2373.900 ;
        RECT 3067.300 2369.780 3110.300 2371.180 ;
        RECT 3062.500 2367.060 3104.300 2368.460 ;
        RECT 3057.800 2364.340 3098.300 2365.740 ;
        RECT 22.865 2356.180 114.865 2357.580 ;
        RECT 28.800 2353.460 110.100 2354.860 ;
        RECT 34.800 2350.740 81.300 2352.140 ;
        RECT 40.800 2348.020 86.100 2349.420 ;
        RECT 46.800 2345.300 90.850 2346.700 ;
        RECT 52.800 2342.580 95.800 2343.980 ;
        RECT 58.800 2339.860 100.600 2341.260 ;
        RECT 64.800 2337.140 105.300 2338.540 ;
        RECT 3048.235 2318.100 3140.235 2319.500 ;
        RECT 3053.000 2315.380 3134.300 2316.780 ;
        RECT 3081.800 2312.660 3128.300 2314.060 ;
        RECT 3077.000 2309.940 3122.300 2311.340 ;
        RECT 3072.250 2307.220 3116.300 2308.620 ;
        RECT 3067.300 2304.500 3110.300 2305.900 ;
        RECT 22.865 2301.780 114.865 2303.180 ;
        RECT 3062.500 2301.780 3104.300 2303.180 ;
        RECT 28.800 2299.060 110.100 2300.460 ;
        RECT 3057.800 2299.060 3098.300 2300.460 ;
        RECT 34.800 2296.340 81.300 2297.740 ;
        RECT 40.800 2293.620 86.100 2295.020 ;
        RECT 46.800 2290.900 90.850 2292.300 ;
        RECT 52.800 2288.180 95.800 2289.580 ;
        RECT 58.800 2285.460 100.600 2286.860 ;
        RECT 64.800 2282.740 105.300 2284.140 ;
        RECT 3048.235 2252.820 3140.235 2254.220 ;
        RECT 3053.000 2250.100 3134.300 2251.500 ;
        RECT 3081.800 2247.380 3128.300 2248.780 ;
        RECT 3077.000 2244.660 3122.300 2246.060 ;
        RECT 3072.250 2241.940 3116.300 2243.340 ;
        RECT 3067.300 2239.220 3110.300 2240.620 ;
        RECT 22.865 2236.500 114.865 2237.900 ;
        RECT 3062.500 2236.500 3104.300 2237.900 ;
        RECT 28.800 2233.780 110.100 2235.180 ;
        RECT 3057.800 2233.780 3098.300 2235.180 ;
        RECT 34.800 2231.060 81.300 2232.460 ;
        RECT 40.800 2228.340 86.100 2229.740 ;
        RECT 46.800 2225.620 90.850 2227.020 ;
        RECT 52.800 2222.900 95.800 2224.300 ;
        RECT 58.800 2220.180 100.600 2221.580 ;
        RECT 64.800 2217.460 105.300 2218.860 ;
        RECT 3048.235 2187.540 3140.235 2188.940 ;
        RECT 3053.000 2184.820 3134.300 2186.220 ;
        RECT 3081.800 2182.100 3128.300 2183.500 ;
        RECT 3077.000 2179.380 3122.300 2180.780 ;
        RECT 3072.250 2176.660 3116.300 2178.060 ;
        RECT 3067.300 2173.940 3110.300 2175.340 ;
        RECT 22.865 2171.220 114.865 2172.620 ;
        RECT 3062.500 2171.220 3104.300 2172.620 ;
        RECT 28.800 2168.500 110.100 2169.900 ;
        RECT 3057.800 2168.500 3098.300 2169.900 ;
        RECT 34.800 2165.780 81.300 2167.180 ;
        RECT 40.800 2163.060 86.100 2164.460 ;
        RECT 46.800 2160.340 90.850 2161.740 ;
        RECT 52.800 2157.620 95.800 2159.020 ;
        RECT 58.800 2154.900 100.600 2156.300 ;
        RECT 64.800 2152.180 105.300 2153.580 ;
        RECT 3048.235 2122.260 3140.235 2123.660 ;
        RECT 3053.000 2119.540 3134.300 2120.940 ;
        RECT 3081.800 2116.820 3128.300 2118.220 ;
        RECT 3077.000 2114.100 3122.300 2115.500 ;
        RECT 3072.250 2111.380 3116.300 2112.780 ;
        RECT 3067.300 2108.660 3110.300 2110.060 ;
        RECT 22.865 2105.940 114.865 2107.340 ;
        RECT 3062.500 2105.940 3104.300 2107.340 ;
        RECT 28.800 2103.220 110.100 2104.620 ;
        RECT 3057.800 2103.220 3098.300 2104.620 ;
        RECT 34.800 2100.500 81.300 2101.900 ;
        RECT 40.800 2097.780 86.100 2099.180 ;
        RECT 46.800 2095.060 90.850 2096.460 ;
        RECT 52.800 2092.340 95.800 2093.740 ;
        RECT 58.800 2089.620 100.600 2091.020 ;
        RECT 64.800 2086.900 105.300 2088.300 ;
        RECT 3048.235 2056.980 3140.235 2058.380 ;
        RECT 3053.000 2054.260 3134.300 2055.660 ;
        RECT 3081.800 2051.540 3128.300 2052.940 ;
        RECT 3077.000 2048.820 3122.300 2050.220 ;
        RECT 3072.250 2046.100 3116.300 2047.500 ;
        RECT 3067.300 2043.380 3110.300 2044.780 ;
        RECT 22.865 2040.660 114.865 2042.060 ;
        RECT 3062.500 2040.660 3104.300 2042.060 ;
        RECT 28.800 2037.940 110.100 2039.340 ;
        RECT 3057.800 2037.940 3098.300 2039.340 ;
        RECT 34.800 2035.220 81.300 2036.620 ;
        RECT 40.800 2032.500 86.100 2033.900 ;
        RECT 46.800 2029.780 90.850 2031.180 ;
        RECT 52.800 2027.060 95.800 2028.460 ;
        RECT 58.800 2024.340 100.600 2025.740 ;
        RECT 64.800 2021.620 105.300 2023.020 ;
        RECT 3048.235 1991.700 3140.235 1993.100 ;
        RECT 3053.000 1988.980 3134.300 1990.380 ;
        RECT 3081.800 1986.260 3128.300 1987.660 ;
        RECT 3077.000 1983.540 3122.300 1984.940 ;
        RECT 3072.250 1980.820 3116.300 1982.220 ;
        RECT 3067.300 1978.100 3110.300 1979.500 ;
        RECT 22.865 1975.380 114.865 1976.780 ;
        RECT 3062.500 1975.380 3104.300 1976.780 ;
        RECT 28.800 1972.660 110.100 1974.060 ;
        RECT 3057.800 1972.660 3098.300 1974.060 ;
        RECT 34.800 1969.940 81.300 1971.340 ;
        RECT 40.800 1967.220 86.100 1968.620 ;
        RECT 46.800 1964.500 90.850 1965.900 ;
        RECT 52.800 1961.780 95.800 1963.180 ;
        RECT 58.800 1959.060 100.600 1960.460 ;
        RECT 64.800 1956.340 105.300 1957.740 ;
        RECT 3048.235 1926.420 3140.235 1927.820 ;
        RECT 3053.000 1923.700 3134.300 1925.100 ;
        RECT 3081.800 1920.980 3128.300 1922.380 ;
        RECT 3077.000 1918.260 3122.300 1919.660 ;
        RECT 3072.250 1915.540 3116.300 1916.940 ;
        RECT 3067.300 1912.820 3110.300 1914.220 ;
        RECT 22.865 1910.100 114.865 1911.500 ;
        RECT 3062.500 1910.100 3104.300 1911.500 ;
        RECT 28.800 1907.380 110.100 1908.780 ;
        RECT 3057.800 1907.380 3098.300 1908.780 ;
        RECT 34.800 1904.660 81.300 1906.060 ;
        RECT 40.800 1901.940 86.100 1903.340 ;
        RECT 46.800 1899.220 90.850 1900.620 ;
        RECT 52.800 1896.500 95.800 1897.900 ;
        RECT 58.800 1893.780 100.600 1895.180 ;
        RECT 64.800 1891.060 105.300 1892.460 ;
        RECT 22.865 1844.820 114.865 1846.220 ;
        RECT 3048.235 1844.820 3140.235 1846.220 ;
        RECT 28.800 1842.100 110.100 1843.500 ;
        RECT 3053.000 1842.100 3134.300 1843.500 ;
        RECT 34.800 1839.380 81.300 1840.780 ;
        RECT 3081.800 1839.380 3128.300 1840.780 ;
        RECT 40.800 1836.660 86.100 1838.060 ;
        RECT 3077.000 1836.660 3122.300 1838.060 ;
        RECT 46.800 1833.940 90.850 1835.340 ;
        RECT 3072.250 1833.940 3116.300 1835.340 ;
        RECT 52.800 1831.220 95.800 1832.620 ;
        RECT 3067.300 1831.220 3110.300 1832.620 ;
        RECT 58.800 1828.500 100.600 1829.900 ;
        RECT 3062.500 1828.500 3104.300 1829.900 ;
        RECT 64.800 1825.780 105.300 1827.180 ;
        RECT 3057.800 1825.780 3098.300 1827.180 ;
        RECT 22.865 1779.540 114.865 1780.940 ;
        RECT 3048.235 1779.540 3140.235 1780.940 ;
        RECT 28.800 1776.820 110.100 1778.220 ;
        RECT 3053.000 1776.820 3134.300 1778.220 ;
        RECT 34.800 1774.100 81.300 1775.500 ;
        RECT 3081.800 1774.100 3128.300 1775.500 ;
        RECT 40.800 1771.380 86.100 1772.780 ;
        RECT 3077.000 1771.380 3122.300 1772.780 ;
        RECT 46.800 1768.660 90.850 1770.060 ;
        RECT 3072.250 1768.660 3116.300 1770.060 ;
        RECT 52.800 1765.940 95.800 1767.340 ;
        RECT 3067.300 1765.940 3110.300 1767.340 ;
        RECT 58.800 1763.220 100.600 1764.620 ;
        RECT 3062.500 1763.220 3104.300 1764.620 ;
        RECT 64.800 1760.500 105.300 1761.900 ;
        RECT 3057.800 1760.500 3098.300 1761.900 ;
        RECT 3048.235 1714.260 3140.235 1715.660 ;
        RECT 3053.000 1711.540 3134.300 1712.940 ;
        RECT 3081.800 1708.820 3128.300 1710.220 ;
        RECT 3077.000 1706.100 3122.300 1707.500 ;
        RECT 22.865 1703.380 114.865 1704.780 ;
        RECT 3072.250 1703.380 3116.300 1704.780 ;
        RECT 28.800 1700.660 110.100 1702.060 ;
        RECT 3067.300 1700.660 3110.300 1702.060 ;
        RECT 34.800 1697.940 81.300 1699.340 ;
        RECT 3062.500 1697.940 3104.300 1699.340 ;
        RECT 40.800 1695.220 86.100 1696.620 ;
        RECT 3057.800 1695.220 3098.300 1696.620 ;
        RECT 46.800 1692.500 90.850 1693.900 ;
        RECT 52.800 1689.780 95.800 1691.180 ;
        RECT 58.800 1687.060 100.600 1688.460 ;
        RECT 64.800 1684.340 105.300 1685.740 ;
        RECT 22.865 1648.980 114.865 1650.380 ;
        RECT 3048.235 1648.980 3140.235 1650.380 ;
        RECT 28.800 1646.260 110.100 1647.660 ;
        RECT 3053.000 1646.260 3134.300 1647.660 ;
        RECT 34.800 1643.540 81.300 1644.940 ;
        RECT 3081.800 1643.540 3128.300 1644.940 ;
        RECT 40.800 1640.820 86.100 1642.220 ;
        RECT 3077.000 1640.820 3122.300 1642.220 ;
        RECT 46.800 1638.100 90.850 1639.500 ;
        RECT 3072.250 1638.100 3116.300 1639.500 ;
        RECT 52.800 1635.380 95.800 1636.780 ;
        RECT 3067.300 1635.380 3110.300 1636.780 ;
        RECT 58.800 1632.660 100.600 1634.060 ;
        RECT 3062.500 1632.660 3104.300 1634.060 ;
        RECT 64.800 1629.940 105.300 1631.340 ;
        RECT 3057.800 1629.940 3098.300 1631.340 ;
        RECT 3048.235 1591.860 3140.235 1593.260 ;
        RECT 3053.000 1589.140 3134.300 1590.540 ;
        RECT 3081.800 1586.420 3128.300 1587.820 ;
        RECT 22.865 1583.700 114.865 1585.100 ;
        RECT 3077.000 1583.700 3122.300 1585.100 ;
        RECT 28.800 1580.980 110.100 1582.380 ;
        RECT 3072.250 1580.980 3116.300 1582.380 ;
        RECT 34.800 1578.260 81.300 1579.660 ;
        RECT 3067.300 1578.260 3110.300 1579.660 ;
        RECT 40.800 1575.540 86.100 1576.940 ;
        RECT 3062.500 1575.540 3104.300 1576.940 ;
        RECT 46.800 1572.820 90.850 1574.220 ;
        RECT 3057.800 1572.820 3098.300 1574.220 ;
        RECT 52.800 1570.100 95.800 1571.500 ;
        RECT 58.800 1567.380 100.600 1568.780 ;
        RECT 64.800 1564.660 105.300 1566.060 ;
        RECT 22.865 1529.300 114.865 1530.700 ;
        RECT 28.800 1526.580 110.100 1527.980 ;
        RECT 34.800 1523.860 81.300 1525.260 ;
        RECT 40.800 1521.140 86.100 1522.540 ;
        RECT 46.800 1518.420 90.850 1519.820 ;
        RECT 3048.235 1518.420 3140.235 1519.820 ;
        RECT 52.800 1515.700 95.800 1517.100 ;
        RECT 3053.000 1515.700 3134.300 1517.100 ;
        RECT 58.800 1512.980 100.600 1514.380 ;
        RECT 3081.800 1512.980 3128.300 1514.380 ;
        RECT 64.800 1510.260 105.300 1511.660 ;
        RECT 3077.000 1510.260 3122.300 1511.660 ;
        RECT 3072.250 1507.540 3116.300 1508.940 ;
        RECT 3067.300 1504.820 3110.300 1506.220 ;
        RECT 3062.500 1502.100 3104.300 1503.500 ;
        RECT 3057.800 1499.380 3098.300 1500.780 ;
        RECT 22.865 1453.140 114.865 1454.540 ;
        RECT 3048.235 1453.140 3140.235 1454.540 ;
        RECT 28.800 1450.420 110.100 1451.820 ;
        RECT 3053.000 1450.420 3134.300 1451.820 ;
        RECT 34.800 1447.700 81.300 1449.100 ;
        RECT 3081.800 1447.700 3128.300 1449.100 ;
        RECT 40.800 1444.980 86.100 1446.380 ;
        RECT 3077.000 1444.980 3122.300 1446.380 ;
        RECT 46.800 1442.260 90.850 1443.660 ;
        RECT 3072.250 1442.260 3116.300 1443.660 ;
        RECT 52.800 1439.540 95.800 1440.940 ;
        RECT 3067.300 1439.540 3110.300 1440.940 ;
        RECT 58.800 1436.820 100.600 1438.220 ;
        RECT 3062.500 1436.820 3104.300 1438.220 ;
        RECT 64.800 1434.100 105.300 1435.500 ;
        RECT 3057.800 1434.100 3098.300 1435.500 ;
        RECT 22.865 1387.860 114.865 1389.260 ;
        RECT 3048.235 1387.860 3140.235 1389.260 ;
        RECT 28.800 1385.140 110.100 1386.540 ;
        RECT 3053.000 1385.140 3134.300 1386.540 ;
        RECT 34.800 1382.420 81.300 1383.820 ;
        RECT 3081.800 1382.420 3128.300 1383.820 ;
        RECT 40.800 1379.700 86.100 1381.100 ;
        RECT 3077.000 1379.700 3122.300 1381.100 ;
        RECT 46.800 1376.980 90.850 1378.380 ;
        RECT 3072.250 1376.980 3116.300 1378.380 ;
        RECT 52.800 1374.260 95.800 1375.660 ;
        RECT 3067.300 1374.260 3110.300 1375.660 ;
        RECT 58.800 1371.540 100.600 1372.940 ;
        RECT 3062.500 1371.540 3104.300 1372.940 ;
        RECT 64.800 1368.820 105.300 1370.220 ;
        RECT 3057.800 1368.820 3098.300 1370.220 ;
        RECT 22.865 1333.460 114.865 1334.860 ;
        RECT 28.800 1330.740 110.100 1332.140 ;
        RECT 34.800 1328.020 81.300 1329.420 ;
        RECT 40.800 1325.300 86.100 1326.700 ;
        RECT 46.800 1322.580 90.850 1323.980 ;
        RECT 52.800 1319.860 95.800 1321.260 ;
        RECT 58.800 1317.140 100.600 1318.540 ;
        RECT 64.800 1314.420 105.300 1315.820 ;
        RECT 3048.235 1314.420 3140.235 1315.820 ;
        RECT 3053.000 1311.700 3134.300 1313.100 ;
        RECT 3081.800 1308.980 3128.300 1310.380 ;
        RECT 3077.000 1306.260 3122.300 1307.660 ;
        RECT 3072.250 1303.540 3116.300 1304.940 ;
        RECT 3067.300 1300.820 3110.300 1302.220 ;
        RECT 3062.500 1298.100 3104.300 1299.500 ;
        RECT 3057.800 1295.380 3098.300 1296.780 ;
        RECT 22.865 1257.300 114.865 1258.700 ;
        RECT 3048.235 1257.300 3140.235 1258.700 ;
        RECT 28.800 1254.580 110.100 1255.980 ;
        RECT 3053.000 1254.580 3134.300 1255.980 ;
        RECT 34.800 1251.860 81.300 1253.260 ;
        RECT 3081.800 1251.860 3128.300 1253.260 ;
        RECT 40.800 1249.140 86.100 1250.540 ;
        RECT 3077.000 1249.140 3122.300 1250.540 ;
        RECT 46.800 1246.420 90.850 1247.820 ;
        RECT 3072.250 1246.420 3116.300 1247.820 ;
        RECT 52.800 1243.700 95.800 1245.100 ;
        RECT 3067.300 1243.700 3110.300 1245.100 ;
        RECT 58.800 1240.980 100.600 1242.380 ;
        RECT 3062.500 1240.980 3104.300 1242.380 ;
        RECT 64.800 1238.260 105.300 1239.660 ;
        RECT 3057.800 1238.260 3098.300 1239.660 ;
        RECT 22.865 1192.020 114.865 1193.420 ;
        RECT 3048.235 1192.020 3140.235 1193.420 ;
        RECT 28.800 1189.300 110.100 1190.700 ;
        RECT 3053.000 1189.300 3134.300 1190.700 ;
        RECT 34.800 1186.580 81.300 1187.980 ;
        RECT 3081.800 1186.580 3128.300 1187.980 ;
        RECT 40.800 1183.860 86.100 1185.260 ;
        RECT 3077.000 1183.860 3122.300 1185.260 ;
        RECT 46.800 1181.140 90.850 1182.540 ;
        RECT 3072.250 1181.140 3116.300 1182.540 ;
        RECT 52.800 1178.420 95.800 1179.820 ;
        RECT 3067.300 1178.420 3110.300 1179.820 ;
        RECT 58.800 1175.700 100.600 1177.100 ;
        RECT 3062.500 1175.700 3104.300 1177.100 ;
        RECT 64.800 1172.980 105.300 1174.380 ;
        RECT 3057.800 1172.980 3098.300 1174.380 ;
        RECT 22.865 1126.740 114.865 1128.140 ;
        RECT 3048.235 1126.740 3140.235 1128.140 ;
        RECT 28.800 1124.020 110.100 1125.420 ;
        RECT 3053.000 1124.020 3134.300 1125.420 ;
        RECT 34.800 1121.300 81.300 1122.700 ;
        RECT 3081.800 1121.300 3128.300 1122.700 ;
        RECT 40.800 1118.580 86.100 1119.980 ;
        RECT 3077.000 1118.580 3122.300 1119.980 ;
        RECT 46.800 1115.860 90.850 1117.260 ;
        RECT 3072.250 1115.860 3116.300 1117.260 ;
        RECT 52.800 1113.140 95.800 1114.540 ;
        RECT 3067.300 1113.140 3110.300 1114.540 ;
        RECT 58.800 1110.420 100.600 1111.820 ;
        RECT 3062.500 1110.420 3104.300 1111.820 ;
        RECT 64.800 1107.700 105.300 1109.100 ;
        RECT 3057.800 1107.700 3098.300 1109.100 ;
        RECT 3048.235 1061.460 3140.235 1062.860 ;
        RECT 3053.000 1058.740 3134.300 1060.140 ;
        RECT 22.865 1056.020 114.865 1057.420 ;
        RECT 3081.800 1056.020 3128.300 1057.420 ;
        RECT 28.800 1053.300 110.100 1054.700 ;
        RECT 3077.000 1053.300 3122.300 1054.700 ;
        RECT 34.800 1050.580 81.300 1051.980 ;
        RECT 3072.250 1050.580 3116.300 1051.980 ;
        RECT 40.800 1047.860 86.100 1049.260 ;
        RECT 3067.300 1047.860 3110.300 1049.260 ;
        RECT 46.800 1045.140 90.850 1046.540 ;
        RECT 3062.500 1045.140 3104.300 1046.540 ;
        RECT 52.800 1042.420 95.800 1043.820 ;
        RECT 3057.800 1042.420 3098.300 1043.820 ;
        RECT 58.800 1039.700 100.600 1041.100 ;
        RECT 64.800 1036.980 105.300 1038.380 ;
        RECT 1040.720 135.270 1063.515 136.865 ;
        RECT 1135.120 134.500 1138.320 134.680 ;
        RECT 1117.920 133.265 1138.320 134.500 ;
        RECT 1135.120 133.095 1138.320 133.265 ;
        RECT 654.720 37.800 699.880 39.405 ;
        RECT 661.520 34.470 693.390 36.070 ;
      LAYER via3 ;
        RECT 3048.480 4554.080 3051.200 4555.200 ;
        RECT 3135.320 4554.080 3140.040 4555.200 ;
        RECT 3053.280 4551.360 3056.000 4552.480 ;
        RECT 3129.320 4551.360 3134.040 4552.480 ;
        RECT 3082.080 4548.640 3084.800 4549.760 ;
        RECT 3123.320 4548.640 3128.040 4549.760 ;
        RECT 3077.280 4545.920 3080.000 4547.040 ;
        RECT 3117.320 4545.920 3122.040 4547.040 ;
        RECT 3072.480 4543.200 3075.200 4544.320 ;
        RECT 3111.320 4543.200 3116.040 4544.320 ;
        RECT 3067.680 4540.480 3070.400 4541.600 ;
        RECT 3105.320 4540.480 3110.040 4541.600 ;
        RECT 3062.880 4537.760 3065.600 4538.880 ;
        RECT 3099.320 4537.760 3104.040 4538.880 ;
        RECT 3058.080 4535.040 3060.800 4536.160 ;
        RECT 3093.320 4535.040 3098.040 4536.160 ;
        RECT 23.060 4529.600 27.780 4530.720 ;
        RECT 111.900 4529.600 114.620 4530.720 ;
        RECT 29.060 4526.880 33.780 4528.000 ;
        RECT 107.100 4526.880 109.820 4528.000 ;
        RECT 35.060 4524.160 39.780 4525.280 ;
        RECT 78.300 4524.160 81.020 4525.280 ;
        RECT 41.060 4521.440 45.780 4522.560 ;
        RECT 83.100 4521.440 85.820 4522.560 ;
        RECT 47.060 4518.720 51.780 4519.840 ;
        RECT 87.900 4518.720 90.620 4519.840 ;
        RECT 53.060 4516.000 57.780 4517.120 ;
        RECT 92.700 4516.000 95.420 4517.120 ;
        RECT 59.060 4513.280 63.780 4514.400 ;
        RECT 97.500 4513.280 100.220 4514.400 ;
        RECT 65.060 4510.560 69.780 4511.680 ;
        RECT 102.300 4510.560 105.020 4511.680 ;
        RECT 3048.480 4480.640 3051.200 4481.760 ;
        RECT 3135.320 4480.640 3140.040 4481.760 ;
        RECT 3053.280 4477.920 3056.000 4479.040 ;
        RECT 3129.320 4477.920 3134.040 4479.040 ;
        RECT 3082.080 4475.200 3084.800 4476.320 ;
        RECT 3123.320 4475.200 3128.040 4476.320 ;
        RECT 3077.280 4472.480 3080.000 4473.600 ;
        RECT 3117.320 4472.480 3122.040 4473.600 ;
        RECT 3072.480 4469.760 3075.200 4470.880 ;
        RECT 3111.320 4469.760 3116.040 4470.880 ;
        RECT 3067.680 4467.040 3070.400 4468.160 ;
        RECT 3105.320 4467.040 3110.040 4468.160 ;
        RECT 3062.880 4464.320 3065.600 4465.440 ;
        RECT 3099.320 4464.320 3104.040 4465.440 ;
        RECT 3058.080 4461.600 3060.800 4462.720 ;
        RECT 3093.320 4461.600 3098.040 4462.720 ;
        RECT 23.060 4456.160 27.780 4457.280 ;
        RECT 111.900 4456.160 114.620 4457.280 ;
        RECT 29.060 4453.440 33.780 4454.560 ;
        RECT 107.100 4453.440 109.820 4454.560 ;
        RECT 35.060 4450.720 39.780 4451.840 ;
        RECT 78.300 4450.720 81.020 4451.840 ;
        RECT 41.060 4448.000 45.780 4449.120 ;
        RECT 83.100 4448.000 85.820 4449.120 ;
        RECT 47.060 4445.280 51.780 4446.400 ;
        RECT 87.900 4445.280 90.620 4446.400 ;
        RECT 53.060 4442.560 57.780 4443.680 ;
        RECT 92.700 4442.560 95.420 4443.680 ;
        RECT 59.060 4439.840 63.780 4440.960 ;
        RECT 97.500 4439.840 100.220 4440.960 ;
        RECT 65.060 4437.120 69.780 4438.240 ;
        RECT 102.300 4437.120 105.020 4438.240 ;
        RECT 3048.480 4423.520 3051.200 4424.640 ;
        RECT 3135.320 4423.520 3140.040 4424.640 ;
        RECT 3053.280 4420.800 3056.000 4421.920 ;
        RECT 3129.320 4420.800 3134.040 4421.920 ;
        RECT 3082.080 4418.080 3084.800 4419.200 ;
        RECT 3123.320 4418.080 3128.040 4419.200 ;
        RECT 3077.280 4415.360 3080.000 4416.480 ;
        RECT 3117.320 4415.360 3122.040 4416.480 ;
        RECT 3072.480 4412.640 3075.200 4413.760 ;
        RECT 3111.320 4412.640 3116.040 4413.760 ;
        RECT 3067.680 4409.920 3070.400 4411.040 ;
        RECT 3105.320 4409.920 3110.040 4411.040 ;
        RECT 3062.880 4407.200 3065.600 4408.320 ;
        RECT 3099.320 4407.200 3104.040 4408.320 ;
        RECT 3058.080 4404.480 3060.800 4405.600 ;
        RECT 3093.320 4404.480 3098.040 4405.600 ;
        RECT 23.060 4390.880 27.780 4392.000 ;
        RECT 111.900 4390.880 114.620 4392.000 ;
        RECT 29.060 4388.160 33.780 4389.280 ;
        RECT 107.100 4388.160 109.820 4389.280 ;
        RECT 35.060 4385.440 39.780 4386.560 ;
        RECT 78.300 4385.440 81.020 4386.560 ;
        RECT 41.060 4382.720 45.780 4383.840 ;
        RECT 83.100 4382.720 85.820 4383.840 ;
        RECT 47.060 4380.000 51.780 4381.120 ;
        RECT 87.900 4380.000 90.620 4381.120 ;
        RECT 53.060 4377.280 57.780 4378.400 ;
        RECT 92.700 4377.280 95.420 4378.400 ;
        RECT 59.060 4374.560 63.780 4375.680 ;
        RECT 97.500 4374.560 100.220 4375.680 ;
        RECT 65.060 4371.840 69.780 4372.960 ;
        RECT 102.300 4371.840 105.020 4372.960 ;
        RECT 3048.480 4358.240 3051.200 4359.360 ;
        RECT 3135.320 4358.240 3140.040 4359.360 ;
        RECT 3053.280 4355.520 3056.000 4356.640 ;
        RECT 3129.320 4355.520 3134.040 4356.640 ;
        RECT 3082.080 4352.800 3084.800 4353.920 ;
        RECT 3123.320 4352.800 3128.040 4353.920 ;
        RECT 3077.280 4350.080 3080.000 4351.200 ;
        RECT 3117.320 4350.080 3122.040 4351.200 ;
        RECT 3072.480 4347.360 3075.200 4348.480 ;
        RECT 3111.320 4347.360 3116.040 4348.480 ;
        RECT 3067.680 4344.640 3070.400 4345.760 ;
        RECT 3105.320 4344.640 3110.040 4345.760 ;
        RECT 3062.880 4341.920 3065.600 4343.040 ;
        RECT 3099.320 4341.920 3104.040 4343.040 ;
        RECT 3058.080 4339.200 3060.800 4340.320 ;
        RECT 3093.320 4339.200 3098.040 4340.320 ;
        RECT 23.060 4325.600 27.780 4326.720 ;
        RECT 111.900 4325.600 114.620 4326.720 ;
        RECT 29.060 4322.880 33.780 4324.000 ;
        RECT 107.100 4322.880 109.820 4324.000 ;
        RECT 35.060 4320.160 39.780 4321.280 ;
        RECT 78.300 4320.160 81.020 4321.280 ;
        RECT 41.060 4317.440 45.780 4318.560 ;
        RECT 83.100 4317.440 85.820 4318.560 ;
        RECT 47.060 4314.720 51.780 4315.840 ;
        RECT 87.900 4314.720 90.620 4315.840 ;
        RECT 53.060 4312.000 57.780 4313.120 ;
        RECT 92.700 4312.000 95.420 4313.120 ;
        RECT 59.060 4309.280 63.780 4310.400 ;
        RECT 97.500 4309.280 100.220 4310.400 ;
        RECT 65.060 4306.560 69.780 4307.680 ;
        RECT 102.300 4306.560 105.020 4307.680 ;
        RECT 3048.480 4292.960 3051.200 4294.080 ;
        RECT 3135.320 4292.960 3140.040 4294.080 ;
        RECT 3053.280 4290.240 3056.000 4291.360 ;
        RECT 3129.320 4290.240 3134.040 4291.360 ;
        RECT 3082.080 4287.520 3084.800 4288.640 ;
        RECT 3123.320 4287.520 3128.040 4288.640 ;
        RECT 3077.280 4284.800 3080.000 4285.920 ;
        RECT 3117.320 4284.800 3122.040 4285.920 ;
        RECT 3072.480 4282.080 3075.200 4283.200 ;
        RECT 3111.320 4282.080 3116.040 4283.200 ;
        RECT 3067.680 4279.360 3070.400 4280.480 ;
        RECT 3105.320 4279.360 3110.040 4280.480 ;
        RECT 3062.880 4276.640 3065.600 4277.760 ;
        RECT 3099.320 4276.640 3104.040 4277.760 ;
        RECT 3058.080 4273.920 3060.800 4275.040 ;
        RECT 3093.320 4273.920 3098.040 4275.040 ;
        RECT 23.060 4260.320 27.780 4261.440 ;
        RECT 111.900 4260.320 114.620 4261.440 ;
        RECT 29.060 4257.600 33.780 4258.720 ;
        RECT 107.100 4257.600 109.820 4258.720 ;
        RECT 35.060 4254.880 39.780 4256.000 ;
        RECT 78.300 4254.880 81.020 4256.000 ;
        RECT 41.060 4252.160 45.780 4253.280 ;
        RECT 83.100 4252.160 85.820 4253.280 ;
        RECT 47.060 4249.440 51.780 4250.560 ;
        RECT 87.900 4249.440 90.620 4250.560 ;
        RECT 53.060 4246.720 57.780 4247.840 ;
        RECT 92.700 4246.720 95.420 4247.840 ;
        RECT 59.060 4244.000 63.780 4245.120 ;
        RECT 97.500 4244.000 100.220 4245.120 ;
        RECT 65.060 4241.280 69.780 4242.400 ;
        RECT 102.300 4241.280 105.020 4242.400 ;
        RECT 3048.480 4227.680 3051.200 4228.800 ;
        RECT 3135.320 4227.680 3140.040 4228.800 ;
        RECT 3053.280 4224.960 3056.000 4226.080 ;
        RECT 3129.320 4224.960 3134.040 4226.080 ;
        RECT 3082.080 4222.240 3084.800 4223.360 ;
        RECT 3123.320 4222.240 3128.040 4223.360 ;
        RECT 3077.280 4219.520 3080.000 4220.640 ;
        RECT 3117.320 4219.520 3122.040 4220.640 ;
        RECT 3072.480 4216.800 3075.200 4217.920 ;
        RECT 3111.320 4216.800 3116.040 4217.920 ;
        RECT 3067.680 4214.080 3070.400 4215.200 ;
        RECT 3105.320 4214.080 3110.040 4215.200 ;
        RECT 3062.880 4211.360 3065.600 4212.480 ;
        RECT 3099.320 4211.360 3104.040 4212.480 ;
        RECT 3058.080 4208.640 3060.800 4209.760 ;
        RECT 3093.320 4208.640 3098.040 4209.760 ;
        RECT 23.060 4195.040 27.780 4196.160 ;
        RECT 111.900 4195.040 114.620 4196.160 ;
        RECT 29.060 4192.320 33.780 4193.440 ;
        RECT 107.100 4192.320 109.820 4193.440 ;
        RECT 35.060 4189.600 39.780 4190.720 ;
        RECT 78.300 4189.600 81.020 4190.720 ;
        RECT 41.060 4186.880 45.780 4188.000 ;
        RECT 83.100 4186.880 85.820 4188.000 ;
        RECT 47.060 4184.160 51.780 4185.280 ;
        RECT 87.900 4184.160 90.620 4185.280 ;
        RECT 53.060 4181.440 57.780 4182.560 ;
        RECT 92.700 4181.440 95.420 4182.560 ;
        RECT 59.060 4178.720 63.780 4179.840 ;
        RECT 97.500 4178.720 100.220 4179.840 ;
        RECT 65.060 4176.000 69.780 4177.120 ;
        RECT 102.300 4176.000 105.020 4177.120 ;
        RECT 3048.480 4162.400 3051.200 4163.520 ;
        RECT 3135.320 4162.400 3140.040 4163.520 ;
        RECT 3053.280 4159.680 3056.000 4160.800 ;
        RECT 3129.320 4159.680 3134.040 4160.800 ;
        RECT 3082.080 4156.960 3084.800 4158.080 ;
        RECT 3123.320 4156.960 3128.040 4158.080 ;
        RECT 3077.280 4154.240 3080.000 4155.360 ;
        RECT 3117.320 4154.240 3122.040 4155.360 ;
        RECT 3072.480 4151.520 3075.200 4152.640 ;
        RECT 3111.320 4151.520 3116.040 4152.640 ;
        RECT 3067.680 4148.800 3070.400 4149.920 ;
        RECT 3105.320 4148.800 3110.040 4149.920 ;
        RECT 3062.880 4146.080 3065.600 4147.200 ;
        RECT 3099.320 4146.080 3104.040 4147.200 ;
        RECT 3058.080 4143.360 3060.800 4144.480 ;
        RECT 3093.320 4143.360 3098.040 4144.480 ;
        RECT 23.060 4129.760 27.780 4130.880 ;
        RECT 111.900 4129.760 114.620 4130.880 ;
        RECT 29.060 4127.040 33.780 4128.160 ;
        RECT 107.100 4127.040 109.820 4128.160 ;
        RECT 35.060 4124.320 39.780 4125.440 ;
        RECT 78.300 4124.320 81.020 4125.440 ;
        RECT 41.060 4121.600 45.780 4122.720 ;
        RECT 83.100 4121.600 85.820 4122.720 ;
        RECT 47.060 4118.880 51.780 4120.000 ;
        RECT 87.900 4118.880 90.620 4120.000 ;
        RECT 53.060 4116.160 57.780 4117.280 ;
        RECT 92.700 4116.160 95.420 4117.280 ;
        RECT 59.060 4113.440 63.780 4114.560 ;
        RECT 97.500 4113.440 100.220 4114.560 ;
        RECT 65.060 4110.720 69.780 4111.840 ;
        RECT 102.300 4110.720 105.020 4111.840 ;
        RECT 3048.480 4097.120 3051.200 4098.240 ;
        RECT 3135.320 4097.120 3140.040 4098.240 ;
        RECT 3053.280 4094.400 3056.000 4095.520 ;
        RECT 3129.320 4094.400 3134.040 4095.520 ;
        RECT 3082.080 4091.680 3084.800 4092.800 ;
        RECT 3123.320 4091.680 3128.040 4092.800 ;
        RECT 3077.280 4088.960 3080.000 4090.080 ;
        RECT 3117.320 4088.960 3122.040 4090.080 ;
        RECT 3072.480 4086.240 3075.200 4087.360 ;
        RECT 3111.320 4086.240 3116.040 4087.360 ;
        RECT 3067.680 4083.520 3070.400 4084.640 ;
        RECT 3105.320 4083.520 3110.040 4084.640 ;
        RECT 3062.880 4080.800 3065.600 4081.920 ;
        RECT 3099.320 4080.800 3104.040 4081.920 ;
        RECT 3058.080 4078.080 3060.800 4079.200 ;
        RECT 3093.320 4078.080 3098.040 4079.200 ;
        RECT 23.060 4064.480 27.780 4065.600 ;
        RECT 111.900 4064.480 114.620 4065.600 ;
        RECT 29.060 4061.760 33.780 4062.880 ;
        RECT 107.100 4061.760 109.820 4062.880 ;
        RECT 35.060 4059.040 39.780 4060.160 ;
        RECT 78.300 4059.040 81.020 4060.160 ;
        RECT 41.060 4056.320 45.780 4057.440 ;
        RECT 83.100 4056.320 85.820 4057.440 ;
        RECT 47.060 4053.600 51.780 4054.720 ;
        RECT 87.900 4053.600 90.620 4054.720 ;
        RECT 53.060 4050.880 57.780 4052.000 ;
        RECT 92.700 4050.880 95.420 4052.000 ;
        RECT 59.060 4048.160 63.780 4049.280 ;
        RECT 97.500 4048.160 100.220 4049.280 ;
        RECT 65.060 4045.440 69.780 4046.560 ;
        RECT 102.300 4045.440 105.020 4046.560 ;
        RECT 3048.480 4031.840 3051.200 4032.960 ;
        RECT 3135.320 4031.840 3140.040 4032.960 ;
        RECT 3053.280 4029.120 3056.000 4030.240 ;
        RECT 3129.320 4029.120 3134.040 4030.240 ;
        RECT 3082.080 4026.400 3084.800 4027.520 ;
        RECT 3123.320 4026.400 3128.040 4027.520 ;
        RECT 3077.280 4023.680 3080.000 4024.800 ;
        RECT 3117.320 4023.680 3122.040 4024.800 ;
        RECT 3072.480 4020.960 3075.200 4022.080 ;
        RECT 3111.320 4020.960 3116.040 4022.080 ;
        RECT 3067.680 4018.240 3070.400 4019.360 ;
        RECT 3105.320 4018.240 3110.040 4019.360 ;
        RECT 3062.880 4015.520 3065.600 4016.640 ;
        RECT 3099.320 4015.520 3104.040 4016.640 ;
        RECT 3058.080 4012.800 3060.800 4013.920 ;
        RECT 3093.320 4012.800 3098.040 4013.920 ;
        RECT 23.060 3999.200 27.780 4000.320 ;
        RECT 111.900 3999.200 114.620 4000.320 ;
        RECT 29.060 3996.480 33.780 3997.600 ;
        RECT 107.100 3996.480 109.820 3997.600 ;
        RECT 35.060 3993.760 39.780 3994.880 ;
        RECT 78.300 3993.760 81.020 3994.880 ;
        RECT 41.060 3991.040 45.780 3992.160 ;
        RECT 83.100 3991.040 85.820 3992.160 ;
        RECT 47.060 3988.320 51.780 3989.440 ;
        RECT 87.900 3988.320 90.620 3989.440 ;
        RECT 53.060 3985.600 57.780 3986.720 ;
        RECT 92.700 3985.600 95.420 3986.720 ;
        RECT 59.060 3982.880 63.780 3984.000 ;
        RECT 97.500 3982.880 100.220 3984.000 ;
        RECT 65.060 3980.160 69.780 3981.280 ;
        RECT 102.300 3980.160 105.020 3981.280 ;
        RECT 3048.480 3966.560 3051.200 3967.680 ;
        RECT 3135.320 3966.560 3140.040 3967.680 ;
        RECT 3053.280 3963.840 3056.000 3964.960 ;
        RECT 3129.320 3963.840 3134.040 3964.960 ;
        RECT 3082.080 3961.120 3084.800 3962.240 ;
        RECT 3123.320 3961.120 3128.040 3962.240 ;
        RECT 3077.280 3958.400 3080.000 3959.520 ;
        RECT 3117.320 3958.400 3122.040 3959.520 ;
        RECT 3072.480 3955.680 3075.200 3956.800 ;
        RECT 3111.320 3955.680 3116.040 3956.800 ;
        RECT 3067.680 3952.960 3070.400 3954.080 ;
        RECT 3105.320 3952.960 3110.040 3954.080 ;
        RECT 3062.880 3950.240 3065.600 3951.360 ;
        RECT 3099.320 3950.240 3104.040 3951.360 ;
        RECT 3058.080 3947.520 3060.800 3948.640 ;
        RECT 3093.320 3947.520 3098.040 3948.640 ;
        RECT 23.060 3933.920 27.780 3935.040 ;
        RECT 111.900 3933.920 114.620 3935.040 ;
        RECT 29.060 3931.200 33.780 3932.320 ;
        RECT 107.100 3931.200 109.820 3932.320 ;
        RECT 35.060 3928.480 39.780 3929.600 ;
        RECT 78.300 3928.480 81.020 3929.600 ;
        RECT 41.060 3925.760 45.780 3926.880 ;
        RECT 83.100 3925.760 85.820 3926.880 ;
        RECT 47.060 3923.040 51.780 3924.160 ;
        RECT 87.900 3923.040 90.620 3924.160 ;
        RECT 53.060 3920.320 57.780 3921.440 ;
        RECT 92.700 3920.320 95.420 3921.440 ;
        RECT 59.060 3917.600 63.780 3918.720 ;
        RECT 97.500 3917.600 100.220 3918.720 ;
        RECT 65.060 3914.880 69.780 3916.000 ;
        RECT 102.300 3914.880 105.020 3916.000 ;
        RECT 3048.480 3901.280 3051.200 3902.400 ;
        RECT 3135.320 3901.280 3140.040 3902.400 ;
        RECT 3053.280 3898.560 3056.000 3899.680 ;
        RECT 3129.320 3898.560 3134.040 3899.680 ;
        RECT 3082.080 3895.840 3084.800 3896.960 ;
        RECT 3123.320 3895.840 3128.040 3896.960 ;
        RECT 3077.280 3893.120 3080.000 3894.240 ;
        RECT 3117.320 3893.120 3122.040 3894.240 ;
        RECT 3072.480 3890.400 3075.200 3891.520 ;
        RECT 3111.320 3890.400 3116.040 3891.520 ;
        RECT 3067.680 3887.680 3070.400 3888.800 ;
        RECT 3105.320 3887.680 3110.040 3888.800 ;
        RECT 3062.880 3884.960 3065.600 3886.080 ;
        RECT 3099.320 3884.960 3104.040 3886.080 ;
        RECT 3058.080 3882.240 3060.800 3883.360 ;
        RECT 3093.320 3882.240 3098.040 3883.360 ;
        RECT 23.060 3868.640 27.780 3869.760 ;
        RECT 111.900 3868.640 114.620 3869.760 ;
        RECT 29.060 3865.920 33.780 3867.040 ;
        RECT 107.100 3865.920 109.820 3867.040 ;
        RECT 35.060 3863.200 39.780 3864.320 ;
        RECT 78.300 3863.200 81.020 3864.320 ;
        RECT 41.060 3860.480 45.780 3861.600 ;
        RECT 83.100 3860.480 85.820 3861.600 ;
        RECT 47.060 3857.760 51.780 3858.880 ;
        RECT 87.900 3857.760 90.620 3858.880 ;
        RECT 53.060 3855.040 57.780 3856.160 ;
        RECT 92.700 3855.040 95.420 3856.160 ;
        RECT 59.060 3852.320 63.780 3853.440 ;
        RECT 97.500 3852.320 100.220 3853.440 ;
        RECT 65.060 3849.600 69.780 3850.720 ;
        RECT 102.300 3849.600 105.020 3850.720 ;
        RECT 3048.480 3836.000 3051.200 3837.120 ;
        RECT 3135.320 3836.000 3140.040 3837.120 ;
        RECT 3053.280 3833.280 3056.000 3834.400 ;
        RECT 3129.320 3833.280 3134.040 3834.400 ;
        RECT 3082.080 3830.560 3084.800 3831.680 ;
        RECT 3123.320 3830.560 3128.040 3831.680 ;
        RECT 3077.280 3827.840 3080.000 3828.960 ;
        RECT 3117.320 3827.840 3122.040 3828.960 ;
        RECT 3072.480 3825.120 3075.200 3826.240 ;
        RECT 3111.320 3825.120 3116.040 3826.240 ;
        RECT 3067.680 3822.400 3070.400 3823.520 ;
        RECT 3105.320 3822.400 3110.040 3823.520 ;
        RECT 3062.880 3819.680 3065.600 3820.800 ;
        RECT 3099.320 3819.680 3104.040 3820.800 ;
        RECT 3058.080 3816.960 3060.800 3818.080 ;
        RECT 3093.320 3816.960 3098.040 3818.080 ;
        RECT 23.060 3803.360 27.780 3804.480 ;
        RECT 111.900 3803.360 114.620 3804.480 ;
        RECT 29.060 3800.640 33.780 3801.760 ;
        RECT 107.100 3800.640 109.820 3801.760 ;
        RECT 35.060 3797.920 39.780 3799.040 ;
        RECT 78.300 3797.920 81.020 3799.040 ;
        RECT 41.060 3795.200 45.780 3796.320 ;
        RECT 83.100 3795.200 85.820 3796.320 ;
        RECT 47.060 3792.480 51.780 3793.600 ;
        RECT 87.900 3792.480 90.620 3793.600 ;
        RECT 53.060 3789.760 57.780 3790.880 ;
        RECT 92.700 3789.760 95.420 3790.880 ;
        RECT 59.060 3787.040 63.780 3788.160 ;
        RECT 97.500 3787.040 100.220 3788.160 ;
        RECT 65.060 3784.320 69.780 3785.440 ;
        RECT 102.300 3784.320 105.020 3785.440 ;
        RECT 3048.480 3770.720 3051.200 3771.840 ;
        RECT 3135.320 3770.720 3140.040 3771.840 ;
        RECT 3053.280 3768.000 3056.000 3769.120 ;
        RECT 3129.320 3768.000 3134.040 3769.120 ;
        RECT 3082.080 3765.280 3084.800 3766.400 ;
        RECT 3123.320 3765.280 3128.040 3766.400 ;
        RECT 3077.280 3762.560 3080.000 3763.680 ;
        RECT 3117.320 3762.560 3122.040 3763.680 ;
        RECT 3072.480 3759.840 3075.200 3760.960 ;
        RECT 3111.320 3759.840 3116.040 3760.960 ;
        RECT 3067.680 3757.120 3070.400 3758.240 ;
        RECT 3105.320 3757.120 3110.040 3758.240 ;
        RECT 3062.880 3754.400 3065.600 3755.520 ;
        RECT 3099.320 3754.400 3104.040 3755.520 ;
        RECT 3058.080 3751.680 3060.800 3752.800 ;
        RECT 3093.320 3751.680 3098.040 3752.800 ;
        RECT 23.060 3738.080 27.780 3739.200 ;
        RECT 111.900 3738.080 114.620 3739.200 ;
        RECT 29.060 3735.360 33.780 3736.480 ;
        RECT 107.100 3735.360 109.820 3736.480 ;
        RECT 35.060 3732.640 39.780 3733.760 ;
        RECT 78.300 3732.640 81.020 3733.760 ;
        RECT 41.060 3729.920 45.780 3731.040 ;
        RECT 83.100 3729.920 85.820 3731.040 ;
        RECT 47.060 3727.200 51.780 3728.320 ;
        RECT 87.900 3727.200 90.620 3728.320 ;
        RECT 53.060 3724.480 57.780 3725.600 ;
        RECT 92.700 3724.480 95.420 3725.600 ;
        RECT 59.060 3721.760 63.780 3722.880 ;
        RECT 97.500 3721.760 100.220 3722.880 ;
        RECT 65.060 3719.040 69.780 3720.160 ;
        RECT 102.300 3719.040 105.020 3720.160 ;
        RECT 3048.480 3705.440 3051.200 3706.560 ;
        RECT 3135.320 3705.440 3140.040 3706.560 ;
        RECT 3053.280 3702.720 3056.000 3703.840 ;
        RECT 3129.320 3702.720 3134.040 3703.840 ;
        RECT 3082.080 3700.000 3084.800 3701.120 ;
        RECT 3123.320 3700.000 3128.040 3701.120 ;
        RECT 3077.280 3697.280 3080.000 3698.400 ;
        RECT 3117.320 3697.280 3122.040 3698.400 ;
        RECT 3072.480 3694.560 3075.200 3695.680 ;
        RECT 3111.320 3694.560 3116.040 3695.680 ;
        RECT 3067.680 3691.840 3070.400 3692.960 ;
        RECT 3105.320 3691.840 3110.040 3692.960 ;
        RECT 3062.880 3689.120 3065.600 3690.240 ;
        RECT 3099.320 3689.120 3104.040 3690.240 ;
        RECT 3058.080 3686.400 3060.800 3687.520 ;
        RECT 3093.320 3686.400 3098.040 3687.520 ;
        RECT 23.060 3680.960 27.780 3682.080 ;
        RECT 111.900 3680.960 114.620 3682.080 ;
        RECT 29.060 3678.240 33.780 3679.360 ;
        RECT 107.100 3678.240 109.820 3679.360 ;
        RECT 35.060 3675.520 39.780 3676.640 ;
        RECT 78.300 3675.520 81.020 3676.640 ;
        RECT 41.060 3672.800 45.780 3673.920 ;
        RECT 83.100 3672.800 85.820 3673.920 ;
        RECT 47.060 3670.080 51.780 3671.200 ;
        RECT 87.900 3670.080 90.620 3671.200 ;
        RECT 53.060 3667.360 57.780 3668.480 ;
        RECT 92.700 3667.360 95.420 3668.480 ;
        RECT 59.060 3664.640 63.780 3665.760 ;
        RECT 97.500 3664.640 100.220 3665.760 ;
        RECT 65.060 3661.920 69.780 3663.040 ;
        RECT 102.300 3661.920 105.020 3663.040 ;
        RECT 3048.480 3640.160 3051.200 3641.280 ;
        RECT 3135.320 3640.160 3140.040 3641.280 ;
        RECT 3053.280 3637.440 3056.000 3638.560 ;
        RECT 3129.320 3637.440 3134.040 3638.560 ;
        RECT 3082.080 3634.720 3084.800 3635.840 ;
        RECT 3123.320 3634.720 3128.040 3635.840 ;
        RECT 3077.280 3632.000 3080.000 3633.120 ;
        RECT 3117.320 3632.000 3122.040 3633.120 ;
        RECT 3072.480 3629.280 3075.200 3630.400 ;
        RECT 3111.320 3629.280 3116.040 3630.400 ;
        RECT 3067.680 3626.560 3070.400 3627.680 ;
        RECT 3105.320 3626.560 3110.040 3627.680 ;
        RECT 3062.880 3623.840 3065.600 3624.960 ;
        RECT 3099.320 3623.840 3104.040 3624.960 ;
        RECT 3058.080 3621.120 3060.800 3622.240 ;
        RECT 3093.320 3621.120 3098.040 3622.240 ;
        RECT 23.060 3607.520 27.780 3608.640 ;
        RECT 111.900 3607.520 114.620 3608.640 ;
        RECT 29.060 3604.800 33.780 3605.920 ;
        RECT 107.100 3604.800 109.820 3605.920 ;
        RECT 35.060 3602.080 39.780 3603.200 ;
        RECT 78.300 3602.080 81.020 3603.200 ;
        RECT 41.060 3599.360 45.780 3600.480 ;
        RECT 83.100 3599.360 85.820 3600.480 ;
        RECT 47.060 3596.640 51.780 3597.760 ;
        RECT 87.900 3596.640 90.620 3597.760 ;
        RECT 53.060 3593.920 57.780 3595.040 ;
        RECT 92.700 3593.920 95.420 3595.040 ;
        RECT 59.060 3591.200 63.780 3592.320 ;
        RECT 97.500 3591.200 100.220 3592.320 ;
        RECT 65.060 3588.480 69.780 3589.600 ;
        RECT 102.300 3588.480 105.020 3589.600 ;
        RECT 3048.480 3566.720 3051.200 3567.840 ;
        RECT 3135.320 3566.720 3140.040 3567.840 ;
        RECT 3053.280 3564.000 3056.000 3565.120 ;
        RECT 3129.320 3564.000 3134.040 3565.120 ;
        RECT 3082.080 3561.280 3084.800 3562.400 ;
        RECT 3123.320 3561.280 3128.040 3562.400 ;
        RECT 3077.280 3558.560 3080.000 3559.680 ;
        RECT 3117.320 3558.560 3122.040 3559.680 ;
        RECT 3072.480 3555.840 3075.200 3556.960 ;
        RECT 3111.320 3555.840 3116.040 3556.960 ;
        RECT 3067.680 3553.120 3070.400 3554.240 ;
        RECT 3105.320 3553.120 3110.040 3554.240 ;
        RECT 3062.880 3550.400 3065.600 3551.520 ;
        RECT 3099.320 3550.400 3104.040 3551.520 ;
        RECT 3058.080 3547.680 3060.800 3548.800 ;
        RECT 3093.320 3547.680 3098.040 3548.800 ;
        RECT 23.060 3542.240 27.780 3543.360 ;
        RECT 111.900 3542.240 114.620 3543.360 ;
        RECT 29.060 3539.520 33.780 3540.640 ;
        RECT 107.100 3539.520 109.820 3540.640 ;
        RECT 35.060 3536.800 39.780 3537.920 ;
        RECT 78.300 3536.800 81.020 3537.920 ;
        RECT 41.060 3534.080 45.780 3535.200 ;
        RECT 83.100 3534.080 85.820 3535.200 ;
        RECT 47.060 3531.360 51.780 3532.480 ;
        RECT 87.900 3531.360 90.620 3532.480 ;
        RECT 53.060 3528.640 57.780 3529.760 ;
        RECT 92.700 3528.640 95.420 3529.760 ;
        RECT 59.060 3525.920 63.780 3527.040 ;
        RECT 97.500 3525.920 100.220 3527.040 ;
        RECT 65.060 3523.200 69.780 3524.320 ;
        RECT 102.300 3523.200 105.020 3524.320 ;
        RECT 3048.480 3509.600 3051.200 3510.720 ;
        RECT 3135.320 3509.600 3140.040 3510.720 ;
        RECT 3053.280 3506.880 3056.000 3508.000 ;
        RECT 3129.320 3506.880 3134.040 3508.000 ;
        RECT 3082.080 3504.160 3084.800 3505.280 ;
        RECT 3123.320 3504.160 3128.040 3505.280 ;
        RECT 3077.280 3501.440 3080.000 3502.560 ;
        RECT 3117.320 3501.440 3122.040 3502.560 ;
        RECT 3072.480 3498.720 3075.200 3499.840 ;
        RECT 3111.320 3498.720 3116.040 3499.840 ;
        RECT 3067.680 3496.000 3070.400 3497.120 ;
        RECT 3105.320 3496.000 3110.040 3497.120 ;
        RECT 3062.880 3493.280 3065.600 3494.400 ;
        RECT 3099.320 3493.280 3104.040 3494.400 ;
        RECT 3058.080 3490.560 3060.800 3491.680 ;
        RECT 3093.320 3490.560 3098.040 3491.680 ;
        RECT 23.060 3460.640 27.780 3461.760 ;
        RECT 111.900 3460.640 114.620 3461.760 ;
        RECT 29.060 3457.920 33.780 3459.040 ;
        RECT 107.100 3457.920 109.820 3459.040 ;
        RECT 35.060 3455.200 39.780 3456.320 ;
        RECT 78.300 3455.200 81.020 3456.320 ;
        RECT 41.060 3452.480 45.780 3453.600 ;
        RECT 83.100 3452.480 85.820 3453.600 ;
        RECT 47.060 3449.760 51.780 3450.880 ;
        RECT 87.900 3449.760 90.620 3450.880 ;
        RECT 53.060 3447.040 57.780 3448.160 ;
        RECT 92.700 3447.040 95.420 3448.160 ;
        RECT 59.060 3444.320 63.780 3445.440 ;
        RECT 97.500 3444.320 100.220 3445.440 ;
        RECT 3048.480 3444.320 3051.200 3445.440 ;
        RECT 3135.320 3444.320 3140.040 3445.440 ;
        RECT 65.060 3441.600 69.780 3442.720 ;
        RECT 102.300 3441.600 105.020 3442.720 ;
        RECT 3053.280 3441.600 3056.000 3442.720 ;
        RECT 3129.320 3441.600 3134.040 3442.720 ;
        RECT 3082.080 3438.880 3084.800 3440.000 ;
        RECT 3123.320 3438.880 3128.040 3440.000 ;
        RECT 3077.280 3436.160 3080.000 3437.280 ;
        RECT 3117.320 3436.160 3122.040 3437.280 ;
        RECT 3072.480 3433.440 3075.200 3434.560 ;
        RECT 3111.320 3433.440 3116.040 3434.560 ;
        RECT 3067.680 3430.720 3070.400 3431.840 ;
        RECT 3105.320 3430.720 3110.040 3431.840 ;
        RECT 3062.880 3428.000 3065.600 3429.120 ;
        RECT 3099.320 3428.000 3104.040 3429.120 ;
        RECT 3058.080 3425.280 3060.800 3426.400 ;
        RECT 3093.320 3425.280 3098.040 3426.400 ;
        RECT 23.060 3411.680 27.780 3412.800 ;
        RECT 111.900 3411.680 114.620 3412.800 ;
        RECT 29.060 3408.960 33.780 3410.080 ;
        RECT 107.100 3408.960 109.820 3410.080 ;
        RECT 35.060 3406.240 39.780 3407.360 ;
        RECT 78.300 3406.240 81.020 3407.360 ;
        RECT 41.060 3403.520 45.780 3404.640 ;
        RECT 83.100 3403.520 85.820 3404.640 ;
        RECT 47.060 3400.800 51.780 3401.920 ;
        RECT 87.900 3400.800 90.620 3401.920 ;
        RECT 53.060 3398.080 57.780 3399.200 ;
        RECT 92.700 3398.080 95.420 3399.200 ;
        RECT 59.060 3395.360 63.780 3396.480 ;
        RECT 97.500 3395.360 100.220 3396.480 ;
        RECT 65.060 3392.640 69.780 3393.760 ;
        RECT 102.300 3392.640 105.020 3393.760 ;
        RECT 3048.480 3379.040 3051.200 3380.160 ;
        RECT 3135.320 3379.040 3140.040 3380.160 ;
        RECT 3053.280 3376.320 3056.000 3377.440 ;
        RECT 3129.320 3376.320 3134.040 3377.440 ;
        RECT 3082.080 3373.600 3084.800 3374.720 ;
        RECT 3123.320 3373.600 3128.040 3374.720 ;
        RECT 3077.280 3370.880 3080.000 3372.000 ;
        RECT 3117.320 3370.880 3122.040 3372.000 ;
        RECT 3072.480 3368.160 3075.200 3369.280 ;
        RECT 3111.320 3368.160 3116.040 3369.280 ;
        RECT 3067.680 3365.440 3070.400 3366.560 ;
        RECT 3105.320 3365.440 3110.040 3366.560 ;
        RECT 3062.880 3362.720 3065.600 3363.840 ;
        RECT 3099.320 3362.720 3104.040 3363.840 ;
        RECT 3058.080 3360.000 3060.800 3361.120 ;
        RECT 3093.320 3360.000 3098.040 3361.120 ;
        RECT 23.060 3346.400 27.780 3347.520 ;
        RECT 111.900 3346.400 114.620 3347.520 ;
        RECT 29.060 3343.680 33.780 3344.800 ;
        RECT 107.100 3343.680 109.820 3344.800 ;
        RECT 35.060 3340.960 39.780 3342.080 ;
        RECT 78.300 3340.960 81.020 3342.080 ;
        RECT 41.060 3338.240 45.780 3339.360 ;
        RECT 83.100 3338.240 85.820 3339.360 ;
        RECT 47.060 3335.520 51.780 3336.640 ;
        RECT 87.900 3335.520 90.620 3336.640 ;
        RECT 53.060 3332.800 57.780 3333.920 ;
        RECT 92.700 3332.800 95.420 3333.920 ;
        RECT 59.060 3330.080 63.780 3331.200 ;
        RECT 97.500 3330.080 100.220 3331.200 ;
        RECT 65.060 3327.360 69.780 3328.480 ;
        RECT 102.300 3327.360 105.020 3328.480 ;
        RECT 3048.480 3313.760 3051.200 3314.880 ;
        RECT 3135.320 3313.760 3140.040 3314.880 ;
        RECT 3053.280 3311.040 3056.000 3312.160 ;
        RECT 3129.320 3311.040 3134.040 3312.160 ;
        RECT 3082.080 3308.320 3084.800 3309.440 ;
        RECT 3123.320 3308.320 3128.040 3309.440 ;
        RECT 3077.280 3305.600 3080.000 3306.720 ;
        RECT 3117.320 3305.600 3122.040 3306.720 ;
        RECT 3072.480 3302.880 3075.200 3304.000 ;
        RECT 3111.320 3302.880 3116.040 3304.000 ;
        RECT 3067.680 3300.160 3070.400 3301.280 ;
        RECT 3105.320 3300.160 3110.040 3301.280 ;
        RECT 3062.880 3297.440 3065.600 3298.560 ;
        RECT 3099.320 3297.440 3104.040 3298.560 ;
        RECT 3058.080 3294.720 3060.800 3295.840 ;
        RECT 3093.320 3294.720 3098.040 3295.840 ;
        RECT 23.060 3281.120 27.780 3282.240 ;
        RECT 111.900 3281.120 114.620 3282.240 ;
        RECT 29.060 3278.400 33.780 3279.520 ;
        RECT 107.100 3278.400 109.820 3279.520 ;
        RECT 35.060 3275.680 39.780 3276.800 ;
        RECT 78.300 3275.680 81.020 3276.800 ;
        RECT 41.060 3272.960 45.780 3274.080 ;
        RECT 83.100 3272.960 85.820 3274.080 ;
        RECT 47.060 3270.240 51.780 3271.360 ;
        RECT 87.900 3270.240 90.620 3271.360 ;
        RECT 53.060 3267.520 57.780 3268.640 ;
        RECT 92.700 3267.520 95.420 3268.640 ;
        RECT 59.060 3264.800 63.780 3265.920 ;
        RECT 97.500 3264.800 100.220 3265.920 ;
        RECT 65.060 3262.080 69.780 3263.200 ;
        RECT 102.300 3262.080 105.020 3263.200 ;
        RECT 3048.480 3248.480 3051.200 3249.600 ;
        RECT 3135.320 3248.480 3140.040 3249.600 ;
        RECT 3053.280 3245.760 3056.000 3246.880 ;
        RECT 3129.320 3245.760 3134.040 3246.880 ;
        RECT 3082.080 3243.040 3084.800 3244.160 ;
        RECT 3123.320 3243.040 3128.040 3244.160 ;
        RECT 3077.280 3240.320 3080.000 3241.440 ;
        RECT 3117.320 3240.320 3122.040 3241.440 ;
        RECT 3072.480 3237.600 3075.200 3238.720 ;
        RECT 3111.320 3237.600 3116.040 3238.720 ;
        RECT 3067.680 3234.880 3070.400 3236.000 ;
        RECT 3105.320 3234.880 3110.040 3236.000 ;
        RECT 3062.880 3232.160 3065.600 3233.280 ;
        RECT 3099.320 3232.160 3104.040 3233.280 ;
        RECT 3058.080 3229.440 3060.800 3230.560 ;
        RECT 3093.320 3229.440 3098.040 3230.560 ;
        RECT 23.060 3207.680 27.780 3208.800 ;
        RECT 111.900 3207.680 114.620 3208.800 ;
        RECT 29.060 3204.960 33.780 3206.080 ;
        RECT 107.100 3204.960 109.820 3206.080 ;
        RECT 35.060 3202.240 39.780 3203.360 ;
        RECT 78.300 3202.240 81.020 3203.360 ;
        RECT 41.060 3199.520 45.780 3200.640 ;
        RECT 83.100 3199.520 85.820 3200.640 ;
        RECT 47.060 3196.800 51.780 3197.920 ;
        RECT 87.900 3196.800 90.620 3197.920 ;
        RECT 53.060 3194.080 57.780 3195.200 ;
        RECT 92.700 3194.080 95.420 3195.200 ;
        RECT 59.060 3191.360 63.780 3192.480 ;
        RECT 97.500 3191.360 100.220 3192.480 ;
        RECT 65.060 3188.640 69.780 3189.760 ;
        RECT 102.300 3188.640 105.020 3189.760 ;
        RECT 3048.480 3183.200 3051.200 3184.320 ;
        RECT 3135.320 3183.200 3140.040 3184.320 ;
        RECT 3053.280 3180.480 3056.000 3181.600 ;
        RECT 3129.320 3180.480 3134.040 3181.600 ;
        RECT 3082.080 3177.760 3084.800 3178.880 ;
        RECT 3123.320 3177.760 3128.040 3178.880 ;
        RECT 3077.280 3175.040 3080.000 3176.160 ;
        RECT 3117.320 3175.040 3122.040 3176.160 ;
        RECT 3072.480 3172.320 3075.200 3173.440 ;
        RECT 3111.320 3172.320 3116.040 3173.440 ;
        RECT 3067.680 3169.600 3070.400 3170.720 ;
        RECT 3105.320 3169.600 3110.040 3170.720 ;
        RECT 3062.880 3166.880 3065.600 3168.000 ;
        RECT 3099.320 3166.880 3104.040 3168.000 ;
        RECT 3058.080 3164.160 3060.800 3165.280 ;
        RECT 3093.320 3164.160 3098.040 3165.280 ;
        RECT 23.060 3150.560 27.780 3151.680 ;
        RECT 111.900 3150.560 114.620 3151.680 ;
        RECT 29.060 3147.840 33.780 3148.960 ;
        RECT 107.100 3147.840 109.820 3148.960 ;
        RECT 35.060 3145.120 39.780 3146.240 ;
        RECT 78.300 3145.120 81.020 3146.240 ;
        RECT 41.060 3142.400 45.780 3143.520 ;
        RECT 83.100 3142.400 85.820 3143.520 ;
        RECT 47.060 3139.680 51.780 3140.800 ;
        RECT 87.900 3139.680 90.620 3140.800 ;
        RECT 53.060 3136.960 57.780 3138.080 ;
        RECT 92.700 3136.960 95.420 3138.080 ;
        RECT 59.060 3134.240 63.780 3135.360 ;
        RECT 97.500 3134.240 100.220 3135.360 ;
        RECT 65.060 3131.520 69.780 3132.640 ;
        RECT 102.300 3131.520 105.020 3132.640 ;
        RECT 3048.480 3117.920 3051.200 3119.040 ;
        RECT 3135.320 3117.920 3140.040 3119.040 ;
        RECT 3053.280 3115.200 3056.000 3116.320 ;
        RECT 3129.320 3115.200 3134.040 3116.320 ;
        RECT 3082.080 3112.480 3084.800 3113.600 ;
        RECT 3123.320 3112.480 3128.040 3113.600 ;
        RECT 3077.280 3109.760 3080.000 3110.880 ;
        RECT 3117.320 3109.760 3122.040 3110.880 ;
        RECT 3072.480 3107.040 3075.200 3108.160 ;
        RECT 3111.320 3107.040 3116.040 3108.160 ;
        RECT 3067.680 3104.320 3070.400 3105.440 ;
        RECT 3105.320 3104.320 3110.040 3105.440 ;
        RECT 3062.880 3101.600 3065.600 3102.720 ;
        RECT 3099.320 3101.600 3104.040 3102.720 ;
        RECT 3058.080 3098.880 3060.800 3100.000 ;
        RECT 3093.320 3098.880 3098.040 3100.000 ;
        RECT 23.060 3085.280 27.780 3086.400 ;
        RECT 111.900 3085.280 114.620 3086.400 ;
        RECT 29.060 3082.560 33.780 3083.680 ;
        RECT 107.100 3082.560 109.820 3083.680 ;
        RECT 35.060 3079.840 39.780 3080.960 ;
        RECT 78.300 3079.840 81.020 3080.960 ;
        RECT 41.060 3077.120 45.780 3078.240 ;
        RECT 83.100 3077.120 85.820 3078.240 ;
        RECT 47.060 3074.400 51.780 3075.520 ;
        RECT 87.900 3074.400 90.620 3075.520 ;
        RECT 53.060 3071.680 57.780 3072.800 ;
        RECT 92.700 3071.680 95.420 3072.800 ;
        RECT 59.060 3068.960 63.780 3070.080 ;
        RECT 97.500 3068.960 100.220 3070.080 ;
        RECT 65.060 3066.240 69.780 3067.360 ;
        RECT 102.300 3066.240 105.020 3067.360 ;
        RECT 3048.480 3052.640 3051.200 3053.760 ;
        RECT 3135.320 3052.640 3140.040 3053.760 ;
        RECT 3053.280 3049.920 3056.000 3051.040 ;
        RECT 3129.320 3049.920 3134.040 3051.040 ;
        RECT 3082.080 3047.200 3084.800 3048.320 ;
        RECT 3123.320 3047.200 3128.040 3048.320 ;
        RECT 3077.280 3044.480 3080.000 3045.600 ;
        RECT 3117.320 3044.480 3122.040 3045.600 ;
        RECT 3072.480 3041.760 3075.200 3042.880 ;
        RECT 3111.320 3041.760 3116.040 3042.880 ;
        RECT 3067.680 3039.040 3070.400 3040.160 ;
        RECT 3105.320 3039.040 3110.040 3040.160 ;
        RECT 3062.880 3036.320 3065.600 3037.440 ;
        RECT 3099.320 3036.320 3104.040 3037.440 ;
        RECT 3058.080 3033.600 3060.800 3034.720 ;
        RECT 3093.320 3033.600 3098.040 3034.720 ;
        RECT 23.060 3030.880 27.780 3032.000 ;
        RECT 111.900 3030.880 114.620 3032.000 ;
        RECT 29.060 3028.160 33.780 3029.280 ;
        RECT 107.100 3028.160 109.820 3029.280 ;
        RECT 35.060 3025.440 39.780 3026.560 ;
        RECT 78.300 3025.440 81.020 3026.560 ;
        RECT 41.060 3022.720 45.780 3023.840 ;
        RECT 83.100 3022.720 85.820 3023.840 ;
        RECT 47.060 3020.000 51.780 3021.120 ;
        RECT 87.900 3020.000 90.620 3021.120 ;
        RECT 53.060 3017.280 57.780 3018.400 ;
        RECT 92.700 3017.280 95.420 3018.400 ;
        RECT 59.060 3014.560 63.780 3015.680 ;
        RECT 97.500 3014.560 100.220 3015.680 ;
        RECT 65.060 3011.840 69.780 3012.960 ;
        RECT 102.300 3011.840 105.020 3012.960 ;
        RECT 3048.480 2987.360 3051.200 2988.480 ;
        RECT 3135.320 2987.360 3140.040 2988.480 ;
        RECT 3053.280 2984.640 3056.000 2985.760 ;
        RECT 3129.320 2984.640 3134.040 2985.760 ;
        RECT 3082.080 2981.920 3084.800 2983.040 ;
        RECT 3123.320 2981.920 3128.040 2983.040 ;
        RECT 3077.280 2979.200 3080.000 2980.320 ;
        RECT 3117.320 2979.200 3122.040 2980.320 ;
        RECT 3072.480 2976.480 3075.200 2977.600 ;
        RECT 3111.320 2976.480 3116.040 2977.600 ;
        RECT 3067.680 2973.760 3070.400 2974.880 ;
        RECT 3105.320 2973.760 3110.040 2974.880 ;
        RECT 3062.880 2971.040 3065.600 2972.160 ;
        RECT 3099.320 2971.040 3104.040 2972.160 ;
        RECT 3058.080 2968.320 3060.800 2969.440 ;
        RECT 3093.320 2968.320 3098.040 2969.440 ;
        RECT 23.060 2954.720 27.780 2955.840 ;
        RECT 111.900 2954.720 114.620 2955.840 ;
        RECT 29.060 2952.000 33.780 2953.120 ;
        RECT 107.100 2952.000 109.820 2953.120 ;
        RECT 35.060 2949.280 39.780 2950.400 ;
        RECT 78.300 2949.280 81.020 2950.400 ;
        RECT 41.060 2946.560 45.780 2947.680 ;
        RECT 83.100 2946.560 85.820 2947.680 ;
        RECT 47.060 2943.840 51.780 2944.960 ;
        RECT 87.900 2943.840 90.620 2944.960 ;
        RECT 53.060 2941.120 57.780 2942.240 ;
        RECT 92.700 2941.120 95.420 2942.240 ;
        RECT 59.060 2938.400 63.780 2939.520 ;
        RECT 97.500 2938.400 100.220 2939.520 ;
        RECT 65.060 2935.680 69.780 2936.800 ;
        RECT 102.300 2935.680 105.020 2936.800 ;
        RECT 3048.480 2922.080 3051.200 2923.200 ;
        RECT 3135.320 2922.080 3140.040 2923.200 ;
        RECT 3053.280 2919.360 3056.000 2920.480 ;
        RECT 3129.320 2919.360 3134.040 2920.480 ;
        RECT 3082.080 2916.640 3084.800 2917.760 ;
        RECT 3123.320 2916.640 3128.040 2917.760 ;
        RECT 3077.280 2913.920 3080.000 2915.040 ;
        RECT 3117.320 2913.920 3122.040 2915.040 ;
        RECT 3072.480 2911.200 3075.200 2912.320 ;
        RECT 3111.320 2911.200 3116.040 2912.320 ;
        RECT 3067.680 2908.480 3070.400 2909.600 ;
        RECT 3105.320 2908.480 3110.040 2909.600 ;
        RECT 3062.880 2905.760 3065.600 2906.880 ;
        RECT 3099.320 2905.760 3104.040 2906.880 ;
        RECT 3058.080 2903.040 3060.800 2904.160 ;
        RECT 3093.320 2903.040 3098.040 2904.160 ;
        RECT 23.060 2889.440 27.780 2890.560 ;
        RECT 111.900 2889.440 114.620 2890.560 ;
        RECT 29.060 2886.720 33.780 2887.840 ;
        RECT 107.100 2886.720 109.820 2887.840 ;
        RECT 35.060 2884.000 39.780 2885.120 ;
        RECT 78.300 2884.000 81.020 2885.120 ;
        RECT 41.060 2881.280 45.780 2882.400 ;
        RECT 83.100 2881.280 85.820 2882.400 ;
        RECT 47.060 2878.560 51.780 2879.680 ;
        RECT 87.900 2878.560 90.620 2879.680 ;
        RECT 53.060 2875.840 57.780 2876.960 ;
        RECT 92.700 2875.840 95.420 2876.960 ;
        RECT 59.060 2873.120 63.780 2874.240 ;
        RECT 97.500 2873.120 100.220 2874.240 ;
        RECT 65.060 2870.400 69.780 2871.520 ;
        RECT 102.300 2870.400 105.020 2871.520 ;
        RECT 3048.480 2856.800 3051.200 2857.920 ;
        RECT 3135.320 2856.800 3140.040 2857.920 ;
        RECT 3053.280 2854.080 3056.000 2855.200 ;
        RECT 3129.320 2854.080 3134.040 2855.200 ;
        RECT 3082.080 2851.360 3084.800 2852.480 ;
        RECT 3123.320 2851.360 3128.040 2852.480 ;
        RECT 3077.280 2848.640 3080.000 2849.760 ;
        RECT 3117.320 2848.640 3122.040 2849.760 ;
        RECT 3072.480 2845.920 3075.200 2847.040 ;
        RECT 3111.320 2845.920 3116.040 2847.040 ;
        RECT 3067.680 2843.200 3070.400 2844.320 ;
        RECT 3105.320 2843.200 3110.040 2844.320 ;
        RECT 3062.880 2840.480 3065.600 2841.600 ;
        RECT 3099.320 2840.480 3104.040 2841.600 ;
        RECT 3058.080 2837.760 3060.800 2838.880 ;
        RECT 3093.320 2837.760 3098.040 2838.880 ;
        RECT 23.060 2835.040 27.780 2836.160 ;
        RECT 111.900 2835.040 114.620 2836.160 ;
        RECT 29.060 2832.320 33.780 2833.440 ;
        RECT 107.100 2832.320 109.820 2833.440 ;
        RECT 35.060 2829.600 39.780 2830.720 ;
        RECT 78.300 2829.600 81.020 2830.720 ;
        RECT 41.060 2826.880 45.780 2828.000 ;
        RECT 83.100 2826.880 85.820 2828.000 ;
        RECT 47.060 2824.160 51.780 2825.280 ;
        RECT 87.900 2824.160 90.620 2825.280 ;
        RECT 53.060 2821.440 57.780 2822.560 ;
        RECT 92.700 2821.440 95.420 2822.560 ;
        RECT 59.060 2818.720 63.780 2819.840 ;
        RECT 97.500 2818.720 100.220 2819.840 ;
        RECT 65.060 2816.000 69.780 2817.120 ;
        RECT 102.300 2816.000 105.020 2817.120 ;
        RECT 3048.480 2791.520 3051.200 2792.640 ;
        RECT 3135.320 2791.520 3140.040 2792.640 ;
        RECT 3053.280 2788.800 3056.000 2789.920 ;
        RECT 3129.320 2788.800 3134.040 2789.920 ;
        RECT 3082.080 2786.080 3084.800 2787.200 ;
        RECT 3123.320 2786.080 3128.040 2787.200 ;
        RECT 3077.280 2783.360 3080.000 2784.480 ;
        RECT 3117.320 2783.360 3122.040 2784.480 ;
        RECT 3072.480 2780.640 3075.200 2781.760 ;
        RECT 3111.320 2780.640 3116.040 2781.760 ;
        RECT 3067.680 2777.920 3070.400 2779.040 ;
        RECT 3105.320 2777.920 3110.040 2779.040 ;
        RECT 3062.880 2775.200 3065.600 2776.320 ;
        RECT 3099.320 2775.200 3104.040 2776.320 ;
        RECT 3058.080 2772.480 3060.800 2773.600 ;
        RECT 3093.320 2772.480 3098.040 2773.600 ;
        RECT 23.060 2758.880 27.780 2760.000 ;
        RECT 111.900 2758.880 114.620 2760.000 ;
        RECT 29.060 2756.160 33.780 2757.280 ;
        RECT 107.100 2756.160 109.820 2757.280 ;
        RECT 35.060 2753.440 39.780 2754.560 ;
        RECT 78.300 2753.440 81.020 2754.560 ;
        RECT 41.060 2750.720 45.780 2751.840 ;
        RECT 83.100 2750.720 85.820 2751.840 ;
        RECT 47.060 2748.000 51.780 2749.120 ;
        RECT 87.900 2748.000 90.620 2749.120 ;
        RECT 53.060 2745.280 57.780 2746.400 ;
        RECT 92.700 2745.280 95.420 2746.400 ;
        RECT 59.060 2742.560 63.780 2743.680 ;
        RECT 97.500 2742.560 100.220 2743.680 ;
        RECT 65.060 2739.840 69.780 2740.960 ;
        RECT 102.300 2739.840 105.020 2740.960 ;
        RECT 3072.480 2715.360 3075.200 2716.480 ;
        RECT 3111.320 2715.360 3116.040 2716.480 ;
        RECT 3067.680 2712.640 3070.400 2713.760 ;
        RECT 3105.320 2712.640 3110.040 2713.760 ;
        RECT 3062.880 2709.920 3065.600 2711.040 ;
        RECT 3099.320 2709.920 3104.040 2711.040 ;
        RECT 3058.080 2707.200 3060.800 2708.320 ;
        RECT 3093.320 2707.200 3098.040 2708.320 ;
        RECT 23.060 2693.600 27.780 2694.720 ;
        RECT 111.900 2693.600 114.620 2694.720 ;
        RECT 29.060 2690.880 33.780 2692.000 ;
        RECT 107.100 2690.880 109.820 2692.000 ;
        RECT 35.060 2688.160 39.780 2689.280 ;
        RECT 78.300 2688.160 81.020 2689.280 ;
        RECT 41.060 2685.440 45.780 2686.560 ;
        RECT 83.100 2685.440 85.820 2686.560 ;
        RECT 47.060 2682.720 51.780 2683.840 ;
        RECT 87.900 2682.720 90.620 2683.840 ;
        RECT 53.060 2680.000 57.780 2681.120 ;
        RECT 92.700 2680.000 95.420 2681.120 ;
        RECT 59.060 2677.280 63.780 2678.400 ;
        RECT 97.500 2677.280 100.220 2678.400 ;
        RECT 65.060 2674.560 69.780 2675.680 ;
        RECT 102.300 2674.560 105.020 2675.680 ;
        RECT 3048.480 2652.800 3051.200 2653.920 ;
        RECT 3135.320 2652.800 3140.040 2653.920 ;
        RECT 3053.280 2650.080 3056.000 2651.200 ;
        RECT 3129.320 2650.080 3134.040 2651.200 ;
        RECT 3082.080 2647.360 3084.800 2648.480 ;
        RECT 3123.320 2647.360 3128.040 2648.480 ;
        RECT 3077.280 2644.640 3080.000 2645.760 ;
        RECT 3117.320 2644.640 3122.040 2645.760 ;
        RECT 3072.480 2641.920 3075.200 2643.040 ;
        RECT 3111.320 2641.920 3116.040 2643.040 ;
        RECT 3067.680 2639.200 3070.400 2640.320 ;
        RECT 3105.320 2639.200 3110.040 2640.320 ;
        RECT 3062.880 2636.480 3065.600 2637.600 ;
        RECT 3099.320 2636.480 3104.040 2637.600 ;
        RECT 3058.080 2633.760 3060.800 2634.880 ;
        RECT 3093.320 2633.760 3098.040 2634.880 ;
        RECT 23.060 2628.320 27.780 2629.440 ;
        RECT 111.900 2628.320 114.620 2629.440 ;
        RECT 29.060 2625.600 33.780 2626.720 ;
        RECT 107.100 2625.600 109.820 2626.720 ;
        RECT 35.060 2622.880 39.780 2624.000 ;
        RECT 78.300 2622.880 81.020 2624.000 ;
        RECT 41.060 2620.160 45.780 2621.280 ;
        RECT 83.100 2620.160 85.820 2621.280 ;
        RECT 47.060 2617.440 51.780 2618.560 ;
        RECT 87.900 2617.440 90.620 2618.560 ;
        RECT 53.060 2614.720 57.780 2615.840 ;
        RECT 92.700 2614.720 95.420 2615.840 ;
        RECT 59.060 2612.000 63.780 2613.120 ;
        RECT 97.500 2612.000 100.220 2613.120 ;
        RECT 65.060 2609.280 69.780 2610.400 ;
        RECT 102.300 2609.280 105.020 2610.400 ;
        RECT 3048.480 2587.520 3051.200 2588.640 ;
        RECT 3135.320 2587.520 3140.040 2588.640 ;
        RECT 3053.280 2584.800 3056.000 2585.920 ;
        RECT 3129.320 2584.800 3134.040 2585.920 ;
        RECT 3082.080 2582.080 3084.800 2583.200 ;
        RECT 3123.320 2582.080 3128.040 2583.200 ;
        RECT 3077.280 2579.360 3080.000 2580.480 ;
        RECT 3117.320 2579.360 3122.040 2580.480 ;
        RECT 3072.480 2576.640 3075.200 2577.760 ;
        RECT 3111.320 2576.640 3116.040 2577.760 ;
        RECT 3067.680 2573.920 3070.400 2575.040 ;
        RECT 3105.320 2573.920 3110.040 2575.040 ;
        RECT 3062.880 2571.200 3065.600 2572.320 ;
        RECT 3099.320 2571.200 3104.040 2572.320 ;
        RECT 3058.080 2568.480 3060.800 2569.600 ;
        RECT 3093.320 2568.480 3098.040 2569.600 ;
        RECT 23.060 2563.040 27.780 2564.160 ;
        RECT 111.900 2563.040 114.620 2564.160 ;
        RECT 29.060 2560.320 33.780 2561.440 ;
        RECT 107.100 2560.320 109.820 2561.440 ;
        RECT 35.060 2557.600 39.780 2558.720 ;
        RECT 78.300 2557.600 81.020 2558.720 ;
        RECT 41.060 2554.880 45.780 2556.000 ;
        RECT 83.100 2554.880 85.820 2556.000 ;
        RECT 47.060 2552.160 51.780 2553.280 ;
        RECT 87.900 2552.160 90.620 2553.280 ;
        RECT 53.060 2549.440 57.780 2550.560 ;
        RECT 92.700 2549.440 95.420 2550.560 ;
        RECT 59.060 2546.720 63.780 2547.840 ;
        RECT 97.500 2546.720 100.220 2547.840 ;
        RECT 65.060 2544.000 69.780 2545.120 ;
        RECT 102.300 2544.000 105.020 2545.120 ;
        RECT 3048.480 2522.240 3051.200 2523.360 ;
        RECT 3135.320 2522.240 3140.040 2523.360 ;
        RECT 3053.280 2519.520 3056.000 2520.640 ;
        RECT 3129.320 2519.520 3134.040 2520.640 ;
        RECT 3082.080 2516.800 3084.800 2517.920 ;
        RECT 3123.320 2516.800 3128.040 2517.920 ;
        RECT 3077.280 2514.080 3080.000 2515.200 ;
        RECT 3117.320 2514.080 3122.040 2515.200 ;
        RECT 3072.480 2511.360 3075.200 2512.480 ;
        RECT 3111.320 2511.360 3116.040 2512.480 ;
        RECT 3067.680 2508.640 3070.400 2509.760 ;
        RECT 3105.320 2508.640 3110.040 2509.760 ;
        RECT 3062.880 2505.920 3065.600 2507.040 ;
        RECT 3099.320 2505.920 3104.040 2507.040 ;
        RECT 3058.080 2503.200 3060.800 2504.320 ;
        RECT 3093.320 2503.200 3098.040 2504.320 ;
        RECT 23.060 2497.760 27.780 2498.880 ;
        RECT 111.900 2497.760 114.620 2498.880 ;
        RECT 29.060 2495.040 33.780 2496.160 ;
        RECT 107.100 2495.040 109.820 2496.160 ;
        RECT 35.060 2492.320 39.780 2493.440 ;
        RECT 78.300 2492.320 81.020 2493.440 ;
        RECT 41.060 2489.600 45.780 2490.720 ;
        RECT 83.100 2489.600 85.820 2490.720 ;
        RECT 47.060 2486.880 51.780 2488.000 ;
        RECT 87.900 2486.880 90.620 2488.000 ;
        RECT 53.060 2484.160 57.780 2485.280 ;
        RECT 92.700 2484.160 95.420 2485.280 ;
        RECT 59.060 2481.440 63.780 2482.560 ;
        RECT 97.500 2481.440 100.220 2482.560 ;
        RECT 65.060 2478.720 69.780 2479.840 ;
        RECT 102.300 2478.720 105.020 2479.840 ;
        RECT 3048.480 2456.960 3051.200 2458.080 ;
        RECT 3135.320 2456.960 3140.040 2458.080 ;
        RECT 3053.280 2454.240 3056.000 2455.360 ;
        RECT 3129.320 2454.240 3134.040 2455.360 ;
        RECT 3082.080 2451.520 3084.800 2452.640 ;
        RECT 3123.320 2451.520 3128.040 2452.640 ;
        RECT 3077.280 2448.800 3080.000 2449.920 ;
        RECT 3117.320 2448.800 3122.040 2449.920 ;
        RECT 3072.480 2446.080 3075.200 2447.200 ;
        RECT 3111.320 2446.080 3116.040 2447.200 ;
        RECT 3067.680 2443.360 3070.400 2444.480 ;
        RECT 3105.320 2443.360 3110.040 2444.480 ;
        RECT 3062.880 2440.640 3065.600 2441.760 ;
        RECT 3099.320 2440.640 3104.040 2441.760 ;
        RECT 3058.080 2437.920 3060.800 2439.040 ;
        RECT 3093.320 2437.920 3098.040 2439.040 ;
        RECT 23.060 2432.480 27.780 2433.600 ;
        RECT 111.900 2432.480 114.620 2433.600 ;
        RECT 29.060 2429.760 33.780 2430.880 ;
        RECT 107.100 2429.760 109.820 2430.880 ;
        RECT 35.060 2427.040 39.780 2428.160 ;
        RECT 78.300 2427.040 81.020 2428.160 ;
        RECT 41.060 2424.320 45.780 2425.440 ;
        RECT 83.100 2424.320 85.820 2425.440 ;
        RECT 47.060 2421.600 51.780 2422.720 ;
        RECT 87.900 2421.600 90.620 2422.720 ;
        RECT 53.060 2418.880 57.780 2420.000 ;
        RECT 92.700 2418.880 95.420 2420.000 ;
        RECT 59.060 2416.160 63.780 2417.280 ;
        RECT 97.500 2416.160 100.220 2417.280 ;
        RECT 65.060 2413.440 69.780 2414.560 ;
        RECT 102.300 2413.440 105.020 2414.560 ;
        RECT 3048.480 2383.520 3051.200 2384.640 ;
        RECT 3135.320 2383.520 3140.040 2384.640 ;
        RECT 3053.280 2380.800 3056.000 2381.920 ;
        RECT 3129.320 2380.800 3134.040 2381.920 ;
        RECT 3082.080 2378.080 3084.800 2379.200 ;
        RECT 3123.320 2378.080 3128.040 2379.200 ;
        RECT 3077.280 2375.360 3080.000 2376.480 ;
        RECT 3117.320 2375.360 3122.040 2376.480 ;
        RECT 3072.480 2372.640 3075.200 2373.760 ;
        RECT 3111.320 2372.640 3116.040 2373.760 ;
        RECT 3067.680 2369.920 3070.400 2371.040 ;
        RECT 3105.320 2369.920 3110.040 2371.040 ;
        RECT 3062.880 2367.200 3065.600 2368.320 ;
        RECT 3099.320 2367.200 3104.040 2368.320 ;
        RECT 3058.080 2364.480 3060.800 2365.600 ;
        RECT 3093.320 2364.480 3098.040 2365.600 ;
        RECT 23.060 2356.320 27.780 2357.440 ;
        RECT 111.900 2356.320 114.620 2357.440 ;
        RECT 29.060 2353.600 33.780 2354.720 ;
        RECT 107.100 2353.600 109.820 2354.720 ;
        RECT 35.060 2350.880 39.780 2352.000 ;
        RECT 78.300 2350.880 81.020 2352.000 ;
        RECT 41.060 2348.160 45.780 2349.280 ;
        RECT 83.100 2348.160 85.820 2349.280 ;
        RECT 47.060 2345.440 51.780 2346.560 ;
        RECT 87.900 2345.440 90.620 2346.560 ;
        RECT 53.060 2342.720 57.780 2343.840 ;
        RECT 92.700 2342.720 95.420 2343.840 ;
        RECT 59.060 2340.000 63.780 2341.120 ;
        RECT 97.500 2340.000 100.220 2341.120 ;
        RECT 65.060 2337.280 69.780 2338.400 ;
        RECT 102.300 2337.280 105.020 2338.400 ;
        RECT 3048.480 2318.240 3051.200 2319.360 ;
        RECT 3135.320 2318.240 3140.040 2319.360 ;
        RECT 3053.280 2315.520 3056.000 2316.640 ;
        RECT 3129.320 2315.520 3134.040 2316.640 ;
        RECT 3082.080 2312.800 3084.800 2313.920 ;
        RECT 3123.320 2312.800 3128.040 2313.920 ;
        RECT 3077.280 2310.080 3080.000 2311.200 ;
        RECT 3117.320 2310.080 3122.040 2311.200 ;
        RECT 3072.480 2307.360 3075.200 2308.480 ;
        RECT 3111.320 2307.360 3116.040 2308.480 ;
        RECT 3067.680 2304.640 3070.400 2305.760 ;
        RECT 3105.320 2304.640 3110.040 2305.760 ;
        RECT 23.060 2301.920 27.780 2303.040 ;
        RECT 111.900 2301.920 114.620 2303.040 ;
        RECT 3062.880 2301.920 3065.600 2303.040 ;
        RECT 3099.320 2301.920 3104.040 2303.040 ;
        RECT 29.060 2299.200 33.780 2300.320 ;
        RECT 107.100 2299.200 109.820 2300.320 ;
        RECT 3058.080 2299.200 3060.800 2300.320 ;
        RECT 3093.320 2299.200 3098.040 2300.320 ;
        RECT 35.060 2296.480 39.780 2297.600 ;
        RECT 78.300 2296.480 81.020 2297.600 ;
        RECT 41.060 2293.760 45.780 2294.880 ;
        RECT 83.100 2293.760 85.820 2294.880 ;
        RECT 47.060 2291.040 51.780 2292.160 ;
        RECT 87.900 2291.040 90.620 2292.160 ;
        RECT 53.060 2288.320 57.780 2289.440 ;
        RECT 92.700 2288.320 95.420 2289.440 ;
        RECT 59.060 2285.600 63.780 2286.720 ;
        RECT 97.500 2285.600 100.220 2286.720 ;
        RECT 65.060 2282.880 69.780 2284.000 ;
        RECT 102.300 2282.880 105.020 2284.000 ;
        RECT 3048.480 2252.960 3051.200 2254.080 ;
        RECT 3135.320 2252.960 3140.040 2254.080 ;
        RECT 3053.280 2250.240 3056.000 2251.360 ;
        RECT 3129.320 2250.240 3134.040 2251.360 ;
        RECT 3082.080 2247.520 3084.800 2248.640 ;
        RECT 3123.320 2247.520 3128.040 2248.640 ;
        RECT 3077.280 2244.800 3080.000 2245.920 ;
        RECT 3117.320 2244.800 3122.040 2245.920 ;
        RECT 3072.480 2242.080 3075.200 2243.200 ;
        RECT 3111.320 2242.080 3116.040 2243.200 ;
        RECT 3067.680 2239.360 3070.400 2240.480 ;
        RECT 3105.320 2239.360 3110.040 2240.480 ;
        RECT 23.060 2236.640 27.780 2237.760 ;
        RECT 111.900 2236.640 114.620 2237.760 ;
        RECT 3062.880 2236.640 3065.600 2237.760 ;
        RECT 3099.320 2236.640 3104.040 2237.760 ;
        RECT 29.060 2233.920 33.780 2235.040 ;
        RECT 107.100 2233.920 109.820 2235.040 ;
        RECT 3058.080 2233.920 3060.800 2235.040 ;
        RECT 3093.320 2233.920 3098.040 2235.040 ;
        RECT 35.060 2231.200 39.780 2232.320 ;
        RECT 78.300 2231.200 81.020 2232.320 ;
        RECT 41.060 2228.480 45.780 2229.600 ;
        RECT 83.100 2228.480 85.820 2229.600 ;
        RECT 47.060 2225.760 51.780 2226.880 ;
        RECT 87.900 2225.760 90.620 2226.880 ;
        RECT 53.060 2223.040 57.780 2224.160 ;
        RECT 92.700 2223.040 95.420 2224.160 ;
        RECT 59.060 2220.320 63.780 2221.440 ;
        RECT 97.500 2220.320 100.220 2221.440 ;
        RECT 65.060 2217.600 69.780 2218.720 ;
        RECT 102.300 2217.600 105.020 2218.720 ;
        RECT 3048.480 2187.680 3051.200 2188.800 ;
        RECT 3135.320 2187.680 3140.040 2188.800 ;
        RECT 3053.280 2184.960 3056.000 2186.080 ;
        RECT 3129.320 2184.960 3134.040 2186.080 ;
        RECT 3082.080 2182.240 3084.800 2183.360 ;
        RECT 3123.320 2182.240 3128.040 2183.360 ;
        RECT 3077.280 2179.520 3080.000 2180.640 ;
        RECT 3117.320 2179.520 3122.040 2180.640 ;
        RECT 3072.480 2176.800 3075.200 2177.920 ;
        RECT 3111.320 2176.800 3116.040 2177.920 ;
        RECT 3067.680 2174.080 3070.400 2175.200 ;
        RECT 3105.320 2174.080 3110.040 2175.200 ;
        RECT 23.060 2171.360 27.780 2172.480 ;
        RECT 111.900 2171.360 114.620 2172.480 ;
        RECT 3062.880 2171.360 3065.600 2172.480 ;
        RECT 3099.320 2171.360 3104.040 2172.480 ;
        RECT 29.060 2168.640 33.780 2169.760 ;
        RECT 107.100 2168.640 109.820 2169.760 ;
        RECT 3058.080 2168.640 3060.800 2169.760 ;
        RECT 3093.320 2168.640 3098.040 2169.760 ;
        RECT 35.060 2165.920 39.780 2167.040 ;
        RECT 78.300 2165.920 81.020 2167.040 ;
        RECT 41.060 2163.200 45.780 2164.320 ;
        RECT 83.100 2163.200 85.820 2164.320 ;
        RECT 47.060 2160.480 51.780 2161.600 ;
        RECT 87.900 2160.480 90.620 2161.600 ;
        RECT 53.060 2157.760 57.780 2158.880 ;
        RECT 92.700 2157.760 95.420 2158.880 ;
        RECT 59.060 2155.040 63.780 2156.160 ;
        RECT 97.500 2155.040 100.220 2156.160 ;
        RECT 65.060 2152.320 69.780 2153.440 ;
        RECT 102.300 2152.320 105.020 2153.440 ;
        RECT 3048.480 2122.400 3051.200 2123.520 ;
        RECT 3135.320 2122.400 3140.040 2123.520 ;
        RECT 3053.280 2119.680 3056.000 2120.800 ;
        RECT 3129.320 2119.680 3134.040 2120.800 ;
        RECT 3082.080 2116.960 3084.800 2118.080 ;
        RECT 3123.320 2116.960 3128.040 2118.080 ;
        RECT 3077.280 2114.240 3080.000 2115.360 ;
        RECT 3117.320 2114.240 3122.040 2115.360 ;
        RECT 3072.480 2111.520 3075.200 2112.640 ;
        RECT 3111.320 2111.520 3116.040 2112.640 ;
        RECT 3067.680 2108.800 3070.400 2109.920 ;
        RECT 3105.320 2108.800 3110.040 2109.920 ;
        RECT 23.060 2106.080 27.780 2107.200 ;
        RECT 111.900 2106.080 114.620 2107.200 ;
        RECT 3062.880 2106.080 3065.600 2107.200 ;
        RECT 3099.320 2106.080 3104.040 2107.200 ;
        RECT 29.060 2103.360 33.780 2104.480 ;
        RECT 107.100 2103.360 109.820 2104.480 ;
        RECT 3058.080 2103.360 3060.800 2104.480 ;
        RECT 3093.320 2103.360 3098.040 2104.480 ;
        RECT 35.060 2100.640 39.780 2101.760 ;
        RECT 78.300 2100.640 81.020 2101.760 ;
        RECT 41.060 2097.920 45.780 2099.040 ;
        RECT 83.100 2097.920 85.820 2099.040 ;
        RECT 47.060 2095.200 51.780 2096.320 ;
        RECT 87.900 2095.200 90.620 2096.320 ;
        RECT 53.060 2092.480 57.780 2093.600 ;
        RECT 92.700 2092.480 95.420 2093.600 ;
        RECT 59.060 2089.760 63.780 2090.880 ;
        RECT 97.500 2089.760 100.220 2090.880 ;
        RECT 65.060 2087.040 69.780 2088.160 ;
        RECT 102.300 2087.040 105.020 2088.160 ;
        RECT 3048.480 2057.120 3051.200 2058.240 ;
        RECT 3135.320 2057.120 3140.040 2058.240 ;
        RECT 3053.280 2054.400 3056.000 2055.520 ;
        RECT 3129.320 2054.400 3134.040 2055.520 ;
        RECT 3082.080 2051.680 3084.800 2052.800 ;
        RECT 3123.320 2051.680 3128.040 2052.800 ;
        RECT 3077.280 2048.960 3080.000 2050.080 ;
        RECT 3117.320 2048.960 3122.040 2050.080 ;
        RECT 3072.480 2046.240 3075.200 2047.360 ;
        RECT 3111.320 2046.240 3116.040 2047.360 ;
        RECT 3067.680 2043.520 3070.400 2044.640 ;
        RECT 3105.320 2043.520 3110.040 2044.640 ;
        RECT 23.060 2040.800 27.780 2041.920 ;
        RECT 111.900 2040.800 114.620 2041.920 ;
        RECT 3062.880 2040.800 3065.600 2041.920 ;
        RECT 3099.320 2040.800 3104.040 2041.920 ;
        RECT 29.060 2038.080 33.780 2039.200 ;
        RECT 107.100 2038.080 109.820 2039.200 ;
        RECT 3058.080 2038.080 3060.800 2039.200 ;
        RECT 3093.320 2038.080 3098.040 2039.200 ;
        RECT 35.060 2035.360 39.780 2036.480 ;
        RECT 78.300 2035.360 81.020 2036.480 ;
        RECT 41.060 2032.640 45.780 2033.760 ;
        RECT 83.100 2032.640 85.820 2033.760 ;
        RECT 47.060 2029.920 51.780 2031.040 ;
        RECT 87.900 2029.920 90.620 2031.040 ;
        RECT 53.060 2027.200 57.780 2028.320 ;
        RECT 92.700 2027.200 95.420 2028.320 ;
        RECT 59.060 2024.480 63.780 2025.600 ;
        RECT 97.500 2024.480 100.220 2025.600 ;
        RECT 65.060 2021.760 69.780 2022.880 ;
        RECT 102.300 2021.760 105.020 2022.880 ;
        RECT 3048.480 1991.840 3051.200 1992.960 ;
        RECT 3135.320 1991.840 3140.040 1992.960 ;
        RECT 3053.280 1989.120 3056.000 1990.240 ;
        RECT 3129.320 1989.120 3134.040 1990.240 ;
        RECT 3082.080 1986.400 3084.800 1987.520 ;
        RECT 3123.320 1986.400 3128.040 1987.520 ;
        RECT 3077.280 1983.680 3080.000 1984.800 ;
        RECT 3117.320 1983.680 3122.040 1984.800 ;
        RECT 3072.480 1980.960 3075.200 1982.080 ;
        RECT 3111.320 1980.960 3116.040 1982.080 ;
        RECT 3067.680 1978.240 3070.400 1979.360 ;
        RECT 3105.320 1978.240 3110.040 1979.360 ;
        RECT 23.060 1975.520 27.780 1976.640 ;
        RECT 111.900 1975.520 114.620 1976.640 ;
        RECT 3062.880 1975.520 3065.600 1976.640 ;
        RECT 3099.320 1975.520 3104.040 1976.640 ;
        RECT 29.060 1972.800 33.780 1973.920 ;
        RECT 107.100 1972.800 109.820 1973.920 ;
        RECT 3058.080 1972.800 3060.800 1973.920 ;
        RECT 3093.320 1972.800 3098.040 1973.920 ;
        RECT 35.060 1970.080 39.780 1971.200 ;
        RECT 78.300 1970.080 81.020 1971.200 ;
        RECT 41.060 1967.360 45.780 1968.480 ;
        RECT 83.100 1967.360 85.820 1968.480 ;
        RECT 47.060 1964.640 51.780 1965.760 ;
        RECT 87.900 1964.640 90.620 1965.760 ;
        RECT 53.060 1961.920 57.780 1963.040 ;
        RECT 92.700 1961.920 95.420 1963.040 ;
        RECT 59.060 1959.200 63.780 1960.320 ;
        RECT 97.500 1959.200 100.220 1960.320 ;
        RECT 65.060 1956.480 69.780 1957.600 ;
        RECT 102.300 1956.480 105.020 1957.600 ;
        RECT 3048.480 1926.560 3051.200 1927.680 ;
        RECT 3135.320 1926.560 3140.040 1927.680 ;
        RECT 3053.280 1923.840 3056.000 1924.960 ;
        RECT 3129.320 1923.840 3134.040 1924.960 ;
        RECT 3082.080 1921.120 3084.800 1922.240 ;
        RECT 3123.320 1921.120 3128.040 1922.240 ;
        RECT 3077.280 1918.400 3080.000 1919.520 ;
        RECT 3117.320 1918.400 3122.040 1919.520 ;
        RECT 3072.480 1915.680 3075.200 1916.800 ;
        RECT 3111.320 1915.680 3116.040 1916.800 ;
        RECT 3067.680 1912.960 3070.400 1914.080 ;
        RECT 3105.320 1912.960 3110.040 1914.080 ;
        RECT 23.060 1910.240 27.780 1911.360 ;
        RECT 111.900 1910.240 114.620 1911.360 ;
        RECT 3062.880 1910.240 3065.600 1911.360 ;
        RECT 3099.320 1910.240 3104.040 1911.360 ;
        RECT 29.060 1907.520 33.780 1908.640 ;
        RECT 107.100 1907.520 109.820 1908.640 ;
        RECT 3058.080 1907.520 3060.800 1908.640 ;
        RECT 3093.320 1907.520 3098.040 1908.640 ;
        RECT 35.060 1904.800 39.780 1905.920 ;
        RECT 78.300 1904.800 81.020 1905.920 ;
        RECT 41.060 1902.080 45.780 1903.200 ;
        RECT 83.100 1902.080 85.820 1903.200 ;
        RECT 47.060 1899.360 51.780 1900.480 ;
        RECT 87.900 1899.360 90.620 1900.480 ;
        RECT 53.060 1896.640 57.780 1897.760 ;
        RECT 92.700 1896.640 95.420 1897.760 ;
        RECT 59.060 1893.920 63.780 1895.040 ;
        RECT 97.500 1893.920 100.220 1895.040 ;
        RECT 65.060 1891.200 69.780 1892.320 ;
        RECT 102.300 1891.200 105.020 1892.320 ;
        RECT 23.060 1844.960 27.780 1846.080 ;
        RECT 111.900 1844.960 114.620 1846.080 ;
        RECT 3048.480 1844.960 3051.200 1846.080 ;
        RECT 3135.320 1844.960 3140.040 1846.080 ;
        RECT 29.060 1842.240 33.780 1843.360 ;
        RECT 107.100 1842.240 109.820 1843.360 ;
        RECT 3053.280 1842.240 3056.000 1843.360 ;
        RECT 3129.320 1842.240 3134.040 1843.360 ;
        RECT 35.060 1839.520 39.780 1840.640 ;
        RECT 78.300 1839.520 81.020 1840.640 ;
        RECT 3082.080 1839.520 3084.800 1840.640 ;
        RECT 3123.320 1839.520 3128.040 1840.640 ;
        RECT 41.060 1836.800 45.780 1837.920 ;
        RECT 83.100 1836.800 85.820 1837.920 ;
        RECT 3077.280 1836.800 3080.000 1837.920 ;
        RECT 3117.320 1836.800 3122.040 1837.920 ;
        RECT 47.060 1834.080 51.780 1835.200 ;
        RECT 87.900 1834.080 90.620 1835.200 ;
        RECT 3072.480 1834.080 3075.200 1835.200 ;
        RECT 3111.320 1834.080 3116.040 1835.200 ;
        RECT 53.060 1831.360 57.780 1832.480 ;
        RECT 92.700 1831.360 95.420 1832.480 ;
        RECT 3067.680 1831.360 3070.400 1832.480 ;
        RECT 3105.320 1831.360 3110.040 1832.480 ;
        RECT 59.060 1828.640 63.780 1829.760 ;
        RECT 97.500 1828.640 100.220 1829.760 ;
        RECT 3062.880 1828.640 3065.600 1829.760 ;
        RECT 3099.320 1828.640 3104.040 1829.760 ;
        RECT 65.060 1825.920 69.780 1827.040 ;
        RECT 102.300 1825.920 105.020 1827.040 ;
        RECT 3058.080 1825.920 3060.800 1827.040 ;
        RECT 3093.320 1825.920 3098.040 1827.040 ;
        RECT 23.060 1779.680 27.780 1780.800 ;
        RECT 111.900 1779.680 114.620 1780.800 ;
        RECT 3048.480 1779.680 3051.200 1780.800 ;
        RECT 3135.320 1779.680 3140.040 1780.800 ;
        RECT 29.060 1776.960 33.780 1778.080 ;
        RECT 107.100 1776.960 109.820 1778.080 ;
        RECT 3053.280 1776.960 3056.000 1778.080 ;
        RECT 3129.320 1776.960 3134.040 1778.080 ;
        RECT 35.060 1774.240 39.780 1775.360 ;
        RECT 78.300 1774.240 81.020 1775.360 ;
        RECT 3082.080 1774.240 3084.800 1775.360 ;
        RECT 3123.320 1774.240 3128.040 1775.360 ;
        RECT 41.060 1771.520 45.780 1772.640 ;
        RECT 83.100 1771.520 85.820 1772.640 ;
        RECT 3077.280 1771.520 3080.000 1772.640 ;
        RECT 3117.320 1771.520 3122.040 1772.640 ;
        RECT 47.060 1768.800 51.780 1769.920 ;
        RECT 87.900 1768.800 90.620 1769.920 ;
        RECT 3072.480 1768.800 3075.200 1769.920 ;
        RECT 3111.320 1768.800 3116.040 1769.920 ;
        RECT 53.060 1766.080 57.780 1767.200 ;
        RECT 92.700 1766.080 95.420 1767.200 ;
        RECT 3067.680 1766.080 3070.400 1767.200 ;
        RECT 3105.320 1766.080 3110.040 1767.200 ;
        RECT 59.060 1763.360 63.780 1764.480 ;
        RECT 97.500 1763.360 100.220 1764.480 ;
        RECT 3062.880 1763.360 3065.600 1764.480 ;
        RECT 3099.320 1763.360 3104.040 1764.480 ;
        RECT 65.060 1760.640 69.780 1761.760 ;
        RECT 102.300 1760.640 105.020 1761.760 ;
        RECT 3058.080 1760.640 3060.800 1761.760 ;
        RECT 3093.320 1760.640 3098.040 1761.760 ;
        RECT 3048.480 1714.400 3051.200 1715.520 ;
        RECT 3135.320 1714.400 3140.040 1715.520 ;
        RECT 3053.280 1711.680 3056.000 1712.800 ;
        RECT 3129.320 1711.680 3134.040 1712.800 ;
        RECT 3082.080 1708.960 3084.800 1710.080 ;
        RECT 3123.320 1708.960 3128.040 1710.080 ;
        RECT 3077.280 1706.240 3080.000 1707.360 ;
        RECT 3117.320 1706.240 3122.040 1707.360 ;
        RECT 23.060 1703.520 27.780 1704.640 ;
        RECT 111.900 1703.520 114.620 1704.640 ;
        RECT 3072.480 1703.520 3075.200 1704.640 ;
        RECT 3111.320 1703.520 3116.040 1704.640 ;
        RECT 29.060 1700.800 33.780 1701.920 ;
        RECT 107.100 1700.800 109.820 1701.920 ;
        RECT 3067.680 1700.800 3070.400 1701.920 ;
        RECT 3105.320 1700.800 3110.040 1701.920 ;
        RECT 35.060 1698.080 39.780 1699.200 ;
        RECT 78.300 1698.080 81.020 1699.200 ;
        RECT 3062.880 1698.080 3065.600 1699.200 ;
        RECT 3099.320 1698.080 3104.040 1699.200 ;
        RECT 41.060 1695.360 45.780 1696.480 ;
        RECT 83.100 1695.360 85.820 1696.480 ;
        RECT 3058.080 1695.360 3060.800 1696.480 ;
        RECT 3093.320 1695.360 3098.040 1696.480 ;
        RECT 47.060 1692.640 51.780 1693.760 ;
        RECT 87.900 1692.640 90.620 1693.760 ;
        RECT 53.060 1689.920 57.780 1691.040 ;
        RECT 92.700 1689.920 95.420 1691.040 ;
        RECT 59.060 1687.200 63.780 1688.320 ;
        RECT 97.500 1687.200 100.220 1688.320 ;
        RECT 65.060 1684.480 69.780 1685.600 ;
        RECT 102.300 1684.480 105.020 1685.600 ;
        RECT 23.060 1649.120 27.780 1650.240 ;
        RECT 111.900 1649.120 114.620 1650.240 ;
        RECT 3048.480 1649.120 3051.200 1650.240 ;
        RECT 3135.320 1649.120 3140.040 1650.240 ;
        RECT 29.060 1646.400 33.780 1647.520 ;
        RECT 107.100 1646.400 109.820 1647.520 ;
        RECT 3053.280 1646.400 3056.000 1647.520 ;
        RECT 3129.320 1646.400 3134.040 1647.520 ;
        RECT 35.060 1643.680 39.780 1644.800 ;
        RECT 78.300 1643.680 81.020 1644.800 ;
        RECT 3082.080 1643.680 3084.800 1644.800 ;
        RECT 3123.320 1643.680 3128.040 1644.800 ;
        RECT 41.060 1640.960 45.780 1642.080 ;
        RECT 83.100 1640.960 85.820 1642.080 ;
        RECT 3077.280 1640.960 3080.000 1642.080 ;
        RECT 3117.320 1640.960 3122.040 1642.080 ;
        RECT 47.060 1638.240 51.780 1639.360 ;
        RECT 87.900 1638.240 90.620 1639.360 ;
        RECT 3072.480 1638.240 3075.200 1639.360 ;
        RECT 3111.320 1638.240 3116.040 1639.360 ;
        RECT 53.060 1635.520 57.780 1636.640 ;
        RECT 92.700 1635.520 95.420 1636.640 ;
        RECT 3067.680 1635.520 3070.400 1636.640 ;
        RECT 3105.320 1635.520 3110.040 1636.640 ;
        RECT 59.060 1632.800 63.780 1633.920 ;
        RECT 97.500 1632.800 100.220 1633.920 ;
        RECT 3062.880 1632.800 3065.600 1633.920 ;
        RECT 3099.320 1632.800 3104.040 1633.920 ;
        RECT 65.060 1630.080 69.780 1631.200 ;
        RECT 102.300 1630.080 105.020 1631.200 ;
        RECT 3058.080 1630.080 3060.800 1631.200 ;
        RECT 3093.320 1630.080 3098.040 1631.200 ;
        RECT 3048.480 1592.000 3051.200 1593.120 ;
        RECT 3135.320 1592.000 3140.040 1593.120 ;
        RECT 3053.280 1589.280 3056.000 1590.400 ;
        RECT 3129.320 1589.280 3134.040 1590.400 ;
        RECT 3082.080 1586.560 3084.800 1587.680 ;
        RECT 3123.320 1586.560 3128.040 1587.680 ;
        RECT 23.060 1583.840 27.780 1584.960 ;
        RECT 111.900 1583.840 114.620 1584.960 ;
        RECT 3077.280 1583.840 3080.000 1584.960 ;
        RECT 3117.320 1583.840 3122.040 1584.960 ;
        RECT 29.060 1581.120 33.780 1582.240 ;
        RECT 107.100 1581.120 109.820 1582.240 ;
        RECT 3072.480 1581.120 3075.200 1582.240 ;
        RECT 3111.320 1581.120 3116.040 1582.240 ;
        RECT 35.060 1578.400 39.780 1579.520 ;
        RECT 78.300 1578.400 81.020 1579.520 ;
        RECT 3067.680 1578.400 3070.400 1579.520 ;
        RECT 3105.320 1578.400 3110.040 1579.520 ;
        RECT 41.060 1575.680 45.780 1576.800 ;
        RECT 83.100 1575.680 85.820 1576.800 ;
        RECT 3062.880 1575.680 3065.600 1576.800 ;
        RECT 3099.320 1575.680 3104.040 1576.800 ;
        RECT 47.060 1572.960 51.780 1574.080 ;
        RECT 87.900 1572.960 90.620 1574.080 ;
        RECT 3058.080 1572.960 3060.800 1574.080 ;
        RECT 3093.320 1572.960 3098.040 1574.080 ;
        RECT 53.060 1570.240 57.780 1571.360 ;
        RECT 92.700 1570.240 95.420 1571.360 ;
        RECT 59.060 1567.520 63.780 1568.640 ;
        RECT 97.500 1567.520 100.220 1568.640 ;
        RECT 65.060 1564.800 69.780 1565.920 ;
        RECT 102.300 1564.800 105.020 1565.920 ;
        RECT 23.060 1529.440 27.780 1530.560 ;
        RECT 111.900 1529.440 114.620 1530.560 ;
        RECT 29.060 1526.720 33.780 1527.840 ;
        RECT 107.100 1526.720 109.820 1527.840 ;
        RECT 35.060 1524.000 39.780 1525.120 ;
        RECT 78.300 1524.000 81.020 1525.120 ;
        RECT 41.060 1521.280 45.780 1522.400 ;
        RECT 83.100 1521.280 85.820 1522.400 ;
        RECT 47.060 1518.560 51.780 1519.680 ;
        RECT 87.900 1518.560 90.620 1519.680 ;
        RECT 3048.480 1518.560 3051.200 1519.680 ;
        RECT 3135.320 1518.560 3140.040 1519.680 ;
        RECT 53.060 1515.840 57.780 1516.960 ;
        RECT 92.700 1515.840 95.420 1516.960 ;
        RECT 3053.280 1515.840 3056.000 1516.960 ;
        RECT 3129.320 1515.840 3134.040 1516.960 ;
        RECT 59.060 1513.120 63.780 1514.240 ;
        RECT 97.500 1513.120 100.220 1514.240 ;
        RECT 3082.080 1513.120 3084.800 1514.240 ;
        RECT 3123.320 1513.120 3128.040 1514.240 ;
        RECT 65.060 1510.400 69.780 1511.520 ;
        RECT 102.300 1510.400 105.020 1511.520 ;
        RECT 3077.280 1510.400 3080.000 1511.520 ;
        RECT 3117.320 1510.400 3122.040 1511.520 ;
        RECT 3072.480 1507.680 3075.200 1508.800 ;
        RECT 3111.320 1507.680 3116.040 1508.800 ;
        RECT 3067.680 1504.960 3070.400 1506.080 ;
        RECT 3105.320 1504.960 3110.040 1506.080 ;
        RECT 3062.880 1502.240 3065.600 1503.360 ;
        RECT 3099.320 1502.240 3104.040 1503.360 ;
        RECT 3058.080 1499.520 3060.800 1500.640 ;
        RECT 3093.320 1499.520 3098.040 1500.640 ;
        RECT 23.060 1453.280 27.780 1454.400 ;
        RECT 111.900 1453.280 114.620 1454.400 ;
        RECT 3048.480 1453.280 3051.200 1454.400 ;
        RECT 3135.320 1453.280 3140.040 1454.400 ;
        RECT 29.060 1450.560 33.780 1451.680 ;
        RECT 107.100 1450.560 109.820 1451.680 ;
        RECT 3053.280 1450.560 3056.000 1451.680 ;
        RECT 3129.320 1450.560 3134.040 1451.680 ;
        RECT 35.060 1447.840 39.780 1448.960 ;
        RECT 78.300 1447.840 81.020 1448.960 ;
        RECT 3082.080 1447.840 3084.800 1448.960 ;
        RECT 3123.320 1447.840 3128.040 1448.960 ;
        RECT 41.060 1445.120 45.780 1446.240 ;
        RECT 83.100 1445.120 85.820 1446.240 ;
        RECT 3077.280 1445.120 3080.000 1446.240 ;
        RECT 3117.320 1445.120 3122.040 1446.240 ;
        RECT 47.060 1442.400 51.780 1443.520 ;
        RECT 87.900 1442.400 90.620 1443.520 ;
        RECT 3072.480 1442.400 3075.200 1443.520 ;
        RECT 3111.320 1442.400 3116.040 1443.520 ;
        RECT 53.060 1439.680 57.780 1440.800 ;
        RECT 92.700 1439.680 95.420 1440.800 ;
        RECT 3067.680 1439.680 3070.400 1440.800 ;
        RECT 3105.320 1439.680 3110.040 1440.800 ;
        RECT 59.060 1436.960 63.780 1438.080 ;
        RECT 97.500 1436.960 100.220 1438.080 ;
        RECT 3062.880 1436.960 3065.600 1438.080 ;
        RECT 3099.320 1436.960 3104.040 1438.080 ;
        RECT 65.060 1434.240 69.780 1435.360 ;
        RECT 102.300 1434.240 105.020 1435.360 ;
        RECT 3058.080 1434.240 3060.800 1435.360 ;
        RECT 3093.320 1434.240 3098.040 1435.360 ;
        RECT 23.060 1388.000 27.780 1389.120 ;
        RECT 111.900 1388.000 114.620 1389.120 ;
        RECT 3048.480 1388.000 3051.200 1389.120 ;
        RECT 3135.320 1388.000 3140.040 1389.120 ;
        RECT 29.060 1385.280 33.780 1386.400 ;
        RECT 107.100 1385.280 109.820 1386.400 ;
        RECT 3053.280 1385.280 3056.000 1386.400 ;
        RECT 3129.320 1385.280 3134.040 1386.400 ;
        RECT 35.060 1382.560 39.780 1383.680 ;
        RECT 78.300 1382.560 81.020 1383.680 ;
        RECT 3082.080 1382.560 3084.800 1383.680 ;
        RECT 3123.320 1382.560 3128.040 1383.680 ;
        RECT 41.060 1379.840 45.780 1380.960 ;
        RECT 83.100 1379.840 85.820 1380.960 ;
        RECT 3077.280 1379.840 3080.000 1380.960 ;
        RECT 3117.320 1379.840 3122.040 1380.960 ;
        RECT 47.060 1377.120 51.780 1378.240 ;
        RECT 87.900 1377.120 90.620 1378.240 ;
        RECT 3072.480 1377.120 3075.200 1378.240 ;
        RECT 3111.320 1377.120 3116.040 1378.240 ;
        RECT 53.060 1374.400 57.780 1375.520 ;
        RECT 92.700 1374.400 95.420 1375.520 ;
        RECT 3067.680 1374.400 3070.400 1375.520 ;
        RECT 3105.320 1374.400 3110.040 1375.520 ;
        RECT 59.060 1371.680 63.780 1372.800 ;
        RECT 97.500 1371.680 100.220 1372.800 ;
        RECT 3062.880 1371.680 3065.600 1372.800 ;
        RECT 3099.320 1371.680 3104.040 1372.800 ;
        RECT 65.060 1368.960 69.780 1370.080 ;
        RECT 102.300 1368.960 105.020 1370.080 ;
        RECT 3058.080 1368.960 3060.800 1370.080 ;
        RECT 3093.320 1368.960 3098.040 1370.080 ;
        RECT 23.060 1333.600 27.780 1334.720 ;
        RECT 111.900 1333.600 114.620 1334.720 ;
        RECT 29.060 1330.880 33.780 1332.000 ;
        RECT 107.100 1330.880 109.820 1332.000 ;
        RECT 35.060 1328.160 39.780 1329.280 ;
        RECT 78.300 1328.160 81.020 1329.280 ;
        RECT 41.060 1325.440 45.780 1326.560 ;
        RECT 83.100 1325.440 85.820 1326.560 ;
        RECT 47.060 1322.720 51.780 1323.840 ;
        RECT 87.900 1322.720 90.620 1323.840 ;
        RECT 53.060 1320.000 57.780 1321.120 ;
        RECT 92.700 1320.000 95.420 1321.120 ;
        RECT 59.060 1317.280 63.780 1318.400 ;
        RECT 97.500 1317.280 100.220 1318.400 ;
        RECT 65.060 1314.560 69.780 1315.680 ;
        RECT 102.300 1314.560 105.020 1315.680 ;
        RECT 3048.480 1314.560 3051.200 1315.680 ;
        RECT 3135.320 1314.560 3140.040 1315.680 ;
        RECT 3053.280 1311.840 3056.000 1312.960 ;
        RECT 3129.320 1311.840 3134.040 1312.960 ;
        RECT 3082.080 1309.120 3084.800 1310.240 ;
        RECT 3123.320 1309.120 3128.040 1310.240 ;
        RECT 3077.280 1306.400 3080.000 1307.520 ;
        RECT 3117.320 1306.400 3122.040 1307.520 ;
        RECT 3072.480 1303.680 3075.200 1304.800 ;
        RECT 3111.320 1303.680 3116.040 1304.800 ;
        RECT 3067.680 1300.960 3070.400 1302.080 ;
        RECT 3105.320 1300.960 3110.040 1302.080 ;
        RECT 3062.880 1298.240 3065.600 1299.360 ;
        RECT 3099.320 1298.240 3104.040 1299.360 ;
        RECT 3058.080 1295.520 3060.800 1296.640 ;
        RECT 3093.320 1295.520 3098.040 1296.640 ;
        RECT 23.060 1257.440 27.780 1258.560 ;
        RECT 111.900 1257.440 114.620 1258.560 ;
        RECT 3048.480 1257.440 3051.200 1258.560 ;
        RECT 3135.320 1257.440 3140.040 1258.560 ;
        RECT 29.060 1254.720 33.780 1255.840 ;
        RECT 107.100 1254.720 109.820 1255.840 ;
        RECT 3053.280 1254.720 3056.000 1255.840 ;
        RECT 3129.320 1254.720 3134.040 1255.840 ;
        RECT 35.060 1252.000 39.780 1253.120 ;
        RECT 78.300 1252.000 81.020 1253.120 ;
        RECT 3082.080 1252.000 3084.800 1253.120 ;
        RECT 3123.320 1252.000 3128.040 1253.120 ;
        RECT 41.060 1249.280 45.780 1250.400 ;
        RECT 83.100 1249.280 85.820 1250.400 ;
        RECT 3077.280 1249.280 3080.000 1250.400 ;
        RECT 3117.320 1249.280 3122.040 1250.400 ;
        RECT 47.060 1246.560 51.780 1247.680 ;
        RECT 87.900 1246.560 90.620 1247.680 ;
        RECT 3072.480 1246.560 3075.200 1247.680 ;
        RECT 3111.320 1246.560 3116.040 1247.680 ;
        RECT 53.060 1243.840 57.780 1244.960 ;
        RECT 92.700 1243.840 95.420 1244.960 ;
        RECT 3067.680 1243.840 3070.400 1244.960 ;
        RECT 3105.320 1243.840 3110.040 1244.960 ;
        RECT 59.060 1241.120 63.780 1242.240 ;
        RECT 97.500 1241.120 100.220 1242.240 ;
        RECT 3062.880 1241.120 3065.600 1242.240 ;
        RECT 3099.320 1241.120 3104.040 1242.240 ;
        RECT 65.060 1238.400 69.780 1239.520 ;
        RECT 102.300 1238.400 105.020 1239.520 ;
        RECT 3058.080 1238.400 3060.800 1239.520 ;
        RECT 3093.320 1238.400 3098.040 1239.520 ;
        RECT 23.060 1192.160 27.780 1193.280 ;
        RECT 111.900 1192.160 114.620 1193.280 ;
        RECT 3048.480 1192.160 3051.200 1193.280 ;
        RECT 3135.320 1192.160 3140.040 1193.280 ;
        RECT 29.060 1189.440 33.780 1190.560 ;
        RECT 107.100 1189.440 109.820 1190.560 ;
        RECT 3053.280 1189.440 3056.000 1190.560 ;
        RECT 3129.320 1189.440 3134.040 1190.560 ;
        RECT 35.060 1186.720 39.780 1187.840 ;
        RECT 78.300 1186.720 81.020 1187.840 ;
        RECT 3082.080 1186.720 3084.800 1187.840 ;
        RECT 3123.320 1186.720 3128.040 1187.840 ;
        RECT 41.060 1184.000 45.780 1185.120 ;
        RECT 83.100 1184.000 85.820 1185.120 ;
        RECT 3077.280 1184.000 3080.000 1185.120 ;
        RECT 3117.320 1184.000 3122.040 1185.120 ;
        RECT 47.060 1181.280 51.780 1182.400 ;
        RECT 87.900 1181.280 90.620 1182.400 ;
        RECT 3072.480 1181.280 3075.200 1182.400 ;
        RECT 3111.320 1181.280 3116.040 1182.400 ;
        RECT 53.060 1178.560 57.780 1179.680 ;
        RECT 92.700 1178.560 95.420 1179.680 ;
        RECT 3067.680 1178.560 3070.400 1179.680 ;
        RECT 3105.320 1178.560 3110.040 1179.680 ;
        RECT 59.060 1175.840 63.780 1176.960 ;
        RECT 97.500 1175.840 100.220 1176.960 ;
        RECT 3062.880 1175.840 3065.600 1176.960 ;
        RECT 3099.320 1175.840 3104.040 1176.960 ;
        RECT 65.060 1173.120 69.780 1174.240 ;
        RECT 102.300 1173.120 105.020 1174.240 ;
        RECT 3058.080 1173.120 3060.800 1174.240 ;
        RECT 3093.320 1173.120 3098.040 1174.240 ;
        RECT 23.060 1126.880 27.780 1128.000 ;
        RECT 111.900 1126.880 114.620 1128.000 ;
        RECT 3048.480 1126.880 3051.200 1128.000 ;
        RECT 3135.320 1126.880 3140.040 1128.000 ;
        RECT 29.060 1124.160 33.780 1125.280 ;
        RECT 107.100 1124.160 109.820 1125.280 ;
        RECT 3053.280 1124.160 3056.000 1125.280 ;
        RECT 3129.320 1124.160 3134.040 1125.280 ;
        RECT 35.060 1121.440 39.780 1122.560 ;
        RECT 78.300 1121.440 81.020 1122.560 ;
        RECT 3082.080 1121.440 3084.800 1122.560 ;
        RECT 3123.320 1121.440 3128.040 1122.560 ;
        RECT 41.060 1118.720 45.780 1119.840 ;
        RECT 83.100 1118.720 85.820 1119.840 ;
        RECT 3077.280 1118.720 3080.000 1119.840 ;
        RECT 3117.320 1118.720 3122.040 1119.840 ;
        RECT 47.060 1116.000 51.780 1117.120 ;
        RECT 87.900 1116.000 90.620 1117.120 ;
        RECT 3072.480 1116.000 3075.200 1117.120 ;
        RECT 3111.320 1116.000 3116.040 1117.120 ;
        RECT 53.060 1113.280 57.780 1114.400 ;
        RECT 92.700 1113.280 95.420 1114.400 ;
        RECT 3067.680 1113.280 3070.400 1114.400 ;
        RECT 3105.320 1113.280 3110.040 1114.400 ;
        RECT 59.060 1110.560 63.780 1111.680 ;
        RECT 97.500 1110.560 100.220 1111.680 ;
        RECT 3062.880 1110.560 3065.600 1111.680 ;
        RECT 3099.320 1110.560 3104.040 1111.680 ;
        RECT 65.060 1107.840 69.780 1108.960 ;
        RECT 102.300 1107.840 105.020 1108.960 ;
        RECT 3058.080 1107.840 3060.800 1108.960 ;
        RECT 3093.320 1107.840 3098.040 1108.960 ;
        RECT 3048.480 1061.600 3051.200 1062.720 ;
        RECT 3135.320 1061.600 3140.040 1062.720 ;
        RECT 3053.280 1058.880 3056.000 1060.000 ;
        RECT 3129.320 1058.880 3134.040 1060.000 ;
        RECT 23.060 1056.160 27.780 1057.280 ;
        RECT 111.900 1056.160 114.620 1057.280 ;
        RECT 3082.080 1056.160 3084.800 1057.280 ;
        RECT 3123.320 1056.160 3128.040 1057.280 ;
        RECT 29.060 1053.440 33.780 1054.560 ;
        RECT 107.100 1053.440 109.820 1054.560 ;
        RECT 3077.280 1053.440 3080.000 1054.560 ;
        RECT 3117.320 1053.440 3122.040 1054.560 ;
        RECT 35.060 1050.720 39.780 1051.840 ;
        RECT 78.300 1050.720 81.020 1051.840 ;
        RECT 3072.480 1050.720 3075.200 1051.840 ;
        RECT 3111.320 1050.720 3116.040 1051.840 ;
        RECT 41.060 1048.000 45.780 1049.120 ;
        RECT 83.100 1048.000 85.820 1049.120 ;
        RECT 3067.680 1048.000 3070.400 1049.120 ;
        RECT 3105.320 1048.000 3110.040 1049.120 ;
        RECT 47.060 1045.280 51.780 1046.400 ;
        RECT 87.900 1045.280 90.620 1046.400 ;
        RECT 3062.880 1045.280 3065.600 1046.400 ;
        RECT 3099.320 1045.280 3104.040 1046.400 ;
        RECT 53.060 1042.560 57.780 1043.680 ;
        RECT 92.700 1042.560 95.420 1043.680 ;
        RECT 3058.080 1042.560 3060.800 1043.680 ;
        RECT 3093.320 1042.560 3098.040 1043.680 ;
        RECT 59.060 1039.840 63.780 1040.960 ;
        RECT 97.500 1039.840 100.220 1040.960 ;
        RECT 65.060 1037.120 69.780 1038.240 ;
        RECT 102.300 1037.120 105.020 1038.240 ;
        RECT 1040.955 135.520 1045.275 136.640 ;
        RECT 1135.355 133.320 1138.075 134.440 ;
        RECT 654.975 38.040 659.295 39.160 ;
        RECT 698.860 37.945 699.580 38.665 ;
        RECT 661.735 34.720 666.055 35.840 ;
        RECT 692.360 35.125 693.080 35.845 ;
      LAYER met4 ;
        RECT 3048.480 4554.080 3051.200 4555.200 ;
        RECT 3135.320 4554.080 3140.040 4555.200 ;
        RECT 3053.280 4551.360 3056.000 4552.480 ;
        RECT 3129.320 4551.360 3134.040 4552.480 ;
        RECT 3082.080 4548.640 3084.800 4549.760 ;
        RECT 3123.320 4548.640 3128.040 4549.760 ;
        RECT 3077.280 4545.920 3080.000 4547.040 ;
        RECT 3117.320 4545.920 3122.040 4547.040 ;
        RECT 3072.480 4543.200 3075.200 4544.320 ;
        RECT 3111.320 4543.200 3116.040 4544.320 ;
        RECT 3067.680 4540.480 3070.400 4541.600 ;
        RECT 3105.320 4540.480 3110.040 4541.600 ;
        RECT 3062.880 4537.760 3065.600 4538.880 ;
        RECT 3099.320 4537.760 3104.040 4538.880 ;
        RECT 3058.080 4535.040 3060.800 4536.160 ;
        RECT 3093.320 4535.040 3098.040 4536.160 ;
        RECT 23.060 4529.600 27.780 4530.720 ;
        RECT 111.900 4529.600 114.620 4530.720 ;
        RECT 29.060 4526.880 33.780 4528.000 ;
        RECT 107.100 4526.880 109.820 4528.000 ;
        RECT 35.060 4524.160 39.780 4525.280 ;
        RECT 78.300 4524.160 81.020 4525.280 ;
        RECT 41.060 4521.440 45.780 4522.560 ;
        RECT 83.100 4521.440 85.820 4522.560 ;
        RECT 47.060 4518.720 51.780 4519.840 ;
        RECT 87.900 4518.720 90.620 4519.840 ;
        RECT 53.060 4516.000 57.780 4517.120 ;
        RECT 92.700 4516.000 95.420 4517.120 ;
        RECT 59.060 4513.280 63.780 4514.400 ;
        RECT 97.500 4513.280 100.220 4514.400 ;
        RECT 65.060 4510.560 69.780 4511.680 ;
        RECT 102.300 4510.560 105.020 4511.680 ;
        RECT 3048.480 4480.640 3051.200 4481.760 ;
        RECT 3135.320 4480.640 3140.040 4481.760 ;
        RECT 3053.280 4477.920 3056.000 4479.040 ;
        RECT 3129.320 4477.920 3134.040 4479.040 ;
        RECT 3082.080 4475.200 3084.800 4476.320 ;
        RECT 3123.320 4475.200 3128.040 4476.320 ;
        RECT 3077.280 4472.480 3080.000 4473.600 ;
        RECT 3117.320 4472.480 3122.040 4473.600 ;
        RECT 3072.480 4469.760 3075.200 4470.880 ;
        RECT 3111.320 4469.760 3116.040 4470.880 ;
        RECT 3067.680 4467.040 3070.400 4468.160 ;
        RECT 3105.320 4467.040 3110.040 4468.160 ;
        RECT 3062.880 4464.320 3065.600 4465.440 ;
        RECT 3099.320 4464.320 3104.040 4465.440 ;
        RECT 3058.080 4461.600 3060.800 4462.720 ;
        RECT 3093.320 4461.600 3098.040 4462.720 ;
        RECT 23.060 4456.160 27.780 4457.280 ;
        RECT 111.900 4456.160 114.620 4457.280 ;
        RECT 29.060 4453.440 33.780 4454.560 ;
        RECT 107.100 4453.440 109.820 4454.560 ;
        RECT 35.060 4450.720 39.780 4451.840 ;
        RECT 78.300 4450.720 81.020 4451.840 ;
        RECT 41.060 4448.000 45.780 4449.120 ;
        RECT 83.100 4448.000 85.820 4449.120 ;
        RECT 47.060 4445.280 51.780 4446.400 ;
        RECT 87.900 4445.280 90.620 4446.400 ;
        RECT 53.060 4442.560 57.780 4443.680 ;
        RECT 92.700 4442.560 95.420 4443.680 ;
        RECT 59.060 4439.840 63.780 4440.960 ;
        RECT 97.500 4439.840 100.220 4440.960 ;
        RECT 65.060 4437.120 69.780 4438.240 ;
        RECT 102.300 4437.120 105.020 4438.240 ;
        RECT 3048.480 4423.520 3051.200 4424.640 ;
        RECT 3135.320 4423.520 3140.040 4424.640 ;
        RECT 3053.280 4420.800 3056.000 4421.920 ;
        RECT 3129.320 4420.800 3134.040 4421.920 ;
        RECT 3082.080 4418.080 3084.800 4419.200 ;
        RECT 3123.320 4418.080 3128.040 4419.200 ;
        RECT 3077.280 4415.360 3080.000 4416.480 ;
        RECT 3117.320 4415.360 3122.040 4416.480 ;
        RECT 3072.480 4412.640 3075.200 4413.760 ;
        RECT 3111.320 4412.640 3116.040 4413.760 ;
        RECT 3067.680 4409.920 3070.400 4411.040 ;
        RECT 3105.320 4409.920 3110.040 4411.040 ;
        RECT 3062.880 4407.200 3065.600 4408.320 ;
        RECT 3099.320 4407.200 3104.040 4408.320 ;
        RECT 3058.080 4404.480 3060.800 4405.600 ;
        RECT 3093.320 4404.480 3098.040 4405.600 ;
        RECT 23.060 4390.880 27.780 4392.000 ;
        RECT 111.900 4390.880 114.620 4392.000 ;
        RECT 29.060 4388.160 33.780 4389.280 ;
        RECT 107.100 4388.160 109.820 4389.280 ;
        RECT 35.060 4385.440 39.780 4386.560 ;
        RECT 78.300 4385.440 81.020 4386.560 ;
        RECT 41.060 4382.720 45.780 4383.840 ;
        RECT 83.100 4382.720 85.820 4383.840 ;
        RECT 47.060 4380.000 51.780 4381.120 ;
        RECT 87.900 4380.000 90.620 4381.120 ;
        RECT 53.060 4377.280 57.780 4378.400 ;
        RECT 92.700 4377.280 95.420 4378.400 ;
        RECT 59.060 4374.560 63.780 4375.680 ;
        RECT 97.500 4374.560 100.220 4375.680 ;
        RECT 65.060 4371.840 69.780 4372.960 ;
        RECT 102.300 4371.840 105.020 4372.960 ;
        RECT 3048.480 4358.240 3051.200 4359.360 ;
        RECT 3135.320 4358.240 3140.040 4359.360 ;
        RECT 3053.280 4355.520 3056.000 4356.640 ;
        RECT 3129.320 4355.520 3134.040 4356.640 ;
        RECT 3082.080 4352.800 3084.800 4353.920 ;
        RECT 3123.320 4352.800 3128.040 4353.920 ;
        RECT 3077.280 4350.080 3080.000 4351.200 ;
        RECT 3117.320 4350.080 3122.040 4351.200 ;
        RECT 3072.480 4347.360 3075.200 4348.480 ;
        RECT 3111.320 4347.360 3116.040 4348.480 ;
        RECT 3067.680 4344.640 3070.400 4345.760 ;
        RECT 3105.320 4344.640 3110.040 4345.760 ;
        RECT 3062.880 4341.920 3065.600 4343.040 ;
        RECT 3099.320 4341.920 3104.040 4343.040 ;
        RECT 3058.080 4339.200 3060.800 4340.320 ;
        RECT 3093.320 4339.200 3098.040 4340.320 ;
        RECT 23.060 4325.600 27.780 4326.720 ;
        RECT 111.900 4325.600 114.620 4326.720 ;
        RECT 29.060 4322.880 33.780 4324.000 ;
        RECT 107.100 4322.880 109.820 4324.000 ;
        RECT 35.060 4320.160 39.780 4321.280 ;
        RECT 78.300 4320.160 81.020 4321.280 ;
        RECT 41.060 4317.440 45.780 4318.560 ;
        RECT 83.100 4317.440 85.820 4318.560 ;
        RECT 47.060 4314.720 51.780 4315.840 ;
        RECT 87.900 4314.720 90.620 4315.840 ;
        RECT 53.060 4312.000 57.780 4313.120 ;
        RECT 92.700 4312.000 95.420 4313.120 ;
        RECT 59.060 4309.280 63.780 4310.400 ;
        RECT 97.500 4309.280 100.220 4310.400 ;
        RECT 65.060 4306.560 69.780 4307.680 ;
        RECT 102.300 4306.560 105.020 4307.680 ;
        RECT 3048.480 4292.960 3051.200 4294.080 ;
        RECT 3135.320 4292.960 3140.040 4294.080 ;
        RECT 3053.280 4290.240 3056.000 4291.360 ;
        RECT 3129.320 4290.240 3134.040 4291.360 ;
        RECT 3082.080 4287.520 3084.800 4288.640 ;
        RECT 3123.320 4287.520 3128.040 4288.640 ;
        RECT 3077.280 4284.800 3080.000 4285.920 ;
        RECT 3117.320 4284.800 3122.040 4285.920 ;
        RECT 3072.480 4282.080 3075.200 4283.200 ;
        RECT 3111.320 4282.080 3116.040 4283.200 ;
        RECT 3067.680 4279.360 3070.400 4280.480 ;
        RECT 3105.320 4279.360 3110.040 4280.480 ;
        RECT 3062.880 4276.640 3065.600 4277.760 ;
        RECT 3099.320 4276.640 3104.040 4277.760 ;
        RECT 3058.080 4273.920 3060.800 4275.040 ;
        RECT 3093.320 4273.920 3098.040 4275.040 ;
        RECT 23.060 4260.320 27.780 4261.440 ;
        RECT 111.900 4260.320 114.620 4261.440 ;
        RECT 29.060 4257.600 33.780 4258.720 ;
        RECT 107.100 4257.600 109.820 4258.720 ;
        RECT 35.060 4254.880 39.780 4256.000 ;
        RECT 78.300 4254.880 81.020 4256.000 ;
        RECT 41.060 4252.160 45.780 4253.280 ;
        RECT 83.100 4252.160 85.820 4253.280 ;
        RECT 47.060 4249.440 51.780 4250.560 ;
        RECT 87.900 4249.440 90.620 4250.560 ;
        RECT 53.060 4246.720 57.780 4247.840 ;
        RECT 92.700 4246.720 95.420 4247.840 ;
        RECT 59.060 4244.000 63.780 4245.120 ;
        RECT 97.500 4244.000 100.220 4245.120 ;
        RECT 65.060 4241.280 69.780 4242.400 ;
        RECT 102.300 4241.280 105.020 4242.400 ;
        RECT 3048.480 4227.680 3051.200 4228.800 ;
        RECT 3135.320 4227.680 3140.040 4228.800 ;
        RECT 3053.280 4224.960 3056.000 4226.080 ;
        RECT 3129.320 4224.960 3134.040 4226.080 ;
        RECT 3082.080 4222.240 3084.800 4223.360 ;
        RECT 3123.320 4222.240 3128.040 4223.360 ;
        RECT 3077.280 4219.520 3080.000 4220.640 ;
        RECT 3117.320 4219.520 3122.040 4220.640 ;
        RECT 3072.480 4216.800 3075.200 4217.920 ;
        RECT 3111.320 4216.800 3116.040 4217.920 ;
        RECT 3067.680 4214.080 3070.400 4215.200 ;
        RECT 3105.320 4214.080 3110.040 4215.200 ;
        RECT 3062.880 4211.360 3065.600 4212.480 ;
        RECT 3099.320 4211.360 3104.040 4212.480 ;
        RECT 3058.080 4208.640 3060.800 4209.760 ;
        RECT 3093.320 4208.640 3098.040 4209.760 ;
        RECT 23.060 4195.040 27.780 4196.160 ;
        RECT 111.900 4195.040 114.620 4196.160 ;
        RECT 29.060 4192.320 33.780 4193.440 ;
        RECT 107.100 4192.320 109.820 4193.440 ;
        RECT 35.060 4189.600 39.780 4190.720 ;
        RECT 78.300 4189.600 81.020 4190.720 ;
        RECT 41.060 4186.880 45.780 4188.000 ;
        RECT 83.100 4186.880 85.820 4188.000 ;
        RECT 47.060 4184.160 51.780 4185.280 ;
        RECT 87.900 4184.160 90.620 4185.280 ;
        RECT 53.060 4181.440 57.780 4182.560 ;
        RECT 92.700 4181.440 95.420 4182.560 ;
        RECT 59.060 4178.720 63.780 4179.840 ;
        RECT 97.500 4178.720 100.220 4179.840 ;
        RECT 65.060 4176.000 69.780 4177.120 ;
        RECT 102.300 4176.000 105.020 4177.120 ;
        RECT 3048.480 4162.400 3051.200 4163.520 ;
        RECT 3135.320 4162.400 3140.040 4163.520 ;
        RECT 3053.280 4159.680 3056.000 4160.800 ;
        RECT 3129.320 4159.680 3134.040 4160.800 ;
        RECT 3082.080 4156.960 3084.800 4158.080 ;
        RECT 3123.320 4156.960 3128.040 4158.080 ;
        RECT 3077.280 4154.240 3080.000 4155.360 ;
        RECT 3117.320 4154.240 3122.040 4155.360 ;
        RECT 3072.480 4151.520 3075.200 4152.640 ;
        RECT 3111.320 4151.520 3116.040 4152.640 ;
        RECT 3067.680 4148.800 3070.400 4149.920 ;
        RECT 3105.320 4148.800 3110.040 4149.920 ;
        RECT 3062.880 4146.080 3065.600 4147.200 ;
        RECT 3099.320 4146.080 3104.040 4147.200 ;
        RECT 3058.080 4143.360 3060.800 4144.480 ;
        RECT 3093.320 4143.360 3098.040 4144.480 ;
        RECT 23.060 4129.760 27.780 4130.880 ;
        RECT 111.900 4129.760 114.620 4130.880 ;
        RECT 29.060 4127.040 33.780 4128.160 ;
        RECT 107.100 4127.040 109.820 4128.160 ;
        RECT 35.060 4124.320 39.780 4125.440 ;
        RECT 78.300 4124.320 81.020 4125.440 ;
        RECT 41.060 4121.600 45.780 4122.720 ;
        RECT 83.100 4121.600 85.820 4122.720 ;
        RECT 47.060 4118.880 51.780 4120.000 ;
        RECT 87.900 4118.880 90.620 4120.000 ;
        RECT 53.060 4116.160 57.780 4117.280 ;
        RECT 92.700 4116.160 95.420 4117.280 ;
        RECT 59.060 4113.440 63.780 4114.560 ;
        RECT 97.500 4113.440 100.220 4114.560 ;
        RECT 65.060 4110.720 69.780 4111.840 ;
        RECT 102.300 4110.720 105.020 4111.840 ;
        RECT 3048.480 4097.120 3051.200 4098.240 ;
        RECT 3135.320 4097.120 3140.040 4098.240 ;
        RECT 3053.280 4094.400 3056.000 4095.520 ;
        RECT 3129.320 4094.400 3134.040 4095.520 ;
        RECT 3082.080 4091.680 3084.800 4092.800 ;
        RECT 3123.320 4091.680 3128.040 4092.800 ;
        RECT 3077.280 4088.960 3080.000 4090.080 ;
        RECT 3117.320 4088.960 3122.040 4090.080 ;
        RECT 3072.480 4086.240 3075.200 4087.360 ;
        RECT 3111.320 4086.240 3116.040 4087.360 ;
        RECT 3067.680 4083.520 3070.400 4084.640 ;
        RECT 3105.320 4083.520 3110.040 4084.640 ;
        RECT 3062.880 4080.800 3065.600 4081.920 ;
        RECT 3099.320 4080.800 3104.040 4081.920 ;
        RECT 3058.080 4078.080 3060.800 4079.200 ;
        RECT 3093.320 4078.080 3098.040 4079.200 ;
        RECT 23.060 4064.480 27.780 4065.600 ;
        RECT 111.900 4064.480 114.620 4065.600 ;
        RECT 29.060 4061.760 33.780 4062.880 ;
        RECT 107.100 4061.760 109.820 4062.880 ;
        RECT 35.060 4059.040 39.780 4060.160 ;
        RECT 78.300 4059.040 81.020 4060.160 ;
        RECT 41.060 4056.320 45.780 4057.440 ;
        RECT 83.100 4056.320 85.820 4057.440 ;
        RECT 47.060 4053.600 51.780 4054.720 ;
        RECT 87.900 4053.600 90.620 4054.720 ;
        RECT 53.060 4050.880 57.780 4052.000 ;
        RECT 92.700 4050.880 95.420 4052.000 ;
        RECT 59.060 4048.160 63.780 4049.280 ;
        RECT 97.500 4048.160 100.220 4049.280 ;
        RECT 65.060 4045.440 69.780 4046.560 ;
        RECT 102.300 4045.440 105.020 4046.560 ;
        RECT 3048.480 4031.840 3051.200 4032.960 ;
        RECT 3135.320 4031.840 3140.040 4032.960 ;
        RECT 3053.280 4029.120 3056.000 4030.240 ;
        RECT 3129.320 4029.120 3134.040 4030.240 ;
        RECT 3082.080 4026.400 3084.800 4027.520 ;
        RECT 3123.320 4026.400 3128.040 4027.520 ;
        RECT 3077.280 4023.680 3080.000 4024.800 ;
        RECT 3117.320 4023.680 3122.040 4024.800 ;
        RECT 3072.480 4020.960 3075.200 4022.080 ;
        RECT 3111.320 4020.960 3116.040 4022.080 ;
        RECT 3067.680 4018.240 3070.400 4019.360 ;
        RECT 3105.320 4018.240 3110.040 4019.360 ;
        RECT 3062.880 4015.520 3065.600 4016.640 ;
        RECT 3099.320 4015.520 3104.040 4016.640 ;
        RECT 3058.080 4012.800 3060.800 4013.920 ;
        RECT 3093.320 4012.800 3098.040 4013.920 ;
        RECT 23.060 3999.200 27.780 4000.320 ;
        RECT 111.900 3999.200 114.620 4000.320 ;
        RECT 29.060 3996.480 33.780 3997.600 ;
        RECT 107.100 3996.480 109.820 3997.600 ;
        RECT 35.060 3993.760 39.780 3994.880 ;
        RECT 78.300 3993.760 81.020 3994.880 ;
        RECT 41.060 3991.040 45.780 3992.160 ;
        RECT 83.100 3991.040 85.820 3992.160 ;
        RECT 47.060 3988.320 51.780 3989.440 ;
        RECT 87.900 3988.320 90.620 3989.440 ;
        RECT 53.060 3985.600 57.780 3986.720 ;
        RECT 92.700 3985.600 95.420 3986.720 ;
        RECT 59.060 3982.880 63.780 3984.000 ;
        RECT 97.500 3982.880 100.220 3984.000 ;
        RECT 65.060 3980.160 69.780 3981.280 ;
        RECT 102.300 3980.160 105.020 3981.280 ;
        RECT 3048.480 3966.560 3051.200 3967.680 ;
        RECT 3135.320 3966.560 3140.040 3967.680 ;
        RECT 3053.280 3963.840 3056.000 3964.960 ;
        RECT 3129.320 3963.840 3134.040 3964.960 ;
        RECT 3082.080 3961.120 3084.800 3962.240 ;
        RECT 3123.320 3961.120 3128.040 3962.240 ;
        RECT 3077.280 3958.400 3080.000 3959.520 ;
        RECT 3117.320 3958.400 3122.040 3959.520 ;
        RECT 3072.480 3955.680 3075.200 3956.800 ;
        RECT 3111.320 3955.680 3116.040 3956.800 ;
        RECT 3067.680 3952.960 3070.400 3954.080 ;
        RECT 3105.320 3952.960 3110.040 3954.080 ;
        RECT 3062.880 3950.240 3065.600 3951.360 ;
        RECT 3099.320 3950.240 3104.040 3951.360 ;
        RECT 3058.080 3947.520 3060.800 3948.640 ;
        RECT 3093.320 3947.520 3098.040 3948.640 ;
        RECT 23.060 3933.920 27.780 3935.040 ;
        RECT 111.900 3933.920 114.620 3935.040 ;
        RECT 29.060 3931.200 33.780 3932.320 ;
        RECT 107.100 3931.200 109.820 3932.320 ;
        RECT 35.060 3928.480 39.780 3929.600 ;
        RECT 78.300 3928.480 81.020 3929.600 ;
        RECT 41.060 3925.760 45.780 3926.880 ;
        RECT 83.100 3925.760 85.820 3926.880 ;
        RECT 47.060 3923.040 51.780 3924.160 ;
        RECT 87.900 3923.040 90.620 3924.160 ;
        RECT 53.060 3920.320 57.780 3921.440 ;
        RECT 92.700 3920.320 95.420 3921.440 ;
        RECT 59.060 3917.600 63.780 3918.720 ;
        RECT 97.500 3917.600 100.220 3918.720 ;
        RECT 65.060 3914.880 69.780 3916.000 ;
        RECT 102.300 3914.880 105.020 3916.000 ;
        RECT 3048.480 3901.280 3051.200 3902.400 ;
        RECT 3135.320 3901.280 3140.040 3902.400 ;
        RECT 3053.280 3898.560 3056.000 3899.680 ;
        RECT 3129.320 3898.560 3134.040 3899.680 ;
        RECT 3082.080 3895.840 3084.800 3896.960 ;
        RECT 3123.320 3895.840 3128.040 3896.960 ;
        RECT 3077.280 3893.120 3080.000 3894.240 ;
        RECT 3117.320 3893.120 3122.040 3894.240 ;
        RECT 3072.480 3890.400 3075.200 3891.520 ;
        RECT 3111.320 3890.400 3116.040 3891.520 ;
        RECT 3067.680 3887.680 3070.400 3888.800 ;
        RECT 3105.320 3887.680 3110.040 3888.800 ;
        RECT 3062.880 3884.960 3065.600 3886.080 ;
        RECT 3099.320 3884.960 3104.040 3886.080 ;
        RECT 3058.080 3882.240 3060.800 3883.360 ;
        RECT 3093.320 3882.240 3098.040 3883.360 ;
        RECT 23.060 3868.640 27.780 3869.760 ;
        RECT 111.900 3868.640 114.620 3869.760 ;
        RECT 29.060 3865.920 33.780 3867.040 ;
        RECT 107.100 3865.920 109.820 3867.040 ;
        RECT 35.060 3863.200 39.780 3864.320 ;
        RECT 78.300 3863.200 81.020 3864.320 ;
        RECT 41.060 3860.480 45.780 3861.600 ;
        RECT 83.100 3860.480 85.820 3861.600 ;
        RECT 47.060 3857.760 51.780 3858.880 ;
        RECT 87.900 3857.760 90.620 3858.880 ;
        RECT 53.060 3855.040 57.780 3856.160 ;
        RECT 92.700 3855.040 95.420 3856.160 ;
        RECT 59.060 3852.320 63.780 3853.440 ;
        RECT 97.500 3852.320 100.220 3853.440 ;
        RECT 65.060 3849.600 69.780 3850.720 ;
        RECT 102.300 3849.600 105.020 3850.720 ;
        RECT 3048.480 3836.000 3051.200 3837.120 ;
        RECT 3135.320 3836.000 3140.040 3837.120 ;
        RECT 3053.280 3833.280 3056.000 3834.400 ;
        RECT 3129.320 3833.280 3134.040 3834.400 ;
        RECT 3082.080 3830.560 3084.800 3831.680 ;
        RECT 3123.320 3830.560 3128.040 3831.680 ;
        RECT 3077.280 3827.840 3080.000 3828.960 ;
        RECT 3117.320 3827.840 3122.040 3828.960 ;
        RECT 3072.480 3825.120 3075.200 3826.240 ;
        RECT 3111.320 3825.120 3116.040 3826.240 ;
        RECT 3067.680 3822.400 3070.400 3823.520 ;
        RECT 3105.320 3822.400 3110.040 3823.520 ;
        RECT 3062.880 3819.680 3065.600 3820.800 ;
        RECT 3099.320 3819.680 3104.040 3820.800 ;
        RECT 3058.080 3816.960 3060.800 3818.080 ;
        RECT 3093.320 3816.960 3098.040 3818.080 ;
        RECT 23.060 3803.360 27.780 3804.480 ;
        RECT 111.900 3803.360 114.620 3804.480 ;
        RECT 29.060 3800.640 33.780 3801.760 ;
        RECT 107.100 3800.640 109.820 3801.760 ;
        RECT 35.060 3797.920 39.780 3799.040 ;
        RECT 78.300 3797.920 81.020 3799.040 ;
        RECT 41.060 3795.200 45.780 3796.320 ;
        RECT 83.100 3795.200 85.820 3796.320 ;
        RECT 47.060 3792.480 51.780 3793.600 ;
        RECT 87.900 3792.480 90.620 3793.600 ;
        RECT 53.060 3789.760 57.780 3790.880 ;
        RECT 92.700 3789.760 95.420 3790.880 ;
        RECT 59.060 3787.040 63.780 3788.160 ;
        RECT 97.500 3787.040 100.220 3788.160 ;
        RECT 65.060 3784.320 69.780 3785.440 ;
        RECT 102.300 3784.320 105.020 3785.440 ;
        RECT 3048.480 3770.720 3051.200 3771.840 ;
        RECT 3135.320 3770.720 3140.040 3771.840 ;
        RECT 3053.280 3768.000 3056.000 3769.120 ;
        RECT 3129.320 3768.000 3134.040 3769.120 ;
        RECT 3082.080 3765.280 3084.800 3766.400 ;
        RECT 3123.320 3765.280 3128.040 3766.400 ;
        RECT 3077.280 3762.560 3080.000 3763.680 ;
        RECT 3117.320 3762.560 3122.040 3763.680 ;
        RECT 3072.480 3759.840 3075.200 3760.960 ;
        RECT 3111.320 3759.840 3116.040 3760.960 ;
        RECT 3067.680 3757.120 3070.400 3758.240 ;
        RECT 3105.320 3757.120 3110.040 3758.240 ;
        RECT 3062.880 3754.400 3065.600 3755.520 ;
        RECT 3099.320 3754.400 3104.040 3755.520 ;
        RECT 3058.080 3751.680 3060.800 3752.800 ;
        RECT 3093.320 3751.680 3098.040 3752.800 ;
        RECT 23.060 3738.080 27.780 3739.200 ;
        RECT 111.900 3738.080 114.620 3739.200 ;
        RECT 29.060 3735.360 33.780 3736.480 ;
        RECT 107.100 3735.360 109.820 3736.480 ;
        RECT 35.060 3732.640 39.780 3733.760 ;
        RECT 78.300 3732.640 81.020 3733.760 ;
        RECT 41.060 3729.920 45.780 3731.040 ;
        RECT 83.100 3729.920 85.820 3731.040 ;
        RECT 47.060 3727.200 51.780 3728.320 ;
        RECT 87.900 3727.200 90.620 3728.320 ;
        RECT 53.060 3724.480 57.780 3725.600 ;
        RECT 92.700 3724.480 95.420 3725.600 ;
        RECT 59.060 3721.760 63.780 3722.880 ;
        RECT 97.500 3721.760 100.220 3722.880 ;
        RECT 65.060 3719.040 69.780 3720.160 ;
        RECT 102.300 3719.040 105.020 3720.160 ;
        RECT 3048.480 3705.440 3051.200 3706.560 ;
        RECT 3135.320 3705.440 3140.040 3706.560 ;
        RECT 3053.280 3702.720 3056.000 3703.840 ;
        RECT 3129.320 3702.720 3134.040 3703.840 ;
        RECT 3082.080 3700.000 3084.800 3701.120 ;
        RECT 3123.320 3700.000 3128.040 3701.120 ;
        RECT 3077.280 3697.280 3080.000 3698.400 ;
        RECT 3117.320 3697.280 3122.040 3698.400 ;
        RECT 3072.480 3694.560 3075.200 3695.680 ;
        RECT 3111.320 3694.560 3116.040 3695.680 ;
        RECT 3067.680 3691.840 3070.400 3692.960 ;
        RECT 3105.320 3691.840 3110.040 3692.960 ;
        RECT 3062.880 3689.120 3065.600 3690.240 ;
        RECT 3099.320 3689.120 3104.040 3690.240 ;
        RECT 3058.080 3686.400 3060.800 3687.520 ;
        RECT 3093.320 3686.400 3098.040 3687.520 ;
        RECT 23.060 3680.960 27.780 3682.080 ;
        RECT 111.900 3680.960 114.620 3682.080 ;
        RECT 29.060 3678.240 33.780 3679.360 ;
        RECT 107.100 3678.240 109.820 3679.360 ;
        RECT 35.060 3675.520 39.780 3676.640 ;
        RECT 78.300 3675.520 81.020 3676.640 ;
        RECT 41.060 3672.800 45.780 3673.920 ;
        RECT 83.100 3672.800 85.820 3673.920 ;
        RECT 47.060 3670.080 51.780 3671.200 ;
        RECT 87.900 3670.080 90.620 3671.200 ;
        RECT 53.060 3667.360 57.780 3668.480 ;
        RECT 92.700 3667.360 95.420 3668.480 ;
        RECT 59.060 3664.640 63.780 3665.760 ;
        RECT 97.500 3664.640 100.220 3665.760 ;
        RECT 65.060 3661.920 69.780 3663.040 ;
        RECT 102.300 3661.920 105.020 3663.040 ;
        RECT 3048.480 3640.160 3051.200 3641.280 ;
        RECT 3135.320 3640.160 3140.040 3641.280 ;
        RECT 3053.280 3637.440 3056.000 3638.560 ;
        RECT 3129.320 3637.440 3134.040 3638.560 ;
        RECT 3082.080 3634.720 3084.800 3635.840 ;
        RECT 3123.320 3634.720 3128.040 3635.840 ;
        RECT 3077.280 3632.000 3080.000 3633.120 ;
        RECT 3117.320 3632.000 3122.040 3633.120 ;
        RECT 3072.480 3629.280 3075.200 3630.400 ;
        RECT 3111.320 3629.280 3116.040 3630.400 ;
        RECT 3067.680 3626.560 3070.400 3627.680 ;
        RECT 3105.320 3626.560 3110.040 3627.680 ;
        RECT 3062.880 3623.840 3065.600 3624.960 ;
        RECT 3099.320 3623.840 3104.040 3624.960 ;
        RECT 3058.080 3621.120 3060.800 3622.240 ;
        RECT 3093.320 3621.120 3098.040 3622.240 ;
        RECT 23.060 3607.520 27.780 3608.640 ;
        RECT 111.900 3607.520 114.620 3608.640 ;
        RECT 29.060 3604.800 33.780 3605.920 ;
        RECT 107.100 3604.800 109.820 3605.920 ;
        RECT 35.060 3602.080 39.780 3603.200 ;
        RECT 78.300 3602.080 81.020 3603.200 ;
        RECT 41.060 3599.360 45.780 3600.480 ;
        RECT 83.100 3599.360 85.820 3600.480 ;
        RECT 47.060 3596.640 51.780 3597.760 ;
        RECT 87.900 3596.640 90.620 3597.760 ;
        RECT 53.060 3593.920 57.780 3595.040 ;
        RECT 92.700 3593.920 95.420 3595.040 ;
        RECT 59.060 3591.200 63.780 3592.320 ;
        RECT 97.500 3591.200 100.220 3592.320 ;
        RECT 65.060 3588.480 69.780 3589.600 ;
        RECT 102.300 3588.480 105.020 3589.600 ;
        RECT 3048.480 3566.720 3051.200 3567.840 ;
        RECT 3135.320 3566.720 3140.040 3567.840 ;
        RECT 3053.280 3564.000 3056.000 3565.120 ;
        RECT 3129.320 3564.000 3134.040 3565.120 ;
        RECT 3082.080 3561.280 3084.800 3562.400 ;
        RECT 3123.320 3561.280 3128.040 3562.400 ;
        RECT 3077.280 3558.560 3080.000 3559.680 ;
        RECT 3117.320 3558.560 3122.040 3559.680 ;
        RECT 3072.480 3555.840 3075.200 3556.960 ;
        RECT 3111.320 3555.840 3116.040 3556.960 ;
        RECT 3067.680 3553.120 3070.400 3554.240 ;
        RECT 3105.320 3553.120 3110.040 3554.240 ;
        RECT 3062.880 3550.400 3065.600 3551.520 ;
        RECT 3099.320 3550.400 3104.040 3551.520 ;
        RECT 3058.080 3547.680 3060.800 3548.800 ;
        RECT 3093.320 3547.680 3098.040 3548.800 ;
        RECT 23.060 3542.240 27.780 3543.360 ;
        RECT 111.900 3542.240 114.620 3543.360 ;
        RECT 29.060 3539.520 33.780 3540.640 ;
        RECT 107.100 3539.520 109.820 3540.640 ;
        RECT 35.060 3536.800 39.780 3537.920 ;
        RECT 78.300 3536.800 81.020 3537.920 ;
        RECT 41.060 3534.080 45.780 3535.200 ;
        RECT 83.100 3534.080 85.820 3535.200 ;
        RECT 47.060 3531.360 51.780 3532.480 ;
        RECT 87.900 3531.360 90.620 3532.480 ;
        RECT 53.060 3528.640 57.780 3529.760 ;
        RECT 92.700 3528.640 95.420 3529.760 ;
        RECT 59.060 3525.920 63.780 3527.040 ;
        RECT 97.500 3525.920 100.220 3527.040 ;
        RECT 65.060 3523.200 69.780 3524.320 ;
        RECT 102.300 3523.200 105.020 3524.320 ;
        RECT 3048.480 3509.600 3051.200 3510.720 ;
        RECT 3135.320 3509.600 3140.040 3510.720 ;
        RECT 3053.280 3506.880 3056.000 3508.000 ;
        RECT 3129.320 3506.880 3134.040 3508.000 ;
        RECT 3082.080 3504.160 3084.800 3505.280 ;
        RECT 3123.320 3504.160 3128.040 3505.280 ;
        RECT 3077.280 3501.440 3080.000 3502.560 ;
        RECT 3117.320 3501.440 3122.040 3502.560 ;
        RECT 3072.480 3498.720 3075.200 3499.840 ;
        RECT 3111.320 3498.720 3116.040 3499.840 ;
        RECT 3067.680 3496.000 3070.400 3497.120 ;
        RECT 3105.320 3496.000 3110.040 3497.120 ;
        RECT 3062.880 3493.280 3065.600 3494.400 ;
        RECT 3099.320 3493.280 3104.040 3494.400 ;
        RECT 3058.080 3490.560 3060.800 3491.680 ;
        RECT 3093.320 3490.560 3098.040 3491.680 ;
        RECT 23.060 3460.640 27.780 3461.760 ;
        RECT 111.900 3460.640 114.620 3461.760 ;
        RECT 29.060 3457.920 33.780 3459.040 ;
        RECT 107.100 3457.920 109.820 3459.040 ;
        RECT 35.060 3455.200 39.780 3456.320 ;
        RECT 78.300 3455.200 81.020 3456.320 ;
        RECT 41.060 3452.480 45.780 3453.600 ;
        RECT 83.100 3452.480 85.820 3453.600 ;
        RECT 47.060 3449.760 51.780 3450.880 ;
        RECT 87.900 3449.760 90.620 3450.880 ;
        RECT 53.060 3447.040 57.780 3448.160 ;
        RECT 92.700 3447.040 95.420 3448.160 ;
        RECT 59.060 3444.320 63.780 3445.440 ;
        RECT 97.500 3444.320 100.220 3445.440 ;
        RECT 3048.480 3444.320 3051.200 3445.440 ;
        RECT 3135.320 3444.320 3140.040 3445.440 ;
        RECT 65.060 3441.600 69.780 3442.720 ;
        RECT 102.300 3441.600 105.020 3442.720 ;
        RECT 3053.280 3441.600 3056.000 3442.720 ;
        RECT 3129.320 3441.600 3134.040 3442.720 ;
        RECT 3082.080 3438.880 3084.800 3440.000 ;
        RECT 3123.320 3438.880 3128.040 3440.000 ;
        RECT 3077.280 3436.160 3080.000 3437.280 ;
        RECT 3117.320 3436.160 3122.040 3437.280 ;
        RECT 3072.480 3433.440 3075.200 3434.560 ;
        RECT 3111.320 3433.440 3116.040 3434.560 ;
        RECT 3067.680 3430.720 3070.400 3431.840 ;
        RECT 3105.320 3430.720 3110.040 3431.840 ;
        RECT 3062.880 3428.000 3065.600 3429.120 ;
        RECT 3099.320 3428.000 3104.040 3429.120 ;
        RECT 3058.080 3425.280 3060.800 3426.400 ;
        RECT 3093.320 3425.280 3098.040 3426.400 ;
        RECT 23.060 3411.680 27.780 3412.800 ;
        RECT 111.900 3411.680 114.620 3412.800 ;
        RECT 29.060 3408.960 33.780 3410.080 ;
        RECT 107.100 3408.960 109.820 3410.080 ;
        RECT 35.060 3406.240 39.780 3407.360 ;
        RECT 78.300 3406.240 81.020 3407.360 ;
        RECT 41.060 3403.520 45.780 3404.640 ;
        RECT 83.100 3403.520 85.820 3404.640 ;
        RECT 47.060 3400.800 51.780 3401.920 ;
        RECT 87.900 3400.800 90.620 3401.920 ;
        RECT 53.060 3398.080 57.780 3399.200 ;
        RECT 92.700 3398.080 95.420 3399.200 ;
        RECT 59.060 3395.360 63.780 3396.480 ;
        RECT 97.500 3395.360 100.220 3396.480 ;
        RECT 65.060 3392.640 69.780 3393.760 ;
        RECT 102.300 3392.640 105.020 3393.760 ;
        RECT 3048.480 3379.040 3051.200 3380.160 ;
        RECT 3135.320 3379.040 3140.040 3380.160 ;
        RECT 3053.280 3376.320 3056.000 3377.440 ;
        RECT 3129.320 3376.320 3134.040 3377.440 ;
        RECT 3082.080 3373.600 3084.800 3374.720 ;
        RECT 3123.320 3373.600 3128.040 3374.720 ;
        RECT 3077.280 3370.880 3080.000 3372.000 ;
        RECT 3117.320 3370.880 3122.040 3372.000 ;
        RECT 3072.480 3368.160 3075.200 3369.280 ;
        RECT 3111.320 3368.160 3116.040 3369.280 ;
        RECT 3067.680 3365.440 3070.400 3366.560 ;
        RECT 3105.320 3365.440 3110.040 3366.560 ;
        RECT 3062.880 3362.720 3065.600 3363.840 ;
        RECT 3099.320 3362.720 3104.040 3363.840 ;
        RECT 3058.080 3360.000 3060.800 3361.120 ;
        RECT 3093.320 3360.000 3098.040 3361.120 ;
        RECT 23.060 3346.400 27.780 3347.520 ;
        RECT 111.900 3346.400 114.620 3347.520 ;
        RECT 29.060 3343.680 33.780 3344.800 ;
        RECT 107.100 3343.680 109.820 3344.800 ;
        RECT 35.060 3340.960 39.780 3342.080 ;
        RECT 78.300 3340.960 81.020 3342.080 ;
        RECT 41.060 3338.240 45.780 3339.360 ;
        RECT 83.100 3338.240 85.820 3339.360 ;
        RECT 47.060 3335.520 51.780 3336.640 ;
        RECT 87.900 3335.520 90.620 3336.640 ;
        RECT 53.060 3332.800 57.780 3333.920 ;
        RECT 92.700 3332.800 95.420 3333.920 ;
        RECT 59.060 3330.080 63.780 3331.200 ;
        RECT 97.500 3330.080 100.220 3331.200 ;
        RECT 65.060 3327.360 69.780 3328.480 ;
        RECT 102.300 3327.360 105.020 3328.480 ;
        RECT 3048.480 3313.760 3051.200 3314.880 ;
        RECT 3135.320 3313.760 3140.040 3314.880 ;
        RECT 3053.280 3311.040 3056.000 3312.160 ;
        RECT 3129.320 3311.040 3134.040 3312.160 ;
        RECT 3082.080 3308.320 3084.800 3309.440 ;
        RECT 3123.320 3308.320 3128.040 3309.440 ;
        RECT 3077.280 3305.600 3080.000 3306.720 ;
        RECT 3117.320 3305.600 3122.040 3306.720 ;
        RECT 3072.480 3302.880 3075.200 3304.000 ;
        RECT 3111.320 3302.880 3116.040 3304.000 ;
        RECT 3067.680 3300.160 3070.400 3301.280 ;
        RECT 3105.320 3300.160 3110.040 3301.280 ;
        RECT 3062.880 3297.440 3065.600 3298.560 ;
        RECT 3099.320 3297.440 3104.040 3298.560 ;
        RECT 3058.080 3294.720 3060.800 3295.840 ;
        RECT 3093.320 3294.720 3098.040 3295.840 ;
        RECT 23.060 3281.120 27.780 3282.240 ;
        RECT 111.900 3281.120 114.620 3282.240 ;
        RECT 29.060 3278.400 33.780 3279.520 ;
        RECT 107.100 3278.400 109.820 3279.520 ;
        RECT 35.060 3275.680 39.780 3276.800 ;
        RECT 78.300 3275.680 81.020 3276.800 ;
        RECT 41.060 3272.960 45.780 3274.080 ;
        RECT 83.100 3272.960 85.820 3274.080 ;
        RECT 47.060 3270.240 51.780 3271.360 ;
        RECT 87.900 3270.240 90.620 3271.360 ;
        RECT 53.060 3267.520 57.780 3268.640 ;
        RECT 92.700 3267.520 95.420 3268.640 ;
        RECT 59.060 3264.800 63.780 3265.920 ;
        RECT 97.500 3264.800 100.220 3265.920 ;
        RECT 65.060 3262.080 69.780 3263.200 ;
        RECT 102.300 3262.080 105.020 3263.200 ;
        RECT 3048.480 3248.480 3051.200 3249.600 ;
        RECT 3135.320 3248.480 3140.040 3249.600 ;
        RECT 3053.280 3245.760 3056.000 3246.880 ;
        RECT 3129.320 3245.760 3134.040 3246.880 ;
        RECT 3082.080 3243.040 3084.800 3244.160 ;
        RECT 3123.320 3243.040 3128.040 3244.160 ;
        RECT 3077.280 3240.320 3080.000 3241.440 ;
        RECT 3117.320 3240.320 3122.040 3241.440 ;
        RECT 3072.480 3237.600 3075.200 3238.720 ;
        RECT 3111.320 3237.600 3116.040 3238.720 ;
        RECT 3067.680 3234.880 3070.400 3236.000 ;
        RECT 3105.320 3234.880 3110.040 3236.000 ;
        RECT 3062.880 3232.160 3065.600 3233.280 ;
        RECT 3099.320 3232.160 3104.040 3233.280 ;
        RECT 3058.080 3229.440 3060.800 3230.560 ;
        RECT 3093.320 3229.440 3098.040 3230.560 ;
        RECT 23.060 3207.680 27.780 3208.800 ;
        RECT 111.900 3207.680 114.620 3208.800 ;
        RECT 29.060 3204.960 33.780 3206.080 ;
        RECT 107.100 3204.960 109.820 3206.080 ;
        RECT 35.060 3202.240 39.780 3203.360 ;
        RECT 78.300 3202.240 81.020 3203.360 ;
        RECT 41.060 3199.520 45.780 3200.640 ;
        RECT 83.100 3199.520 85.820 3200.640 ;
        RECT 47.060 3196.800 51.780 3197.920 ;
        RECT 87.900 3196.800 90.620 3197.920 ;
        RECT 53.060 3194.080 57.780 3195.200 ;
        RECT 92.700 3194.080 95.420 3195.200 ;
        RECT 59.060 3191.360 63.780 3192.480 ;
        RECT 97.500 3191.360 100.220 3192.480 ;
        RECT 65.060 3188.640 69.780 3189.760 ;
        RECT 102.300 3188.640 105.020 3189.760 ;
        RECT 3048.480 3183.200 3051.200 3184.320 ;
        RECT 3135.320 3183.200 3140.040 3184.320 ;
        RECT 3053.280 3180.480 3056.000 3181.600 ;
        RECT 3129.320 3180.480 3134.040 3181.600 ;
        RECT 3082.080 3177.760 3084.800 3178.880 ;
        RECT 3123.320 3177.760 3128.040 3178.880 ;
        RECT 3077.280 3175.040 3080.000 3176.160 ;
        RECT 3117.320 3175.040 3122.040 3176.160 ;
        RECT 3072.480 3172.320 3075.200 3173.440 ;
        RECT 3111.320 3172.320 3116.040 3173.440 ;
        RECT 3067.680 3169.600 3070.400 3170.720 ;
        RECT 3105.320 3169.600 3110.040 3170.720 ;
        RECT 3062.880 3166.880 3065.600 3168.000 ;
        RECT 3099.320 3166.880 3104.040 3168.000 ;
        RECT 3058.080 3164.160 3060.800 3165.280 ;
        RECT 3093.320 3164.160 3098.040 3165.280 ;
        RECT 23.060 3150.560 27.780 3151.680 ;
        RECT 111.900 3150.560 114.620 3151.680 ;
        RECT 29.060 3147.840 33.780 3148.960 ;
        RECT 107.100 3147.840 109.820 3148.960 ;
        RECT 35.060 3145.120 39.780 3146.240 ;
        RECT 78.300 3145.120 81.020 3146.240 ;
        RECT 41.060 3142.400 45.780 3143.520 ;
        RECT 83.100 3142.400 85.820 3143.520 ;
        RECT 47.060 3139.680 51.780 3140.800 ;
        RECT 87.900 3139.680 90.620 3140.800 ;
        RECT 53.060 3136.960 57.780 3138.080 ;
        RECT 92.700 3136.960 95.420 3138.080 ;
        RECT 59.060 3134.240 63.780 3135.360 ;
        RECT 97.500 3134.240 100.220 3135.360 ;
        RECT 65.060 3131.520 69.780 3132.640 ;
        RECT 102.300 3131.520 105.020 3132.640 ;
        RECT 3048.480 3117.920 3051.200 3119.040 ;
        RECT 3135.320 3117.920 3140.040 3119.040 ;
        RECT 3053.280 3115.200 3056.000 3116.320 ;
        RECT 3129.320 3115.200 3134.040 3116.320 ;
        RECT 3082.080 3112.480 3084.800 3113.600 ;
        RECT 3123.320 3112.480 3128.040 3113.600 ;
        RECT 3077.280 3109.760 3080.000 3110.880 ;
        RECT 3117.320 3109.760 3122.040 3110.880 ;
        RECT 3072.480 3107.040 3075.200 3108.160 ;
        RECT 3111.320 3107.040 3116.040 3108.160 ;
        RECT 3067.680 3104.320 3070.400 3105.440 ;
        RECT 3105.320 3104.320 3110.040 3105.440 ;
        RECT 3062.880 3101.600 3065.600 3102.720 ;
        RECT 3099.320 3101.600 3104.040 3102.720 ;
        RECT 3058.080 3098.880 3060.800 3100.000 ;
        RECT 3093.320 3098.880 3098.040 3100.000 ;
        RECT 23.060 3085.280 27.780 3086.400 ;
        RECT 111.900 3085.280 114.620 3086.400 ;
        RECT 29.060 3082.560 33.780 3083.680 ;
        RECT 107.100 3082.560 109.820 3083.680 ;
        RECT 35.060 3079.840 39.780 3080.960 ;
        RECT 78.300 3079.840 81.020 3080.960 ;
        RECT 41.060 3077.120 45.780 3078.240 ;
        RECT 83.100 3077.120 85.820 3078.240 ;
        RECT 47.060 3074.400 51.780 3075.520 ;
        RECT 87.900 3074.400 90.620 3075.520 ;
        RECT 53.060 3071.680 57.780 3072.800 ;
        RECT 92.700 3071.680 95.420 3072.800 ;
        RECT 59.060 3068.960 63.780 3070.080 ;
        RECT 97.500 3068.960 100.220 3070.080 ;
        RECT 65.060 3066.240 69.780 3067.360 ;
        RECT 102.300 3066.240 105.020 3067.360 ;
        RECT 3048.480 3052.640 3051.200 3053.760 ;
        RECT 3135.320 3052.640 3140.040 3053.760 ;
        RECT 3053.280 3049.920 3056.000 3051.040 ;
        RECT 3129.320 3049.920 3134.040 3051.040 ;
        RECT 3082.080 3047.200 3084.800 3048.320 ;
        RECT 3123.320 3047.200 3128.040 3048.320 ;
        RECT 3077.280 3044.480 3080.000 3045.600 ;
        RECT 3117.320 3044.480 3122.040 3045.600 ;
        RECT 3072.480 3041.760 3075.200 3042.880 ;
        RECT 3111.320 3041.760 3116.040 3042.880 ;
        RECT 3067.680 3039.040 3070.400 3040.160 ;
        RECT 3105.320 3039.040 3110.040 3040.160 ;
        RECT 3062.880 3036.320 3065.600 3037.440 ;
        RECT 3099.320 3036.320 3104.040 3037.440 ;
        RECT 3058.080 3033.600 3060.800 3034.720 ;
        RECT 3093.320 3033.600 3098.040 3034.720 ;
        RECT 23.060 3030.880 27.780 3032.000 ;
        RECT 111.900 3030.880 114.620 3032.000 ;
        RECT 29.060 3028.160 33.780 3029.280 ;
        RECT 107.100 3028.160 109.820 3029.280 ;
        RECT 35.060 3025.440 39.780 3026.560 ;
        RECT 78.300 3025.440 81.020 3026.560 ;
        RECT 41.060 3022.720 45.780 3023.840 ;
        RECT 83.100 3022.720 85.820 3023.840 ;
        RECT 47.060 3020.000 51.780 3021.120 ;
        RECT 87.900 3020.000 90.620 3021.120 ;
        RECT 53.060 3017.280 57.780 3018.400 ;
        RECT 92.700 3017.280 95.420 3018.400 ;
        RECT 59.060 3014.560 63.780 3015.680 ;
        RECT 97.500 3014.560 100.220 3015.680 ;
        RECT 65.060 3011.840 69.780 3012.960 ;
        RECT 102.300 3011.840 105.020 3012.960 ;
        RECT 3048.480 2987.360 3051.200 2988.480 ;
        RECT 3135.320 2987.360 3140.040 2988.480 ;
        RECT 3053.280 2984.640 3056.000 2985.760 ;
        RECT 3129.320 2984.640 3134.040 2985.760 ;
        RECT 3082.080 2981.920 3084.800 2983.040 ;
        RECT 3123.320 2981.920 3128.040 2983.040 ;
        RECT 3077.280 2979.200 3080.000 2980.320 ;
        RECT 3117.320 2979.200 3122.040 2980.320 ;
        RECT 3072.480 2976.480 3075.200 2977.600 ;
        RECT 3111.320 2976.480 3116.040 2977.600 ;
        RECT 3067.680 2973.760 3070.400 2974.880 ;
        RECT 3105.320 2973.760 3110.040 2974.880 ;
        RECT 3062.880 2971.040 3065.600 2972.160 ;
        RECT 3099.320 2971.040 3104.040 2972.160 ;
        RECT 3058.080 2968.320 3060.800 2969.440 ;
        RECT 3093.320 2968.320 3098.040 2969.440 ;
        RECT 23.060 2954.720 27.780 2955.840 ;
        RECT 111.900 2954.720 114.620 2955.840 ;
        RECT 29.060 2952.000 33.780 2953.120 ;
        RECT 107.100 2952.000 109.820 2953.120 ;
        RECT 35.060 2949.280 39.780 2950.400 ;
        RECT 78.300 2949.280 81.020 2950.400 ;
        RECT 41.060 2946.560 45.780 2947.680 ;
        RECT 83.100 2946.560 85.820 2947.680 ;
        RECT 47.060 2943.840 51.780 2944.960 ;
        RECT 87.900 2943.840 90.620 2944.960 ;
        RECT 53.060 2941.120 57.780 2942.240 ;
        RECT 92.700 2941.120 95.420 2942.240 ;
        RECT 59.060 2938.400 63.780 2939.520 ;
        RECT 97.500 2938.400 100.220 2939.520 ;
        RECT 65.060 2935.680 69.780 2936.800 ;
        RECT 102.300 2935.680 105.020 2936.800 ;
        RECT 3048.480 2922.080 3051.200 2923.200 ;
        RECT 3135.320 2922.080 3140.040 2923.200 ;
        RECT 3053.280 2919.360 3056.000 2920.480 ;
        RECT 3129.320 2919.360 3134.040 2920.480 ;
        RECT 3082.080 2916.640 3084.800 2917.760 ;
        RECT 3123.320 2916.640 3128.040 2917.760 ;
        RECT 3077.280 2913.920 3080.000 2915.040 ;
        RECT 3117.320 2913.920 3122.040 2915.040 ;
        RECT 3072.480 2911.200 3075.200 2912.320 ;
        RECT 3111.320 2911.200 3116.040 2912.320 ;
        RECT 3067.680 2908.480 3070.400 2909.600 ;
        RECT 3105.320 2908.480 3110.040 2909.600 ;
        RECT 3062.880 2905.760 3065.600 2906.880 ;
        RECT 3099.320 2905.760 3104.040 2906.880 ;
        RECT 3058.080 2903.040 3060.800 2904.160 ;
        RECT 3093.320 2903.040 3098.040 2904.160 ;
        RECT 23.060 2889.440 27.780 2890.560 ;
        RECT 111.900 2889.440 114.620 2890.560 ;
        RECT 29.060 2886.720 33.780 2887.840 ;
        RECT 107.100 2886.720 109.820 2887.840 ;
        RECT 35.060 2884.000 39.780 2885.120 ;
        RECT 78.300 2884.000 81.020 2885.120 ;
        RECT 41.060 2881.280 45.780 2882.400 ;
        RECT 83.100 2881.280 85.820 2882.400 ;
        RECT 47.060 2878.560 51.780 2879.680 ;
        RECT 87.900 2878.560 90.620 2879.680 ;
        RECT 53.060 2875.840 57.780 2876.960 ;
        RECT 92.700 2875.840 95.420 2876.960 ;
        RECT 59.060 2873.120 63.780 2874.240 ;
        RECT 97.500 2873.120 100.220 2874.240 ;
        RECT 65.060 2870.400 69.780 2871.520 ;
        RECT 102.300 2870.400 105.020 2871.520 ;
        RECT 3048.480 2856.800 3051.200 2857.920 ;
        RECT 3135.320 2856.800 3140.040 2857.920 ;
        RECT 3053.280 2854.080 3056.000 2855.200 ;
        RECT 3129.320 2854.080 3134.040 2855.200 ;
        RECT 3082.080 2851.360 3084.800 2852.480 ;
        RECT 3123.320 2851.360 3128.040 2852.480 ;
        RECT 3077.280 2848.640 3080.000 2849.760 ;
        RECT 3117.320 2848.640 3122.040 2849.760 ;
        RECT 3072.480 2845.920 3075.200 2847.040 ;
        RECT 3111.320 2845.920 3116.040 2847.040 ;
        RECT 3067.680 2843.200 3070.400 2844.320 ;
        RECT 3105.320 2843.200 3110.040 2844.320 ;
        RECT 3062.880 2840.480 3065.600 2841.600 ;
        RECT 3099.320 2840.480 3104.040 2841.600 ;
        RECT 3058.080 2837.760 3060.800 2838.880 ;
        RECT 3093.320 2837.760 3098.040 2838.880 ;
        RECT 23.060 2835.040 27.780 2836.160 ;
        RECT 111.900 2835.040 114.620 2836.160 ;
        RECT 29.060 2832.320 33.780 2833.440 ;
        RECT 107.100 2832.320 109.820 2833.440 ;
        RECT 35.060 2829.600 39.780 2830.720 ;
        RECT 78.300 2829.600 81.020 2830.720 ;
        RECT 41.060 2826.880 45.780 2828.000 ;
        RECT 83.100 2826.880 85.820 2828.000 ;
        RECT 47.060 2824.160 51.780 2825.280 ;
        RECT 87.900 2824.160 90.620 2825.280 ;
        RECT 53.060 2821.440 57.780 2822.560 ;
        RECT 92.700 2821.440 95.420 2822.560 ;
        RECT 59.060 2818.720 63.780 2819.840 ;
        RECT 97.500 2818.720 100.220 2819.840 ;
        RECT 65.060 2816.000 69.780 2817.120 ;
        RECT 102.300 2816.000 105.020 2817.120 ;
        RECT 3048.480 2791.520 3051.200 2792.640 ;
        RECT 3135.320 2791.520 3140.040 2792.640 ;
        RECT 3053.280 2788.800 3056.000 2789.920 ;
        RECT 3129.320 2788.800 3134.040 2789.920 ;
        RECT 3082.080 2786.080 3084.800 2787.200 ;
        RECT 3123.320 2786.080 3128.040 2787.200 ;
        RECT 3077.280 2783.360 3080.000 2784.480 ;
        RECT 3117.320 2783.360 3122.040 2784.480 ;
        RECT 3072.480 2780.640 3075.200 2781.760 ;
        RECT 3111.320 2780.640 3116.040 2781.760 ;
        RECT 3067.680 2777.920 3070.400 2779.040 ;
        RECT 3105.320 2777.920 3110.040 2779.040 ;
        RECT 3062.880 2775.200 3065.600 2776.320 ;
        RECT 3099.320 2775.200 3104.040 2776.320 ;
        RECT 3058.080 2772.480 3060.800 2773.600 ;
        RECT 3093.320 2772.480 3098.040 2773.600 ;
        RECT 23.060 2758.880 27.780 2760.000 ;
        RECT 111.900 2758.880 114.620 2760.000 ;
        RECT 29.060 2756.160 33.780 2757.280 ;
        RECT 107.100 2756.160 109.820 2757.280 ;
        RECT 35.060 2753.440 39.780 2754.560 ;
        RECT 78.300 2753.440 81.020 2754.560 ;
        RECT 41.060 2750.720 45.780 2751.840 ;
        RECT 83.100 2750.720 85.820 2751.840 ;
        RECT 47.060 2748.000 51.780 2749.120 ;
        RECT 87.900 2748.000 90.620 2749.120 ;
        RECT 53.060 2745.280 57.780 2746.400 ;
        RECT 92.700 2745.280 95.420 2746.400 ;
        RECT 59.060 2742.560 63.780 2743.680 ;
        RECT 97.500 2742.560 100.220 2743.680 ;
        RECT 65.060 2739.840 69.780 2740.960 ;
        RECT 102.300 2739.840 105.020 2740.960 ;
        RECT 3072.480 2715.360 3075.200 2716.480 ;
        RECT 3111.320 2715.360 3116.040 2716.480 ;
        RECT 3067.680 2712.640 3070.400 2713.760 ;
        RECT 3105.320 2712.640 3110.040 2713.760 ;
        RECT 3062.880 2709.920 3065.600 2711.040 ;
        RECT 3099.320 2709.920 3104.040 2711.040 ;
        RECT 3058.080 2707.200 3060.800 2708.320 ;
        RECT 3093.320 2707.200 3098.040 2708.320 ;
        RECT 23.060 2693.600 27.780 2694.720 ;
        RECT 111.900 2693.600 114.620 2694.720 ;
        RECT 29.060 2690.880 33.780 2692.000 ;
        RECT 107.100 2690.880 109.820 2692.000 ;
        RECT 35.060 2688.160 39.780 2689.280 ;
        RECT 78.300 2688.160 81.020 2689.280 ;
        RECT 41.060 2685.440 45.780 2686.560 ;
        RECT 83.100 2685.440 85.820 2686.560 ;
        RECT 47.060 2682.720 51.780 2683.840 ;
        RECT 87.900 2682.720 90.620 2683.840 ;
        RECT 53.060 2680.000 57.780 2681.120 ;
        RECT 92.700 2680.000 95.420 2681.120 ;
        RECT 59.060 2677.280 63.780 2678.400 ;
        RECT 97.500 2677.280 100.220 2678.400 ;
        RECT 65.060 2674.560 69.780 2675.680 ;
        RECT 102.300 2674.560 105.020 2675.680 ;
        RECT 3048.480 2652.800 3051.200 2653.920 ;
        RECT 3135.320 2652.800 3140.040 2653.920 ;
        RECT 3053.280 2650.080 3056.000 2651.200 ;
        RECT 3129.320 2650.080 3134.040 2651.200 ;
        RECT 3082.080 2647.360 3084.800 2648.480 ;
        RECT 3123.320 2647.360 3128.040 2648.480 ;
        RECT 3077.280 2644.640 3080.000 2645.760 ;
        RECT 3117.320 2644.640 3122.040 2645.760 ;
        RECT 3072.480 2641.920 3075.200 2643.040 ;
        RECT 3111.320 2641.920 3116.040 2643.040 ;
        RECT 3067.680 2639.200 3070.400 2640.320 ;
        RECT 3105.320 2639.200 3110.040 2640.320 ;
        RECT 3062.880 2636.480 3065.600 2637.600 ;
        RECT 3099.320 2636.480 3104.040 2637.600 ;
        RECT 3058.080 2633.760 3060.800 2634.880 ;
        RECT 3093.320 2633.760 3098.040 2634.880 ;
        RECT 23.060 2628.320 27.780 2629.440 ;
        RECT 111.900 2628.320 114.620 2629.440 ;
        RECT 29.060 2625.600 33.780 2626.720 ;
        RECT 107.100 2625.600 109.820 2626.720 ;
        RECT 35.060 2622.880 39.780 2624.000 ;
        RECT 78.300 2622.880 81.020 2624.000 ;
        RECT 41.060 2620.160 45.780 2621.280 ;
        RECT 83.100 2620.160 85.820 2621.280 ;
        RECT 47.060 2617.440 51.780 2618.560 ;
        RECT 87.900 2617.440 90.620 2618.560 ;
        RECT 53.060 2614.720 57.780 2615.840 ;
        RECT 92.700 2614.720 95.420 2615.840 ;
        RECT 59.060 2612.000 63.780 2613.120 ;
        RECT 97.500 2612.000 100.220 2613.120 ;
        RECT 65.060 2609.280 69.780 2610.400 ;
        RECT 102.300 2609.280 105.020 2610.400 ;
        RECT 3048.480 2587.520 3051.200 2588.640 ;
        RECT 3135.320 2587.520 3140.040 2588.640 ;
        RECT 3053.280 2584.800 3056.000 2585.920 ;
        RECT 3129.320 2584.800 3134.040 2585.920 ;
        RECT 3082.080 2582.080 3084.800 2583.200 ;
        RECT 3123.320 2582.080 3128.040 2583.200 ;
        RECT 3077.280 2579.360 3080.000 2580.480 ;
        RECT 3117.320 2579.360 3122.040 2580.480 ;
        RECT 3072.480 2576.640 3075.200 2577.760 ;
        RECT 3111.320 2576.640 3116.040 2577.760 ;
        RECT 3067.680 2573.920 3070.400 2575.040 ;
        RECT 3105.320 2573.920 3110.040 2575.040 ;
        RECT 3062.880 2571.200 3065.600 2572.320 ;
        RECT 3099.320 2571.200 3104.040 2572.320 ;
        RECT 3058.080 2568.480 3060.800 2569.600 ;
        RECT 3093.320 2568.480 3098.040 2569.600 ;
        RECT 23.060 2563.040 27.780 2564.160 ;
        RECT 111.900 2563.040 114.620 2564.160 ;
        RECT 29.060 2560.320 33.780 2561.440 ;
        RECT 107.100 2560.320 109.820 2561.440 ;
        RECT 35.060 2557.600 39.780 2558.720 ;
        RECT 78.300 2557.600 81.020 2558.720 ;
        RECT 41.060 2554.880 45.780 2556.000 ;
        RECT 83.100 2554.880 85.820 2556.000 ;
        RECT 47.060 2552.160 51.780 2553.280 ;
        RECT 87.900 2552.160 90.620 2553.280 ;
        RECT 53.060 2549.440 57.780 2550.560 ;
        RECT 92.700 2549.440 95.420 2550.560 ;
        RECT 59.060 2546.720 63.780 2547.840 ;
        RECT 97.500 2546.720 100.220 2547.840 ;
        RECT 65.060 2544.000 69.780 2545.120 ;
        RECT 102.300 2544.000 105.020 2545.120 ;
        RECT 3048.480 2522.240 3051.200 2523.360 ;
        RECT 3135.320 2522.240 3140.040 2523.360 ;
        RECT 3053.280 2519.520 3056.000 2520.640 ;
        RECT 3129.320 2519.520 3134.040 2520.640 ;
        RECT 3082.080 2516.800 3084.800 2517.920 ;
        RECT 3123.320 2516.800 3128.040 2517.920 ;
        RECT 3077.280 2514.080 3080.000 2515.200 ;
        RECT 3117.320 2514.080 3122.040 2515.200 ;
        RECT 3072.480 2511.360 3075.200 2512.480 ;
        RECT 3111.320 2511.360 3116.040 2512.480 ;
        RECT 3067.680 2508.640 3070.400 2509.760 ;
        RECT 3105.320 2508.640 3110.040 2509.760 ;
        RECT 3062.880 2505.920 3065.600 2507.040 ;
        RECT 3099.320 2505.920 3104.040 2507.040 ;
        RECT 3058.080 2503.200 3060.800 2504.320 ;
        RECT 3093.320 2503.200 3098.040 2504.320 ;
        RECT 23.060 2497.760 27.780 2498.880 ;
        RECT 111.900 2497.760 114.620 2498.880 ;
        RECT 29.060 2495.040 33.780 2496.160 ;
        RECT 107.100 2495.040 109.820 2496.160 ;
        RECT 35.060 2492.320 39.780 2493.440 ;
        RECT 78.300 2492.320 81.020 2493.440 ;
        RECT 41.060 2489.600 45.780 2490.720 ;
        RECT 83.100 2489.600 85.820 2490.720 ;
        RECT 47.060 2486.880 51.780 2488.000 ;
        RECT 87.900 2486.880 90.620 2488.000 ;
        RECT 53.060 2484.160 57.780 2485.280 ;
        RECT 92.700 2484.160 95.420 2485.280 ;
        RECT 59.060 2481.440 63.780 2482.560 ;
        RECT 97.500 2481.440 100.220 2482.560 ;
        RECT 65.060 2478.720 69.780 2479.840 ;
        RECT 102.300 2478.720 105.020 2479.840 ;
        RECT 3048.480 2456.960 3051.200 2458.080 ;
        RECT 3135.320 2456.960 3140.040 2458.080 ;
        RECT 3053.280 2454.240 3056.000 2455.360 ;
        RECT 3129.320 2454.240 3134.040 2455.360 ;
        RECT 3082.080 2451.520 3084.800 2452.640 ;
        RECT 3123.320 2451.520 3128.040 2452.640 ;
        RECT 3077.280 2448.800 3080.000 2449.920 ;
        RECT 3117.320 2448.800 3122.040 2449.920 ;
        RECT 3072.480 2446.080 3075.200 2447.200 ;
        RECT 3111.320 2446.080 3116.040 2447.200 ;
        RECT 3067.680 2443.360 3070.400 2444.480 ;
        RECT 3105.320 2443.360 3110.040 2444.480 ;
        RECT 3062.880 2440.640 3065.600 2441.760 ;
        RECT 3099.320 2440.640 3104.040 2441.760 ;
        RECT 3058.080 2437.920 3060.800 2439.040 ;
        RECT 3093.320 2437.920 3098.040 2439.040 ;
        RECT 23.060 2432.480 27.780 2433.600 ;
        RECT 111.900 2432.480 114.620 2433.600 ;
        RECT 29.060 2429.760 33.780 2430.880 ;
        RECT 107.100 2429.760 109.820 2430.880 ;
        RECT 35.060 2427.040 39.780 2428.160 ;
        RECT 78.300 2427.040 81.020 2428.160 ;
        RECT 41.060 2424.320 45.780 2425.440 ;
        RECT 83.100 2424.320 85.820 2425.440 ;
        RECT 47.060 2421.600 51.780 2422.720 ;
        RECT 87.900 2421.600 90.620 2422.720 ;
        RECT 53.060 2418.880 57.780 2420.000 ;
        RECT 92.700 2418.880 95.420 2420.000 ;
        RECT 59.060 2416.160 63.780 2417.280 ;
        RECT 97.500 2416.160 100.220 2417.280 ;
        RECT 65.060 2413.440 69.780 2414.560 ;
        RECT 102.300 2413.440 105.020 2414.560 ;
        RECT 3048.480 2383.520 3051.200 2384.640 ;
        RECT 3135.320 2383.520 3140.040 2384.640 ;
        RECT 3053.280 2380.800 3056.000 2381.920 ;
        RECT 3129.320 2380.800 3134.040 2381.920 ;
        RECT 3082.080 2378.080 3084.800 2379.200 ;
        RECT 3123.320 2378.080 3128.040 2379.200 ;
        RECT 3077.280 2375.360 3080.000 2376.480 ;
        RECT 3117.320 2375.360 3122.040 2376.480 ;
        RECT 3072.480 2372.640 3075.200 2373.760 ;
        RECT 3111.320 2372.640 3116.040 2373.760 ;
        RECT 3067.680 2369.920 3070.400 2371.040 ;
        RECT 3105.320 2369.920 3110.040 2371.040 ;
        RECT 3062.880 2367.200 3065.600 2368.320 ;
        RECT 3099.320 2367.200 3104.040 2368.320 ;
        RECT 3058.080 2364.480 3060.800 2365.600 ;
        RECT 3093.320 2364.480 3098.040 2365.600 ;
        RECT 23.060 2356.320 27.780 2357.440 ;
        RECT 111.900 2356.320 114.620 2357.440 ;
        RECT 29.060 2353.600 33.780 2354.720 ;
        RECT 107.100 2353.600 109.820 2354.720 ;
        RECT 35.060 2350.880 39.780 2352.000 ;
        RECT 78.300 2350.880 81.020 2352.000 ;
        RECT 41.060 2348.160 45.780 2349.280 ;
        RECT 83.100 2348.160 85.820 2349.280 ;
        RECT 47.060 2345.440 51.780 2346.560 ;
        RECT 87.900 2345.440 90.620 2346.560 ;
        RECT 53.060 2342.720 57.780 2343.840 ;
        RECT 92.700 2342.720 95.420 2343.840 ;
        RECT 59.060 2340.000 63.780 2341.120 ;
        RECT 97.500 2340.000 100.220 2341.120 ;
        RECT 65.060 2337.280 69.780 2338.400 ;
        RECT 102.300 2337.280 105.020 2338.400 ;
        RECT 3048.480 2318.240 3051.200 2319.360 ;
        RECT 3135.320 2318.240 3140.040 2319.360 ;
        RECT 3053.280 2315.520 3056.000 2316.640 ;
        RECT 3129.320 2315.520 3134.040 2316.640 ;
        RECT 3082.080 2312.800 3084.800 2313.920 ;
        RECT 3123.320 2312.800 3128.040 2313.920 ;
        RECT 3077.280 2310.080 3080.000 2311.200 ;
        RECT 3117.320 2310.080 3122.040 2311.200 ;
        RECT 3072.480 2307.360 3075.200 2308.480 ;
        RECT 3111.320 2307.360 3116.040 2308.480 ;
        RECT 3067.680 2304.640 3070.400 2305.760 ;
        RECT 3105.320 2304.640 3110.040 2305.760 ;
        RECT 23.060 2301.920 27.780 2303.040 ;
        RECT 111.900 2301.920 114.620 2303.040 ;
        RECT 3062.880 2301.920 3065.600 2303.040 ;
        RECT 3099.320 2301.920 3104.040 2303.040 ;
        RECT 29.060 2299.200 33.780 2300.320 ;
        RECT 107.100 2299.200 109.820 2300.320 ;
        RECT 3058.080 2299.200 3060.800 2300.320 ;
        RECT 3093.320 2299.200 3098.040 2300.320 ;
        RECT 35.060 2296.480 39.780 2297.600 ;
        RECT 78.300 2296.480 81.020 2297.600 ;
        RECT 41.060 2293.760 45.780 2294.880 ;
        RECT 83.100 2293.760 85.820 2294.880 ;
        RECT 47.060 2291.040 51.780 2292.160 ;
        RECT 87.900 2291.040 90.620 2292.160 ;
        RECT 53.060 2288.320 57.780 2289.440 ;
        RECT 92.700 2288.320 95.420 2289.440 ;
        RECT 59.060 2285.600 63.780 2286.720 ;
        RECT 97.500 2285.600 100.220 2286.720 ;
        RECT 65.060 2282.880 69.780 2284.000 ;
        RECT 102.300 2282.880 105.020 2284.000 ;
        RECT 3048.480 2252.960 3051.200 2254.080 ;
        RECT 3135.320 2252.960 3140.040 2254.080 ;
        RECT 3053.280 2250.240 3056.000 2251.360 ;
        RECT 3129.320 2250.240 3134.040 2251.360 ;
        RECT 3082.080 2247.520 3084.800 2248.640 ;
        RECT 3123.320 2247.520 3128.040 2248.640 ;
        RECT 3077.280 2244.800 3080.000 2245.920 ;
        RECT 3117.320 2244.800 3122.040 2245.920 ;
        RECT 3072.480 2242.080 3075.200 2243.200 ;
        RECT 3111.320 2242.080 3116.040 2243.200 ;
        RECT 3067.680 2239.360 3070.400 2240.480 ;
        RECT 3105.320 2239.360 3110.040 2240.480 ;
        RECT 23.060 2236.640 27.780 2237.760 ;
        RECT 111.900 2236.640 114.620 2237.760 ;
        RECT 3062.880 2236.640 3065.600 2237.760 ;
        RECT 3099.320 2236.640 3104.040 2237.760 ;
        RECT 29.060 2233.920 33.780 2235.040 ;
        RECT 107.100 2233.920 109.820 2235.040 ;
        RECT 3058.080 2233.920 3060.800 2235.040 ;
        RECT 3093.320 2233.920 3098.040 2235.040 ;
        RECT 35.060 2231.200 39.780 2232.320 ;
        RECT 78.300 2231.200 81.020 2232.320 ;
        RECT 41.060 2228.480 45.780 2229.600 ;
        RECT 83.100 2228.480 85.820 2229.600 ;
        RECT 47.060 2225.760 51.780 2226.880 ;
        RECT 87.900 2225.760 90.620 2226.880 ;
        RECT 53.060 2223.040 57.780 2224.160 ;
        RECT 92.700 2223.040 95.420 2224.160 ;
        RECT 59.060 2220.320 63.780 2221.440 ;
        RECT 97.500 2220.320 100.220 2221.440 ;
        RECT 65.060 2217.600 69.780 2218.720 ;
        RECT 102.300 2217.600 105.020 2218.720 ;
        RECT 3048.480 2187.680 3051.200 2188.800 ;
        RECT 3135.320 2187.680 3140.040 2188.800 ;
        RECT 3053.280 2184.960 3056.000 2186.080 ;
        RECT 3129.320 2184.960 3134.040 2186.080 ;
        RECT 3082.080 2182.240 3084.800 2183.360 ;
        RECT 3123.320 2182.240 3128.040 2183.360 ;
        RECT 3077.280 2179.520 3080.000 2180.640 ;
        RECT 3117.320 2179.520 3122.040 2180.640 ;
        RECT 3072.480 2176.800 3075.200 2177.920 ;
        RECT 3111.320 2176.800 3116.040 2177.920 ;
        RECT 3067.680 2174.080 3070.400 2175.200 ;
        RECT 3105.320 2174.080 3110.040 2175.200 ;
        RECT 23.060 2171.360 27.780 2172.480 ;
        RECT 111.900 2171.360 114.620 2172.480 ;
        RECT 3062.880 2171.360 3065.600 2172.480 ;
        RECT 3099.320 2171.360 3104.040 2172.480 ;
        RECT 29.060 2168.640 33.780 2169.760 ;
        RECT 107.100 2168.640 109.820 2169.760 ;
        RECT 3058.080 2168.640 3060.800 2169.760 ;
        RECT 3093.320 2168.640 3098.040 2169.760 ;
        RECT 35.060 2165.920 39.780 2167.040 ;
        RECT 78.300 2165.920 81.020 2167.040 ;
        RECT 41.060 2163.200 45.780 2164.320 ;
        RECT 83.100 2163.200 85.820 2164.320 ;
        RECT 47.060 2160.480 51.780 2161.600 ;
        RECT 87.900 2160.480 90.620 2161.600 ;
        RECT 53.060 2157.760 57.780 2158.880 ;
        RECT 92.700 2157.760 95.420 2158.880 ;
        RECT 59.060 2155.040 63.780 2156.160 ;
        RECT 97.500 2155.040 100.220 2156.160 ;
        RECT 65.060 2152.320 69.780 2153.440 ;
        RECT 102.300 2152.320 105.020 2153.440 ;
        RECT 3048.480 2122.400 3051.200 2123.520 ;
        RECT 3135.320 2122.400 3140.040 2123.520 ;
        RECT 3053.280 2119.680 3056.000 2120.800 ;
        RECT 3129.320 2119.680 3134.040 2120.800 ;
        RECT 3082.080 2116.960 3084.800 2118.080 ;
        RECT 3123.320 2116.960 3128.040 2118.080 ;
        RECT 3077.280 2114.240 3080.000 2115.360 ;
        RECT 3117.320 2114.240 3122.040 2115.360 ;
        RECT 3072.480 2111.520 3075.200 2112.640 ;
        RECT 3111.320 2111.520 3116.040 2112.640 ;
        RECT 3067.680 2108.800 3070.400 2109.920 ;
        RECT 3105.320 2108.800 3110.040 2109.920 ;
        RECT 23.060 2106.080 27.780 2107.200 ;
        RECT 111.900 2106.080 114.620 2107.200 ;
        RECT 3062.880 2106.080 3065.600 2107.200 ;
        RECT 3099.320 2106.080 3104.040 2107.200 ;
        RECT 29.060 2103.360 33.780 2104.480 ;
        RECT 107.100 2103.360 109.820 2104.480 ;
        RECT 3058.080 2103.360 3060.800 2104.480 ;
        RECT 3093.320 2103.360 3098.040 2104.480 ;
        RECT 35.060 2100.640 39.780 2101.760 ;
        RECT 78.300 2100.640 81.020 2101.760 ;
        RECT 41.060 2097.920 45.780 2099.040 ;
        RECT 83.100 2097.920 85.820 2099.040 ;
        RECT 47.060 2095.200 51.780 2096.320 ;
        RECT 87.900 2095.200 90.620 2096.320 ;
        RECT 53.060 2092.480 57.780 2093.600 ;
        RECT 92.700 2092.480 95.420 2093.600 ;
        RECT 59.060 2089.760 63.780 2090.880 ;
        RECT 97.500 2089.760 100.220 2090.880 ;
        RECT 65.060 2087.040 69.780 2088.160 ;
        RECT 102.300 2087.040 105.020 2088.160 ;
        RECT 3048.480 2057.120 3051.200 2058.240 ;
        RECT 3135.320 2057.120 3140.040 2058.240 ;
        RECT 3053.280 2054.400 3056.000 2055.520 ;
        RECT 3129.320 2054.400 3134.040 2055.520 ;
        RECT 3082.080 2051.680 3084.800 2052.800 ;
        RECT 3123.320 2051.680 3128.040 2052.800 ;
        RECT 3077.280 2048.960 3080.000 2050.080 ;
        RECT 3117.320 2048.960 3122.040 2050.080 ;
        RECT 3072.480 2046.240 3075.200 2047.360 ;
        RECT 3111.320 2046.240 3116.040 2047.360 ;
        RECT 3067.680 2043.520 3070.400 2044.640 ;
        RECT 3105.320 2043.520 3110.040 2044.640 ;
        RECT 23.060 2040.800 27.780 2041.920 ;
        RECT 111.900 2040.800 114.620 2041.920 ;
        RECT 3062.880 2040.800 3065.600 2041.920 ;
        RECT 3099.320 2040.800 3104.040 2041.920 ;
        RECT 29.060 2038.080 33.780 2039.200 ;
        RECT 107.100 2038.080 109.820 2039.200 ;
        RECT 3058.080 2038.080 3060.800 2039.200 ;
        RECT 3093.320 2038.080 3098.040 2039.200 ;
        RECT 35.060 2035.360 39.780 2036.480 ;
        RECT 78.300 2035.360 81.020 2036.480 ;
        RECT 41.060 2032.640 45.780 2033.760 ;
        RECT 83.100 2032.640 85.820 2033.760 ;
        RECT 47.060 2029.920 51.780 2031.040 ;
        RECT 87.900 2029.920 90.620 2031.040 ;
        RECT 53.060 2027.200 57.780 2028.320 ;
        RECT 92.700 2027.200 95.420 2028.320 ;
        RECT 59.060 2024.480 63.780 2025.600 ;
        RECT 97.500 2024.480 100.220 2025.600 ;
        RECT 65.060 2021.760 69.780 2022.880 ;
        RECT 102.300 2021.760 105.020 2022.880 ;
        RECT 3048.480 1991.840 3051.200 1992.960 ;
        RECT 3135.320 1991.840 3140.040 1992.960 ;
        RECT 3053.280 1989.120 3056.000 1990.240 ;
        RECT 3129.320 1989.120 3134.040 1990.240 ;
        RECT 3082.080 1986.400 3084.800 1987.520 ;
        RECT 3123.320 1986.400 3128.040 1987.520 ;
        RECT 3077.280 1983.680 3080.000 1984.800 ;
        RECT 3117.320 1983.680 3122.040 1984.800 ;
        RECT 3072.480 1980.960 3075.200 1982.080 ;
        RECT 3111.320 1980.960 3116.040 1982.080 ;
        RECT 3067.680 1978.240 3070.400 1979.360 ;
        RECT 3105.320 1978.240 3110.040 1979.360 ;
        RECT 23.060 1975.520 27.780 1976.640 ;
        RECT 111.900 1975.520 114.620 1976.640 ;
        RECT 3062.880 1975.520 3065.600 1976.640 ;
        RECT 3099.320 1975.520 3104.040 1976.640 ;
        RECT 29.060 1972.800 33.780 1973.920 ;
        RECT 107.100 1972.800 109.820 1973.920 ;
        RECT 3058.080 1972.800 3060.800 1973.920 ;
        RECT 3093.320 1972.800 3098.040 1973.920 ;
        RECT 35.060 1970.080 39.780 1971.200 ;
        RECT 78.300 1970.080 81.020 1971.200 ;
        RECT 41.060 1967.360 45.780 1968.480 ;
        RECT 83.100 1967.360 85.820 1968.480 ;
        RECT 47.060 1964.640 51.780 1965.760 ;
        RECT 87.900 1964.640 90.620 1965.760 ;
        RECT 53.060 1961.920 57.780 1963.040 ;
        RECT 92.700 1961.920 95.420 1963.040 ;
        RECT 59.060 1959.200 63.780 1960.320 ;
        RECT 97.500 1959.200 100.220 1960.320 ;
        RECT 65.060 1956.480 69.780 1957.600 ;
        RECT 102.300 1956.480 105.020 1957.600 ;
        RECT 3048.480 1926.560 3051.200 1927.680 ;
        RECT 3135.320 1926.560 3140.040 1927.680 ;
        RECT 3053.280 1923.840 3056.000 1924.960 ;
        RECT 3129.320 1923.840 3134.040 1924.960 ;
        RECT 3082.080 1921.120 3084.800 1922.240 ;
        RECT 3123.320 1921.120 3128.040 1922.240 ;
        RECT 3077.280 1918.400 3080.000 1919.520 ;
        RECT 3117.320 1918.400 3122.040 1919.520 ;
        RECT 3072.480 1915.680 3075.200 1916.800 ;
        RECT 3111.320 1915.680 3116.040 1916.800 ;
        RECT 3067.680 1912.960 3070.400 1914.080 ;
        RECT 3105.320 1912.960 3110.040 1914.080 ;
        RECT 23.060 1910.240 27.780 1911.360 ;
        RECT 111.900 1910.240 114.620 1911.360 ;
        RECT 3062.880 1910.240 3065.600 1911.360 ;
        RECT 3099.320 1910.240 3104.040 1911.360 ;
        RECT 29.060 1907.520 33.780 1908.640 ;
        RECT 107.100 1907.520 109.820 1908.640 ;
        RECT 3058.080 1907.520 3060.800 1908.640 ;
        RECT 3093.320 1907.520 3098.040 1908.640 ;
        RECT 35.060 1904.800 39.780 1905.920 ;
        RECT 78.300 1904.800 81.020 1905.920 ;
        RECT 41.060 1902.080 45.780 1903.200 ;
        RECT 83.100 1902.080 85.820 1903.200 ;
        RECT 47.060 1899.360 51.780 1900.480 ;
        RECT 87.900 1899.360 90.620 1900.480 ;
        RECT 53.060 1896.640 57.780 1897.760 ;
        RECT 92.700 1896.640 95.420 1897.760 ;
        RECT 59.060 1893.920 63.780 1895.040 ;
        RECT 97.500 1893.920 100.220 1895.040 ;
        RECT 65.060 1891.200 69.780 1892.320 ;
        RECT 102.300 1891.200 105.020 1892.320 ;
        RECT 23.060 1844.960 27.780 1846.080 ;
        RECT 111.900 1844.960 114.620 1846.080 ;
        RECT 3048.480 1844.960 3051.200 1846.080 ;
        RECT 3135.320 1844.960 3140.040 1846.080 ;
        RECT 29.060 1842.240 33.780 1843.360 ;
        RECT 107.100 1842.240 109.820 1843.360 ;
        RECT 3053.280 1842.240 3056.000 1843.360 ;
        RECT 3129.320 1842.240 3134.040 1843.360 ;
        RECT 35.060 1839.520 39.780 1840.640 ;
        RECT 78.300 1839.520 81.020 1840.640 ;
        RECT 3082.080 1839.520 3084.800 1840.640 ;
        RECT 3123.320 1839.520 3128.040 1840.640 ;
        RECT 41.060 1836.800 45.780 1837.920 ;
        RECT 83.100 1836.800 85.820 1837.920 ;
        RECT 3077.280 1836.800 3080.000 1837.920 ;
        RECT 3117.320 1836.800 3122.040 1837.920 ;
        RECT 47.060 1834.080 51.780 1835.200 ;
        RECT 87.900 1834.080 90.620 1835.200 ;
        RECT 3072.480 1834.080 3075.200 1835.200 ;
        RECT 3111.320 1834.080 3116.040 1835.200 ;
        RECT 53.060 1831.360 57.780 1832.480 ;
        RECT 92.700 1831.360 95.420 1832.480 ;
        RECT 3067.680 1831.360 3070.400 1832.480 ;
        RECT 3105.320 1831.360 3110.040 1832.480 ;
        RECT 59.060 1828.640 63.780 1829.760 ;
        RECT 97.500 1828.640 100.220 1829.760 ;
        RECT 3062.880 1828.640 3065.600 1829.760 ;
        RECT 3099.320 1828.640 3104.040 1829.760 ;
        RECT 65.060 1825.920 69.780 1827.040 ;
        RECT 102.300 1825.920 105.020 1827.040 ;
        RECT 3058.080 1825.920 3060.800 1827.040 ;
        RECT 3093.320 1825.920 3098.040 1827.040 ;
        RECT 23.060 1779.680 27.780 1780.800 ;
        RECT 111.900 1779.680 114.620 1780.800 ;
        RECT 3048.480 1779.680 3051.200 1780.800 ;
        RECT 3135.320 1779.680 3140.040 1780.800 ;
        RECT 29.060 1776.960 33.780 1778.080 ;
        RECT 107.100 1776.960 109.820 1778.080 ;
        RECT 3053.280 1776.960 3056.000 1778.080 ;
        RECT 3129.320 1776.960 3134.040 1778.080 ;
        RECT 35.060 1774.240 39.780 1775.360 ;
        RECT 78.300 1774.240 81.020 1775.360 ;
        RECT 3082.080 1774.240 3084.800 1775.360 ;
        RECT 3123.320 1774.240 3128.040 1775.360 ;
        RECT 41.060 1771.520 45.780 1772.640 ;
        RECT 83.100 1771.520 85.820 1772.640 ;
        RECT 3077.280 1771.520 3080.000 1772.640 ;
        RECT 3117.320 1771.520 3122.040 1772.640 ;
        RECT 47.060 1768.800 51.780 1769.920 ;
        RECT 87.900 1768.800 90.620 1769.920 ;
        RECT 3072.480 1768.800 3075.200 1769.920 ;
        RECT 3111.320 1768.800 3116.040 1769.920 ;
        RECT 53.060 1766.080 57.780 1767.200 ;
        RECT 92.700 1766.080 95.420 1767.200 ;
        RECT 3067.680 1766.080 3070.400 1767.200 ;
        RECT 3105.320 1766.080 3110.040 1767.200 ;
        RECT 59.060 1763.360 63.780 1764.480 ;
        RECT 97.500 1763.360 100.220 1764.480 ;
        RECT 3062.880 1763.360 3065.600 1764.480 ;
        RECT 3099.320 1763.360 3104.040 1764.480 ;
        RECT 65.060 1760.640 69.780 1761.760 ;
        RECT 102.300 1760.640 105.020 1761.760 ;
        RECT 3058.080 1760.640 3060.800 1761.760 ;
        RECT 3093.320 1760.640 3098.040 1761.760 ;
        RECT 3048.480 1714.400 3051.200 1715.520 ;
        RECT 3135.320 1714.400 3140.040 1715.520 ;
        RECT 3053.280 1711.680 3056.000 1712.800 ;
        RECT 3129.320 1711.680 3134.040 1712.800 ;
        RECT 3082.080 1708.960 3084.800 1710.080 ;
        RECT 3123.320 1708.960 3128.040 1710.080 ;
        RECT 3077.280 1706.240 3080.000 1707.360 ;
        RECT 3117.320 1706.240 3122.040 1707.360 ;
        RECT 23.060 1703.520 27.780 1704.640 ;
        RECT 111.900 1703.520 114.620 1704.640 ;
        RECT 3072.480 1703.520 3075.200 1704.640 ;
        RECT 3111.320 1703.520 3116.040 1704.640 ;
        RECT 29.060 1700.800 33.780 1701.920 ;
        RECT 107.100 1700.800 109.820 1701.920 ;
        RECT 3067.680 1700.800 3070.400 1701.920 ;
        RECT 3105.320 1700.800 3110.040 1701.920 ;
        RECT 35.060 1698.080 39.780 1699.200 ;
        RECT 78.300 1698.080 81.020 1699.200 ;
        RECT 3062.880 1698.080 3065.600 1699.200 ;
        RECT 3099.320 1698.080 3104.040 1699.200 ;
        RECT 41.060 1695.360 45.780 1696.480 ;
        RECT 83.100 1695.360 85.820 1696.480 ;
        RECT 3058.080 1695.360 3060.800 1696.480 ;
        RECT 3093.320 1695.360 3098.040 1696.480 ;
        RECT 47.060 1692.640 51.780 1693.760 ;
        RECT 87.900 1692.640 90.620 1693.760 ;
        RECT 53.060 1689.920 57.780 1691.040 ;
        RECT 92.700 1689.920 95.420 1691.040 ;
        RECT 59.060 1687.200 63.780 1688.320 ;
        RECT 97.500 1687.200 100.220 1688.320 ;
        RECT 65.060 1684.480 69.780 1685.600 ;
        RECT 102.300 1684.480 105.020 1685.600 ;
        RECT 23.060 1649.120 27.780 1650.240 ;
        RECT 111.900 1649.120 114.620 1650.240 ;
        RECT 3048.480 1649.120 3051.200 1650.240 ;
        RECT 3135.320 1649.120 3140.040 1650.240 ;
        RECT 29.060 1646.400 33.780 1647.520 ;
        RECT 107.100 1646.400 109.820 1647.520 ;
        RECT 3053.280 1646.400 3056.000 1647.520 ;
        RECT 3129.320 1646.400 3134.040 1647.520 ;
        RECT 35.060 1643.680 39.780 1644.800 ;
        RECT 78.300 1643.680 81.020 1644.800 ;
        RECT 3082.080 1643.680 3084.800 1644.800 ;
        RECT 3123.320 1643.680 3128.040 1644.800 ;
        RECT 41.060 1640.960 45.780 1642.080 ;
        RECT 83.100 1640.960 85.820 1642.080 ;
        RECT 3077.280 1640.960 3080.000 1642.080 ;
        RECT 3117.320 1640.960 3122.040 1642.080 ;
        RECT 47.060 1638.240 51.780 1639.360 ;
        RECT 87.900 1638.240 90.620 1639.360 ;
        RECT 3072.480 1638.240 3075.200 1639.360 ;
        RECT 3111.320 1638.240 3116.040 1639.360 ;
        RECT 53.060 1635.520 57.780 1636.640 ;
        RECT 92.700 1635.520 95.420 1636.640 ;
        RECT 3067.680 1635.520 3070.400 1636.640 ;
        RECT 3105.320 1635.520 3110.040 1636.640 ;
        RECT 59.060 1632.800 63.780 1633.920 ;
        RECT 97.500 1632.800 100.220 1633.920 ;
        RECT 3062.880 1632.800 3065.600 1633.920 ;
        RECT 3099.320 1632.800 3104.040 1633.920 ;
        RECT 65.060 1630.080 69.780 1631.200 ;
        RECT 102.300 1630.080 105.020 1631.200 ;
        RECT 3058.080 1630.080 3060.800 1631.200 ;
        RECT 3093.320 1630.080 3098.040 1631.200 ;
        RECT 3048.480 1592.000 3051.200 1593.120 ;
        RECT 3135.320 1592.000 3140.040 1593.120 ;
        RECT 3053.280 1589.280 3056.000 1590.400 ;
        RECT 3129.320 1589.280 3134.040 1590.400 ;
        RECT 3082.080 1586.560 3084.800 1587.680 ;
        RECT 3123.320 1586.560 3128.040 1587.680 ;
        RECT 23.060 1583.840 27.780 1584.960 ;
        RECT 111.900 1583.840 114.620 1584.960 ;
        RECT 3077.280 1583.840 3080.000 1584.960 ;
        RECT 3117.320 1583.840 3122.040 1584.960 ;
        RECT 29.060 1581.120 33.780 1582.240 ;
        RECT 107.100 1581.120 109.820 1582.240 ;
        RECT 3072.480 1581.120 3075.200 1582.240 ;
        RECT 3111.320 1581.120 3116.040 1582.240 ;
        RECT 35.060 1578.400 39.780 1579.520 ;
        RECT 78.300 1578.400 81.020 1579.520 ;
        RECT 3067.680 1578.400 3070.400 1579.520 ;
        RECT 3105.320 1578.400 3110.040 1579.520 ;
        RECT 41.060 1575.680 45.780 1576.800 ;
        RECT 83.100 1575.680 85.820 1576.800 ;
        RECT 3062.880 1575.680 3065.600 1576.800 ;
        RECT 3099.320 1575.680 3104.040 1576.800 ;
        RECT 47.060 1572.960 51.780 1574.080 ;
        RECT 87.900 1572.960 90.620 1574.080 ;
        RECT 3058.080 1572.960 3060.800 1574.080 ;
        RECT 3093.320 1572.960 3098.040 1574.080 ;
        RECT 53.060 1570.240 57.780 1571.360 ;
        RECT 92.700 1570.240 95.420 1571.360 ;
        RECT 59.060 1567.520 63.780 1568.640 ;
        RECT 97.500 1567.520 100.220 1568.640 ;
        RECT 65.060 1564.800 69.780 1565.920 ;
        RECT 102.300 1564.800 105.020 1565.920 ;
        RECT 23.060 1529.440 27.780 1530.560 ;
        RECT 111.900 1529.440 114.620 1530.560 ;
        RECT 29.060 1526.720 33.780 1527.840 ;
        RECT 107.100 1526.720 109.820 1527.840 ;
        RECT 35.060 1524.000 39.780 1525.120 ;
        RECT 78.300 1524.000 81.020 1525.120 ;
        RECT 41.060 1521.280 45.780 1522.400 ;
        RECT 83.100 1521.280 85.820 1522.400 ;
        RECT 47.060 1518.560 51.780 1519.680 ;
        RECT 87.900 1518.560 90.620 1519.680 ;
        RECT 3048.480 1518.560 3051.200 1519.680 ;
        RECT 3135.320 1518.560 3140.040 1519.680 ;
        RECT 53.060 1515.840 57.780 1516.960 ;
        RECT 92.700 1515.840 95.420 1516.960 ;
        RECT 3053.280 1515.840 3056.000 1516.960 ;
        RECT 3129.320 1515.840 3134.040 1516.960 ;
        RECT 59.060 1513.120 63.780 1514.240 ;
        RECT 97.500 1513.120 100.220 1514.240 ;
        RECT 3082.080 1513.120 3084.800 1514.240 ;
        RECT 3123.320 1513.120 3128.040 1514.240 ;
        RECT 65.060 1510.400 69.780 1511.520 ;
        RECT 102.300 1510.400 105.020 1511.520 ;
        RECT 3077.280 1510.400 3080.000 1511.520 ;
        RECT 3117.320 1510.400 3122.040 1511.520 ;
        RECT 3072.480 1507.680 3075.200 1508.800 ;
        RECT 3111.320 1507.680 3116.040 1508.800 ;
        RECT 3067.680 1504.960 3070.400 1506.080 ;
        RECT 3105.320 1504.960 3110.040 1506.080 ;
        RECT 3062.880 1502.240 3065.600 1503.360 ;
        RECT 3099.320 1502.240 3104.040 1503.360 ;
        RECT 3058.080 1499.520 3060.800 1500.640 ;
        RECT 3093.320 1499.520 3098.040 1500.640 ;
        RECT 23.060 1453.280 27.780 1454.400 ;
        RECT 111.900 1453.280 114.620 1454.400 ;
        RECT 3048.480 1453.280 3051.200 1454.400 ;
        RECT 3135.320 1453.280 3140.040 1454.400 ;
        RECT 29.060 1450.560 33.780 1451.680 ;
        RECT 107.100 1450.560 109.820 1451.680 ;
        RECT 3053.280 1450.560 3056.000 1451.680 ;
        RECT 3129.320 1450.560 3134.040 1451.680 ;
        RECT 35.060 1447.840 39.780 1448.960 ;
        RECT 78.300 1447.840 81.020 1448.960 ;
        RECT 3082.080 1447.840 3084.800 1448.960 ;
        RECT 3123.320 1447.840 3128.040 1448.960 ;
        RECT 41.060 1445.120 45.780 1446.240 ;
        RECT 83.100 1445.120 85.820 1446.240 ;
        RECT 3077.280 1445.120 3080.000 1446.240 ;
        RECT 3117.320 1445.120 3122.040 1446.240 ;
        RECT 47.060 1442.400 51.780 1443.520 ;
        RECT 87.900 1442.400 90.620 1443.520 ;
        RECT 3072.480 1442.400 3075.200 1443.520 ;
        RECT 3111.320 1442.400 3116.040 1443.520 ;
        RECT 53.060 1439.680 57.780 1440.800 ;
        RECT 92.700 1439.680 95.420 1440.800 ;
        RECT 3067.680 1439.680 3070.400 1440.800 ;
        RECT 3105.320 1439.680 3110.040 1440.800 ;
        RECT 59.060 1436.960 63.780 1438.080 ;
        RECT 97.500 1436.960 100.220 1438.080 ;
        RECT 3062.880 1436.960 3065.600 1438.080 ;
        RECT 3099.320 1436.960 3104.040 1438.080 ;
        RECT 65.060 1434.240 69.780 1435.360 ;
        RECT 102.300 1434.240 105.020 1435.360 ;
        RECT 3058.080 1434.240 3060.800 1435.360 ;
        RECT 3093.320 1434.240 3098.040 1435.360 ;
        RECT 23.060 1388.000 27.780 1389.120 ;
        RECT 111.900 1388.000 114.620 1389.120 ;
        RECT 3048.480 1388.000 3051.200 1389.120 ;
        RECT 3135.320 1388.000 3140.040 1389.120 ;
        RECT 29.060 1385.280 33.780 1386.400 ;
        RECT 107.100 1385.280 109.820 1386.400 ;
        RECT 3053.280 1385.280 3056.000 1386.400 ;
        RECT 3129.320 1385.280 3134.040 1386.400 ;
        RECT 35.060 1382.560 39.780 1383.680 ;
        RECT 78.300 1382.560 81.020 1383.680 ;
        RECT 3082.080 1382.560 3084.800 1383.680 ;
        RECT 3123.320 1382.560 3128.040 1383.680 ;
        RECT 41.060 1379.840 45.780 1380.960 ;
        RECT 83.100 1379.840 85.820 1380.960 ;
        RECT 3077.280 1379.840 3080.000 1380.960 ;
        RECT 3117.320 1379.840 3122.040 1380.960 ;
        RECT 47.060 1377.120 51.780 1378.240 ;
        RECT 87.900 1377.120 90.620 1378.240 ;
        RECT 3072.480 1377.120 3075.200 1378.240 ;
        RECT 3111.320 1377.120 3116.040 1378.240 ;
        RECT 53.060 1374.400 57.780 1375.520 ;
        RECT 92.700 1374.400 95.420 1375.520 ;
        RECT 3067.680 1374.400 3070.400 1375.520 ;
        RECT 3105.320 1374.400 3110.040 1375.520 ;
        RECT 59.060 1371.680 63.780 1372.800 ;
        RECT 97.500 1371.680 100.220 1372.800 ;
        RECT 3062.880 1371.680 3065.600 1372.800 ;
        RECT 3099.320 1371.680 3104.040 1372.800 ;
        RECT 65.060 1368.960 69.780 1370.080 ;
        RECT 102.300 1368.960 105.020 1370.080 ;
        RECT 3058.080 1368.960 3060.800 1370.080 ;
        RECT 3093.320 1368.960 3098.040 1370.080 ;
        RECT 23.060 1333.600 27.780 1334.720 ;
        RECT 111.900 1333.600 114.620 1334.720 ;
        RECT 29.060 1330.880 33.780 1332.000 ;
        RECT 107.100 1330.880 109.820 1332.000 ;
        RECT 35.060 1328.160 39.780 1329.280 ;
        RECT 78.300 1328.160 81.020 1329.280 ;
        RECT 41.060 1325.440 45.780 1326.560 ;
        RECT 83.100 1325.440 85.820 1326.560 ;
        RECT 47.060 1322.720 51.780 1323.840 ;
        RECT 87.900 1322.720 90.620 1323.840 ;
        RECT 53.060 1320.000 57.780 1321.120 ;
        RECT 92.700 1320.000 95.420 1321.120 ;
        RECT 59.060 1317.280 63.780 1318.400 ;
        RECT 97.500 1317.280 100.220 1318.400 ;
        RECT 65.060 1314.560 69.780 1315.680 ;
        RECT 102.300 1314.560 105.020 1315.680 ;
        RECT 3048.480 1314.560 3051.200 1315.680 ;
        RECT 3135.320 1314.560 3140.040 1315.680 ;
        RECT 3053.280 1311.840 3056.000 1312.960 ;
        RECT 3129.320 1311.840 3134.040 1312.960 ;
        RECT 3082.080 1309.120 3084.800 1310.240 ;
        RECT 3123.320 1309.120 3128.040 1310.240 ;
        RECT 3077.280 1306.400 3080.000 1307.520 ;
        RECT 3117.320 1306.400 3122.040 1307.520 ;
        RECT 3072.480 1303.680 3075.200 1304.800 ;
        RECT 3111.320 1303.680 3116.040 1304.800 ;
        RECT 3067.680 1300.960 3070.400 1302.080 ;
        RECT 3105.320 1300.960 3110.040 1302.080 ;
        RECT 3062.880 1298.240 3065.600 1299.360 ;
        RECT 3099.320 1298.240 3104.040 1299.360 ;
        RECT 3058.080 1295.520 3060.800 1296.640 ;
        RECT 3093.320 1295.520 3098.040 1296.640 ;
        RECT 23.060 1257.440 27.780 1258.560 ;
        RECT 111.900 1257.440 114.620 1258.560 ;
        RECT 3048.480 1257.440 3051.200 1258.560 ;
        RECT 3135.320 1257.440 3140.040 1258.560 ;
        RECT 29.060 1254.720 33.780 1255.840 ;
        RECT 107.100 1254.720 109.820 1255.840 ;
        RECT 3053.280 1254.720 3056.000 1255.840 ;
        RECT 3129.320 1254.720 3134.040 1255.840 ;
        RECT 35.060 1252.000 39.780 1253.120 ;
        RECT 78.300 1252.000 81.020 1253.120 ;
        RECT 3082.080 1252.000 3084.800 1253.120 ;
        RECT 3123.320 1252.000 3128.040 1253.120 ;
        RECT 41.060 1249.280 45.780 1250.400 ;
        RECT 83.100 1249.280 85.820 1250.400 ;
        RECT 3077.280 1249.280 3080.000 1250.400 ;
        RECT 3117.320 1249.280 3122.040 1250.400 ;
        RECT 47.060 1246.560 51.780 1247.680 ;
        RECT 87.900 1246.560 90.620 1247.680 ;
        RECT 3072.480 1246.560 3075.200 1247.680 ;
        RECT 3111.320 1246.560 3116.040 1247.680 ;
        RECT 53.060 1243.840 57.780 1244.960 ;
        RECT 92.700 1243.840 95.420 1244.960 ;
        RECT 3067.680 1243.840 3070.400 1244.960 ;
        RECT 3105.320 1243.840 3110.040 1244.960 ;
        RECT 59.060 1241.120 63.780 1242.240 ;
        RECT 97.500 1241.120 100.220 1242.240 ;
        RECT 3062.880 1241.120 3065.600 1242.240 ;
        RECT 3099.320 1241.120 3104.040 1242.240 ;
        RECT 65.060 1238.400 69.780 1239.520 ;
        RECT 102.300 1238.400 105.020 1239.520 ;
        RECT 3058.080 1238.400 3060.800 1239.520 ;
        RECT 3093.320 1238.400 3098.040 1239.520 ;
        RECT 23.060 1192.160 27.780 1193.280 ;
        RECT 111.900 1192.160 114.620 1193.280 ;
        RECT 3048.480 1192.160 3051.200 1193.280 ;
        RECT 3135.320 1192.160 3140.040 1193.280 ;
        RECT 29.060 1189.440 33.780 1190.560 ;
        RECT 107.100 1189.440 109.820 1190.560 ;
        RECT 3053.280 1189.440 3056.000 1190.560 ;
        RECT 3129.320 1189.440 3134.040 1190.560 ;
        RECT 35.060 1186.720 39.780 1187.840 ;
        RECT 78.300 1186.720 81.020 1187.840 ;
        RECT 3082.080 1186.720 3084.800 1187.840 ;
        RECT 3123.320 1186.720 3128.040 1187.840 ;
        RECT 41.060 1184.000 45.780 1185.120 ;
        RECT 83.100 1184.000 85.820 1185.120 ;
        RECT 3077.280 1184.000 3080.000 1185.120 ;
        RECT 3117.320 1184.000 3122.040 1185.120 ;
        RECT 47.060 1181.280 51.780 1182.400 ;
        RECT 87.900 1181.280 90.620 1182.400 ;
        RECT 3072.480 1181.280 3075.200 1182.400 ;
        RECT 3111.320 1181.280 3116.040 1182.400 ;
        RECT 53.060 1178.560 57.780 1179.680 ;
        RECT 92.700 1178.560 95.420 1179.680 ;
        RECT 3067.680 1178.560 3070.400 1179.680 ;
        RECT 3105.320 1178.560 3110.040 1179.680 ;
        RECT 59.060 1175.840 63.780 1176.960 ;
        RECT 97.500 1175.840 100.220 1176.960 ;
        RECT 3062.880 1175.840 3065.600 1176.960 ;
        RECT 3099.320 1175.840 3104.040 1176.960 ;
        RECT 65.060 1173.120 69.780 1174.240 ;
        RECT 102.300 1173.120 105.020 1174.240 ;
        RECT 3058.080 1173.120 3060.800 1174.240 ;
        RECT 3093.320 1173.120 3098.040 1174.240 ;
        RECT 23.060 1126.880 27.780 1128.000 ;
        RECT 111.900 1126.880 114.620 1128.000 ;
        RECT 3048.480 1126.880 3051.200 1128.000 ;
        RECT 3135.320 1126.880 3140.040 1128.000 ;
        RECT 29.060 1124.160 33.780 1125.280 ;
        RECT 107.100 1124.160 109.820 1125.280 ;
        RECT 3053.280 1124.160 3056.000 1125.280 ;
        RECT 3129.320 1124.160 3134.040 1125.280 ;
        RECT 35.060 1121.440 39.780 1122.560 ;
        RECT 78.300 1121.440 81.020 1122.560 ;
        RECT 3082.080 1121.440 3084.800 1122.560 ;
        RECT 3123.320 1121.440 3128.040 1122.560 ;
        RECT 41.060 1118.720 45.780 1119.840 ;
        RECT 83.100 1118.720 85.820 1119.840 ;
        RECT 3077.280 1118.720 3080.000 1119.840 ;
        RECT 3117.320 1118.720 3122.040 1119.840 ;
        RECT 47.060 1116.000 51.780 1117.120 ;
        RECT 87.900 1116.000 90.620 1117.120 ;
        RECT 3072.480 1116.000 3075.200 1117.120 ;
        RECT 3111.320 1116.000 3116.040 1117.120 ;
        RECT 53.060 1113.280 57.780 1114.400 ;
        RECT 92.700 1113.280 95.420 1114.400 ;
        RECT 3067.680 1113.280 3070.400 1114.400 ;
        RECT 3105.320 1113.280 3110.040 1114.400 ;
        RECT 59.060 1110.560 63.780 1111.680 ;
        RECT 97.500 1110.560 100.220 1111.680 ;
        RECT 3062.880 1110.560 3065.600 1111.680 ;
        RECT 3099.320 1110.560 3104.040 1111.680 ;
        RECT 65.060 1107.840 69.780 1108.960 ;
        RECT 102.300 1107.840 105.020 1108.960 ;
        RECT 3058.080 1107.840 3060.800 1108.960 ;
        RECT 3093.320 1107.840 3098.040 1108.960 ;
        RECT 3048.480 1061.600 3051.200 1062.720 ;
        RECT 3135.320 1061.600 3140.040 1062.720 ;
        RECT 3053.280 1058.880 3056.000 1060.000 ;
        RECT 3129.320 1058.880 3134.040 1060.000 ;
        RECT 23.060 1056.160 27.780 1057.280 ;
        RECT 111.900 1056.160 114.620 1057.280 ;
        RECT 3082.080 1056.160 3084.800 1057.280 ;
        RECT 3123.320 1056.160 3128.040 1057.280 ;
        RECT 29.060 1053.440 33.780 1054.560 ;
        RECT 107.100 1053.440 109.820 1054.560 ;
        RECT 3077.280 1053.440 3080.000 1054.560 ;
        RECT 3117.320 1053.440 3122.040 1054.560 ;
        RECT 35.060 1050.720 39.780 1051.840 ;
        RECT 78.300 1050.720 81.020 1051.840 ;
        RECT 3072.480 1050.720 3075.200 1051.840 ;
        RECT 3111.320 1050.720 3116.040 1051.840 ;
        RECT 41.060 1048.000 45.780 1049.120 ;
        RECT 83.100 1048.000 85.820 1049.120 ;
        RECT 3067.680 1048.000 3070.400 1049.120 ;
        RECT 3105.320 1048.000 3110.040 1049.120 ;
        RECT 47.060 1045.280 51.780 1046.400 ;
        RECT 87.900 1045.280 90.620 1046.400 ;
        RECT 3062.880 1045.280 3065.600 1046.400 ;
        RECT 3099.320 1045.280 3104.040 1046.400 ;
        RECT 53.060 1042.560 57.780 1043.680 ;
        RECT 92.700 1042.560 95.420 1043.680 ;
        RECT 3058.080 1042.560 3060.800 1043.680 ;
        RECT 3093.320 1042.560 3098.040 1043.680 ;
        RECT 59.060 1039.840 63.780 1040.960 ;
        RECT 97.500 1039.840 100.220 1040.960 ;
        RECT 65.060 1037.120 69.780 1038.240 ;
        RECT 102.300 1037.120 105.020 1038.240 ;
        RECT 1047.520 138.410 1064.310 140.415 ;
        RECT 1040.955 135.520 1045.275 136.640 ;
        RECT 1118.020 135.235 1128.720 136.880 ;
        RECT 1135.355 133.320 1138.075 134.440 ;
        RECT 654.975 38.040 659.295 39.160 ;
        RECT 698.860 37.945 699.580 38.665 ;
        RECT 661.735 34.720 666.055 35.840 ;
        RECT 692.360 35.125 693.080 35.845 ;
        RECT 687.000 22.485 688.955 32.480 ;
        RECT 694.000 10.880 696.410 32.480 ;
      LAYER via4 ;
        RECT 687.380 30.890 688.560 32.070 ;
        RECT 687.380 29.290 688.560 30.470 ;
        RECT 687.380 27.690 688.560 28.870 ;
        RECT 687.380 26.090 688.560 27.270 ;
        RECT 687.380 24.490 688.560 25.670 ;
        RECT 687.380 22.890 688.560 24.070 ;
        RECT 694.660 19.290 695.840 20.470 ;
        RECT 694.660 17.690 695.840 18.870 ;
        RECT 694.660 16.090 695.840 17.270 ;
        RECT 694.660 14.490 695.840 15.670 ;
        RECT 694.660 12.890 695.840 14.070 ;
        RECT 694.660 11.290 695.840 12.470 ;
      LAYER met5 ;
        RECT 687.380 30.890 688.560 32.070 ;
        RECT 687.380 29.290 688.560 30.470 ;
        RECT 687.380 27.690 688.560 28.870 ;
        RECT 687.380 26.090 688.560 27.270 ;
        RECT 687.380 24.490 688.560 25.670 ;
        RECT 687.380 22.890 688.560 24.070 ;
        RECT 694.660 19.290 695.840 20.470 ;
        RECT 694.660 17.690 695.840 18.870 ;
        RECT 694.660 16.090 695.840 17.270 ;
        RECT 694.660 14.490 695.840 15.670 ;
        RECT 694.660 12.890 695.840 14.070 ;
        RECT 694.660 11.290 695.840 12.470 ;
  END
END manual_power_connections
END LIBRARY

