* NGSPICE file created from caravel_clocking.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__274__B1 _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_432_ _351_/Y _432_/D _343_/S VGND VGND VPWR VPWR _432_/Q sky130_fd_sc_hd__dfrtp_4
X_294_ _450_/Q VGND VGND VPWR VPWR _296_/A sky130_fd_sc_hd__inv_2
X_363_ _445_/Q _444_/Q VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__xnor2_1
X_346_ _346_/A VGND VGND VPWR VPWR _410_/S sky130_fd_sc_hd__clkinv_4
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_415_ _411_/A1 _415_/D VGND VGND VPWR VPWR _415_/Q sky130_fd_sc_hd__dfxtp_1
X_277_ _282_/A VGND VGND VPWR VPWR _332_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _411_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ _329_/A _329_/B VGND VGND VPWR VPWR _442_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__443__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_258__3 _464_/CLK VGND VGND VPWR VPWR _457_/CLK sky130_fd_sc_hd__inv_4
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ _448_/Q _326_/B _397_/X VGND VGND VPWR VPWR _293_/Y sky130_fd_sc_hd__nand3b_1
X_362_ _444_/Q VGND VGND VPWR VPWR _362_/Y sky130_fd_sc_hd__clkinv_2
X_431_ _351_/Y _431_/D _343_/S VGND VGND VPWR VPWR _431_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_276_ _443_/Q VGND VGND VPWR VPWR _282_/A sky130_fd_sc_hd__inv_2
X_345_ _345_/A VGND VGND VPWR VPWR _404_/S sky130_fd_sc_hd__clkinv_4
X_414_ _411_/A1 _430_/Q VGND VGND VPWR VPWR _414_/Q sky130_fd_sc_hd__dfxtp_1
X_259_ _263_/A _409_/X VGND VGND VPWR VPWR _261_/A sky130_fd_sc_hd__nand2_1
X_328_ _332_/A _332_/B _442_/Q VGND VGND VPWR VPWR _329_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__310__B1 _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 _393_/X VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_1
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _443_/Q _290_/Y _291_/Y VGND VGND VPWR VPWR _292_/Y sky130_fd_sc_hd__o21bai_1
X_430_ _351_/Y _430_/D _343_/S VGND VGND VPWR VPWR _430_/Q sky130_fd_sc_hd__dfrtp_4
X_361_ _453_/Q _361_/B VGND VGND VPWR VPWR _361_/X sky130_fd_sc_hd__xor2_1
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_344_ _344_/A VGND VGND VPWR VPWR _420_/D sky130_fd_sc_hd__buf_1
X_413_ _455_/Q _413_/A1 _413_/S VGND VGND VPWR VPWR _413_/X sky130_fd_sc_hd__mux2_1
X_275_ _345_/A _275_/B _275_/C VGND VGND VPWR VPWR _281_/A sky130_fd_sc_hd__nand3b_1
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_327_ _335_/A _407_/X VGND VGND VPWR VPWR _329_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__386__A1 _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__439__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput11 _375_/Y VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_2
XANTENNA__422__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ _299_/B VGND VGND VPWR VPWR _291_/Y sky130_fd_sc_hd__inv_2
X_360_ _452_/Q _451_/Q VGND VGND VPWR VPWR _361_/B sky130_fd_sc_hd__nor2_1
X_412_ _412_/A0 _426_/Q _425_/D VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__mux2_1
X_343_ hold1/A _343_/A1 _343_/S VGND VGND VPWR VPWR _344_/A sky130_fd_sc_hd__mux2_2
X_274_ _432_/Q _431_/Q _430_/Q VGND VGND VPWR VPWR _275_/C sky130_fd_sc_hd__o21a_1
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_257_ _257_/A _257_/B VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__nand2_1
X_326_ _332_/A _326_/B VGND VGND VPWR VPWR _335_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_342__7 _393_/X VGND VGND VPWR VPWR _421_/CLK sky130_fd_sc_hd__inv_4
X_309_ _450_/Q _449_/Q VGND VGND VPWR VPWR _309_/Y sky130_fd_sc_hd__nor2_1
Xoutput12 _394_/X VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_1
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A sel[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_290_ _449_/Q _448_/Q VGND VGND VPWR VPWR _290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clkbuf_0_pll_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_273_ _454_/Q VGND VGND VPWR VPWR _275_/B sky130_fd_sc_hd__inv_2
XANTENNA__404__A1 _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_411_ _439_/Q _411_/A1 _411_/S VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__mux2_1
XANTENNA__446__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_256_ _260_/A _260_/B _458_/Q VGND VGND VPWR VPWR _257_/B sky130_fd_sc_hd__nand3_1
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ _321_/Y _324_/Y _283_/Y VGND VGND VPWR VPWR _443_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__468__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ _308_/A _440_/Q VGND VGND VPWR VPWR _308_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_410_ _438_/Q _373_/Y _410_/S VGND VGND VPWR VPWR _410_/X sky130_fd_sc_hd__mux2_1
X_272_ _272_/A _451_/Q VGND VGND VPWR VPWR _345_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_255_ _263_/A _396_/X VGND VGND VPWR VPWR _257_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_324_ _322_/Y _323_/X _275_/C VGND VGND VPWR VPWR _324_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__428__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_238_ _233_/Y _234_/Y _237_/Y _462_/Q VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__a22o_1
X_307_ _442_/Q _441_/Q VGND VGND VPWR VPWR _308_/A sky130_fd_sc_hd__nor2_1
XANTENNA__430__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_271_ _453_/Q _452_/Q VGND VGND VPWR VPWR _272_/A sky130_fd_sc_hd__nor2_1
X_469_ _413_/A1 _469_/D _343_/S VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfrtp_1
X_254_ _260_/A _254_/B VGND VGND VPWR VPWR _263_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_323_ _432_/Q _416_/Q VGND VGND VPWR VPWR _323_/X sky130_fd_sc_hd__and2_1
XANTENNA__434__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_237_ _467_/Q _235_/Y _236_/Y VGND VGND VPWR VPWR _237_/Y sky130_fd_sc_hd__o21bai_1
X_306_ _306_/A _306_/B _406_/S VGND VGND VPWR VPWR _312_/A sky130_fd_sc_hd__nand3_1
XANTENNA__470__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input6_A sel2[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ _270_/A _270_/B VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__nand2_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_468_ _413_/A1 _468_/D _343_/S VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__424__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_399_ _398_/X _432_/Q _443_/Q VGND VGND VPWR VPWR _399_/X sky130_fd_sc_hd__mux2_1
XANTENNA__457__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ _432_/Q _416_/Q VGND VGND VPWR VPWR _322_/Y sky130_fd_sc_hd__nor2_1
X_253_ _253_/A _253_/B _260_/B VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__nand3_1
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_236_ _390_/X VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__inv_2
X_305_ _442_/Q _441_/Q _440_/Q VGND VGND VPWR VPWR _406_/S sky130_fd_sc_hd__nor3b_4
Xclkbuf_1_1_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _413_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__317__S _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_219_ _465_/Q _464_/Q VGND VGND VPWR VPWR _220_/A sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_467_ _413_/A1 _467_/D _343_/S VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfrtp_4
X_398_ _361_/X _432_/Q _404_/S VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__mux2_1
X_252_ _250_/Y _260_/A _248_/B VGND VGND VPWR VPWR _253_/B sky130_fd_sc_hd__o21bai_1
X_321_ _321_/A _321_/B _414_/Q VGND VGND VPWR VPWR _321_/Y sky130_fd_sc_hd__nand3_1
Xclkbuf_1_0_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _464_/CLK sky130_fd_sc_hd__clkbuf_2
X_235_ _461_/Q _460_/Q VGND VGND VPWR VPWR _235_/Y sky130_fd_sc_hd__nor2_1
X_304_ _447_/Q VGND VGND VPWR VPWR _306_/B sky130_fd_sc_hd__inv_2
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ _210_/Y _214_/Y _217_/Y VGND VGND VPWR VPWR _467_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_1_1_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _412_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _453_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_466_ _413_/A1 _466_/D _343_/S VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfstp_1
X_397_ _283_/Y _443_/Q _397_/S VGND VGND VPWR VPWR _397_/X sky130_fd_sc_hd__mux2_4
XANTENNA__423__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__433__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_251_ _437_/Q _438_/Q _436_/Q _234_/Y VGND VGND VPWR VPWR _260_/A sky130_fd_sc_hd__o211ai_4
X_320_ _415_/Q _431_/Q VGND VGND VPWR VPWR _321_/B sky130_fd_sc_hd__or2b_1
X_449_ _449_/CLK _449_/D _343_/S VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfstp_1
X_234_ _462_/Q _461_/Q VGND VGND VPWR VPWR _234_/Y sky130_fd_sc_hd__nor2_2
X_303_ _303_/A _303_/B VGND VGND VPWR VPWR _397_/S sky130_fd_sc_hd__nor2_1
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_217_ _224_/A _254_/B VGND VGND VPWR VPWR _217_/Y sky130_fd_sc_hd__nand2_2
X_302__5 _411_/A1 VGND VGND VPWR VPWR _447_/CLK sky130_fd_sc_hd__inv_4
XANTENNA__458__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_396_ _395_/X _438_/Q _467_/Q VGND VGND VPWR VPWR _396_/X sky130_fd_sc_hd__mux2_1
X_465_ _413_/A1 _465_/D _343_/S VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfrtp_1
X_250_ _250_/A _456_/Q VGND VGND VPWR VPWR _250_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_input4_A sel2[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_379_ _368_/Y _436_/Q _391_/S VGND VGND VPWR VPWR _379_/X sky130_fd_sc_hd__mux2_1
X_448_ _453_/CLK _448_/D _343_/S VGND VGND VPWR VPWR _448_/Q sky130_fd_sc_hd__dfrtn_1
X_233_ _467_/Q _460_/Q _390_/X VGND VGND VPWR VPWR _233_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_216_ _467_/Q VGND VGND VPWR VPWR _254_/B sky130_fd_sc_hd__clkinv_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__427__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_464_ _464_/CLK _464_/D _343_/S VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfstp_1
X_395_ _367_/X _438_/Q _408_/S VGND VGND VPWR VPWR _395_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__452__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__442__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_447_ _447_/CLK _447_/D _343_/S VGND VGND VPWR VPWR _447_/Q sky130_fd_sc_hd__dfstp_1
X_232_ _380_/X _217_/Y _231_/Y VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__a21bo_1
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_301_ _291_/Y _448_/Q _293_/Y VGND VGND VPWR VPWR _448_/D sky130_fd_sc_hd__a21bo_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_215_ _437_/Q _438_/Q _436_/Q VGND VGND VPWR VPWR _224_/A sky130_fd_sc_hd__o21ai_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__467__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_394_ _412_/X _354_/Y _425_/Q VGND VGND VPWR VPWR _394_/X sky130_fd_sc_hd__mux2_1
X_463_ _464_/CLK _463_/D _343_/S VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_377_ _470_/Q _377_/B VGND VGND VPWR VPWR _470_/D sky130_fd_sc_hd__xor2_1
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_446_ _453_/CLK _446_/D _343_/S VGND VGND VPWR VPWR _446_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clkbuf_0_ext_clk/X sky130_fd_sc_hd__clkbuf_16
X_231_ _231_/A _254_/B _463_/Q VGND VGND VPWR VPWR _231_/Y sky130_fd_sc_hd__nand3_1
X_300_ _296_/B _299_/X _292_/Y VGND VGND VPWR VPWR _449_/D sky130_fd_sc_hd__o21ai_1
X_429_ _351_/Y _429_/D _343_/S VGND VGND VPWR VPWR _432_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 ext_clk_sel VGND VGND VPWR VPWR _374_/A sky130_fd_sc_hd__clkbuf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_214_ _211_/Y _212_/X _222_/C VGND VGND VPWR VPWR _214_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__313__A _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__436__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_393_ _412_/X _351_/Y _425_/Q VGND VGND VPWR VPWR _393_/X sky130_fd_sc_hd__mux2_1
X_462_ _464_/CLK _462_/D _343_/S VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__451__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_376_ _469_/Q _436_/Q _468_/Q VGND VGND VPWR VPWR _377_/B sky130_fd_sc_hd__nor3_1
X_445_ _453_/CLK _445_/D _343_/S VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_input2_A ext_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_230_ _392_/X _217_/Y _229_/Y VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__a21bo_1
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__385__A1 _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_428_ _351_/Y _428_/D _343_/S VGND VGND VPWR VPWR _431_/D sky130_fd_sc_hd__dfstp_1
X_359_ _452_/Q _451_/Q VGND VGND VPWR VPWR _359_/Y sky130_fd_sc_hd__xnor2_1
Xinput2 ext_reset VGND VGND VPWR VPWR _375_/A sky130_fd_sc_hd__clkbuf_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ _437_/Q _438_/Q _436_/Q VGND VGND VPWR VPWR _222_/C sky130_fd_sc_hd__o21a_1
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__441__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_392_ _391_/X _437_/Q _467_/Q VGND VGND VPWR VPWR _392_/X sky130_fd_sc_hd__mux2_1
X_461_ _461_/CLK _461_/D _343_/S VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_375_ _375_/A _421_/Q VGND VGND VPWR VPWR _375_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_444_ _453_/CLK _444_/D _343_/S VGND VGND VPWR VPWR _444_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_427_ _351_/Y _427_/D _343_/S VGND VGND VPWR VPWR _430_/D sky130_fd_sc_hd__dfrtp_1
X_358_ _451_/Q VGND VGND VPWR VPWR _358_/Y sky130_fd_sc_hd__clkinv_2
Xinput3 resetb VGND VGND VPWR VPWR _343_/S sky130_fd_sc_hd__buf_12
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ _405_/X _283_/Y _288_/Y VGND VGND VPWR VPWR _451_/D sky130_fd_sc_hd__a21bo_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_212_ _419_/Q _438_/Q VGND VGND VPWR VPWR _212_/X sky130_fd_sc_hd__and2_1
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__464__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__445__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_391_ _369_/Y _437_/Q _391_/S VGND VGND VPWR VPWR _391_/X sky130_fd_sc_hd__mux2_1
X_460_ _464_/CLK _460_/D _343_/S VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__460__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_374_ _374_/A VGND VGND VPWR VPWR _424_/D sky130_fd_sc_hd__clkinv_4
X_443_ _411_/A1 _443_/D _343_/S VGND VGND VPWR VPWR _443_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_426_ _411_/A1 hold1/X _343_/S VGND VGND VPWR VPWR _426_/Q sky130_fd_sc_hd__dfrtp_1
Xinput4 sel2[0] VGND VGND VPWR VPWR _433_/D sky130_fd_sc_hd__clkbuf_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _442_/Q _357_/B VGND VGND VPWR VPWR _357_/X sky130_fd_sc_hd__xor2_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _288_/A _451_/Q _326_/B VGND VGND VPWR VPWR _288_/Y sky130_fd_sc_hd__nand3_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _419_/Q _438_/Q VGND VGND VPWR VPWR _211_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_409_ _408_/X _437_/Q _467_/Q VGND VGND VPWR VPWR _409_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_390_ _217_/Y _467_/Q _390_/S VGND VGND VPWR VPWR _390_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_373_ _469_/Q _468_/Q VGND VGND VPWR VPWR _373_/Y sky130_fd_sc_hd__xnor2_1
X_442_ _411_/A1 _442_/D _343_/S VGND VGND VPWR VPWR _442_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__447__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_425_ _411_/A1 _425_/D _343_/S VGND VGND VPWR VPWR _425_/Q sky130_fd_sc_hd__dfrtp_1
Xinput5 sel2[1] VGND VGND VPWR VPWR _434_/D sky130_fd_sc_hd__clkbuf_1
X_356_ _441_/Q _440_/Q VGND VGND VPWR VPWR _357_/B sky130_fd_sc_hd__nor2_1
X_287_ _402_/X _283_/Y _286_/Y VGND VGND VPWR VPWR _452_/D sky130_fd_sc_hd__a21bo_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_210_ _210_/A _210_/B _417_/Q VGND VGND VPWR VPWR _210_/Y sky130_fd_sc_hd__nand3_1
X_408_ _365_/Y _437_/Q _408_/S VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__mux2_1
X_339_ _439_/Q _339_/B VGND VGND VPWR VPWR _439_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__414__D _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_340__9 _393_/X VGND VGND VPWR VPWR _423_/CLK sky130_fd_sc_hd__inv_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_372_ _468_/Q VGND VGND VPWR VPWR _372_/Y sky130_fd_sc_hd__clkinv_2
X_441_ _441_/CLK _441_/D _343_/S VGND VGND VPWR VPWR _441_/Q sky130_fd_sc_hd__dfstp_2
Xclkbuf_1_0_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _343_/A1 sky130_fd_sc_hd__clkbuf_2
X_424_ _411_/A1 _424_/D _343_/S VGND VGND VPWR VPWR _425_/D sky130_fd_sc_hd__dfrtp_1
X_355_ _441_/Q _440_/Q VGND VGND VPWR VPWR _355_/Y sky130_fd_sc_hd__xnor2_1
X_286_ _288_/A _452_/Q _326_/B VGND VGND VPWR VPWR _286_/Y sky130_fd_sc_hd__nand3_1
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 sel2[2] VGND VGND VPWR VPWR _435_/D sky130_fd_sc_hd__clkbuf_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ _346_/A _269_/B _269_/C VGND VGND VPWR VPWR _270_/B sky130_fd_sc_hd__nand3_1
X_407_ _406_/X _432_/Q _443_/Q VGND VGND VPWR VPWR _407_/X sky130_fd_sc_hd__mux2_1
X_338_ _430_/Q _364_/A _444_/Q VGND VGND VPWR VPWR _339_/B sky130_fd_sc_hd__nand3b_1
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ _465_/Q _371_/B VGND VGND VPWR VPWR _371_/X sky130_fd_sc_hd__xor2_1
X_440_ _411_/A1 _440_/D _343_/S VGND VGND VPWR VPWR _440_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_423_ _423_/CLK _423_/D _343_/S VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfstp_1
X_354_ _269_/B _413_/X _231_/A _353_/Y VGND VGND VPWR VPWR _354_/Y sky130_fd_sc_hd__o2bb2ai_2
X_285_ _399_/X _283_/Y _284_/Y VGND VGND VPWR VPWR _453_/D sky130_fd_sc_hd__a21bo_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__448__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 sel[0] VGND VGND VPWR VPWR _427_/D sky130_fd_sc_hd__clkbuf_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_268_ _346_/A _269_/B _269_/C VGND VGND VPWR VPWR _270_/A sky130_fd_sc_hd__a21o_1
X_406_ _357_/X _432_/Q _406_/S VGND VGND VPWR VPWR _406_/X sky130_fd_sc_hd__mux2_1
X_337_ _446_/Q _445_/Q VGND VGND VPWR VPWR _364_/A sky130_fd_sc_hd__nor2_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__463__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__315__S _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_370_ _464_/Q _463_/Q VGND VGND VPWR VPWR _371_/B sky130_fd_sc_hd__nor2_1
X_422_ _422_/CLK hold2/X _343_/S VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfstp_1
X_353_ _466_/Q _459_/Q VGND VGND VPWR VPWR _353_/Y sky130_fd_sc_hd__xnor2_1
X_284_ _288_/A _453_/Q _332_/B VGND VGND VPWR VPWR _284_/Y sky130_fd_sc_hd__nand3_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 sel[1] VGND VGND VPWR VPWR _428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_267_ _455_/Q VGND VGND VPWR VPWR _269_/C sky130_fd_sc_hd__inv_2
X_336_ _334_/Y _335_/A _335_/Y VGND VGND VPWR VPWR _440_/D sky130_fd_sc_hd__o21ai_1
X_405_ _404_/X _430_/Q _443_/Q VGND VGND VPWR VPWR _405_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_319_ _415_/D _415_/Q VGND VGND VPWR VPWR _321_/A sky130_fd_sc_hd__or2b_1
XANTENNA__432__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__459__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input9_A sel[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_421_ _421_/CLK hold3/X _343_/S VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__338__A_N _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_352_ _437_/Q _438_/Q VGND VGND VPWR VPWR _413_/S sky130_fd_sc_hd__nor2_1
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 sel[2] VGND VGND VPWR VPWR _429_/D sky130_fd_sc_hd__clkbuf_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _303_/A _326_/B VGND VGND VPWR VPWR _283_/Y sky130_fd_sc_hd__nand2_2
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_266_ _436_/Q VGND VGND VPWR VPWR _269_/B sky130_fd_sc_hd__clkinv_4
X_335_ _335_/A _386_/X VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__nand2_1
X_404_ _358_/Y _430_/Q _404_/S VGND VGND VPWR VPWR _404_/X sky130_fd_sc_hd__mux2_1
X_249_ _458_/Q _457_/Q VGND VGND VPWR VPWR _250_/A sky130_fd_sc_hd__nor2_1
X_318_ _318_/A VGND VGND VPWR VPWR _444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_378__13 VGND VGND VPWR VPWR _378__13/HI _423_/D sky130_fd_sc_hd__conb_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_420_ _453_/CLK _420_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_282_ _282_/A VGND VGND VPWR VPWR _326_/B sky130_fd_sc_hd__clkbuf_2
X_351_ _288_/A _349_/Y _350_/X VGND VGND VPWR VPWR _351_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__426__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_334_ _440_/Q VGND VGND VPWR VPWR _334_/Y sky130_fd_sc_hd__inv_2
X_403_ _432_/Q _363_/Y _403_/S VGND VGND VPWR VPWR _403_/X sky130_fd_sc_hd__mux2_1
X_265_ _469_/Q _470_/Q _468_/Q VGND VGND VPWR VPWR _346_/A sky130_fd_sc_hd__nor3b_2
X_248_ _390_/S _248_/B _408_/S VGND VGND VPWR VPWR _253_/A sky130_fd_sc_hd__nand3_1
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_317_ _400_/X _444_/Q _430_/Q VGND VGND VPWR VPWR _318_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ _430_/Q _411_/X VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__and2b_2
X_281_ _281_/A _332_/B _281_/C VGND VGND VPWR VPWR _454_/D sky130_fd_sc_hd__nand3_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_264_ _262_/Y _263_/A _263_/Y VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__o21ai_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_333_ _333_/A _333_/B VGND VGND VPWR VPWR _441_/D sky130_fd_sc_hd__nand2_1
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_402_ _401_/X _415_/D _443_/Q VGND VGND VPWR VPWR _402_/X sky130_fd_sc_hd__mux2_1
X_247_ _458_/Q _457_/Q _456_/Q VGND VGND VPWR VPWR _408_/S sky130_fd_sc_hd__nor3b_2
X_316_ _316_/A VGND VGND VPWR VPWR _445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__431__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ _288_/A _345_/A _275_/B VGND VGND VPWR VPWR _281_/C sky130_fd_sc_hd__o21bai_1
XANTENNA_input7_A sel[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__435__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _263_/A _384_/X VGND VGND VPWR VPWR _263_/Y sky130_fd_sc_hd__nand2_1
X_332_ _332_/A _332_/B _441_/Q VGND VGND VPWR VPWR _333_/B sky130_fd_sc_hd__nand3_1
X_401_ _359_/Y _415_/D _404_/S VGND VGND VPWR VPWR _401_/X sky130_fd_sc_hd__mux2_1
X_246_ _459_/Q VGND VGND VPWR VPWR _248_/B sky130_fd_sc_hd__clkinv_4
X_315_ _403_/X _445_/Q _430_/Q VGND VGND VPWR VPWR _316_/A sky130_fd_sc_hd__mux2_1
XANTENNA__454__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_229_ _231_/A _254_/B _464_/Q VGND VGND VPWR VPWR _229_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__450__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ _456_/Q VGND VGND VPWR VPWR _262_/Y sky130_fd_sc_hd__inv_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _335_/A _382_/X VGND VGND VPWR VPWR _333_/A sky130_fd_sc_hd__nand2_1
X_400_ _415_/D _362_/Y _403_/S VGND VGND VPWR VPWR _400_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_245_ _437_/Q _438_/Q _436_/Q _234_/Y VGND VGND VPWR VPWR _390_/S sky130_fd_sc_hd__o211a_1
X_314_ _446_/Q _314_/B VGND VGND VPWR VPWR _446_/D sky130_fd_sc_hd__xor2_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330__6 _411_/A1 VGND VGND VPWR VPWR _441_/CLK sky130_fd_sc_hd__inv_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_228_ _389_/X _217_/Y _227_/Y VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__a21bo_1
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__429__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__437__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_261_ _261_/A _261_/B VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__nand2_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_459_ _459_/CLK _459_/D _343_/S VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_313_ _430_/Q _445_/Q _444_/Q VGND VGND VPWR VPWR _314_/B sky130_fd_sc_hd__nor3_1
X_227_ _231_/A _260_/B _465_/Q VGND VGND VPWR VPWR _227_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__469__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _260_/A _260_/B _457_/Q VGND VGND VPWR VPWR _261_/B sky130_fd_sc_hd__nand3_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A sel2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_458_ _464_/CLK _458_/D _343_/S VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfrtn_1
X_389_ _388_/X _438_/Q _467_/Q VGND VGND VPWR VPWR _389_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_243_ _236_/Y _460_/Q _233_/Y VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__a21o_1
X_312_ _312_/A _312_/B _332_/B VGND VGND VPWR VPWR _447_/D sky130_fd_sc_hd__nand3_1
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_226_ _226_/A _260_/B _226_/C VGND VGND VPWR VPWR _466_/D sky130_fd_sc_hd__nand3_1
XFILLER_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_209_ _437_/Q _418_/Q VGND VGND VPWR VPWR _210_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__438__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__466__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__453__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__278__B1 _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_457_ _457_/CLK _457_/D _343_/S VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfstp_1
X_388_ _371_/X _438_/Q _391_/S VGND VGND VPWR VPWR _388_/X sky130_fd_sc_hd__mux2_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_242_ _240_/Y _241_/X _237_/Y VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__o21ai_1
X_311_ _308_/Y _332_/A _306_/B VGND VGND VPWR VPWR _312_/B sky130_fd_sc_hd__o21bai_1
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_225_ _231_/A _347_/A _222_/B VGND VGND VPWR VPWR _226_/C sky130_fd_sc_hd__o21bai_1
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_341__8 _393_/X VGND VGND VPWR VPWR _422_/CLK sky130_fd_sc_hd__inv_4
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ _418_/Q _437_/Q VGND VGND VPWR VPWR _210_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_456_ _464_/CLK _456_/D _343_/S VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfrtn_1
X_387_ _437_/Q _372_/Y _410_/S VGND VGND VPWR VPWR _387_/X sky130_fd_sc_hd__mux2_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_310_ _432_/Q _431_/Q _430_/Q _309_/Y VGND VGND VPWR VPWR _332_/A sky130_fd_sc_hd__o211ai_2
X_241_ _460_/Q _390_/X VGND VGND VPWR VPWR _241_/X sky130_fd_sc_hd__and2b_1
X_439_ _453_/CLK _439_/D _343_/S VGND VGND VPWR VPWR _439_/Q sky130_fd_sc_hd__dfstp_1
X_224_ _224_/A VGND VGND VPWR VPWR _231_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__405__A1 _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_207_ _207_/A VGND VGND VPWR VPWR _468_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__449__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_298__4 _453_/CLK VGND VGND VPWR VPWR _449_/CLK sky130_fd_sc_hd__inv_4
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_455_ _413_/A1 _455_/D _343_/S VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__462__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_386_ _385_/X _430_/Q _443_/Q VGND VGND VPWR VPWR _386_/X sky130_fd_sc_hd__mux2_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_240_ _461_/Q VGND VGND VPWR VPWR _240_/Y sky130_fd_sc_hd__inv_2
X_438_ _354_/Y _438_/D _343_/S VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfrtp_4
X_369_ _464_/Q _463_/Q VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__xnor2_1
X_223_ _254_/B VGND VGND VPWR VPWR _260_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_206_ _387_/X _468_/Q _436_/Q VGND VGND VPWR VPWR _207_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__455__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_385_ _334_/Y _430_/Q _406_/S VGND VGND VPWR VPWR _385_/X sky130_fd_sc_hd__mux2_1
X_454_ _411_/A1 _454_/D _343_/S VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfstp_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ _354_/Y _437_/D _343_/S VGND VGND VPWR VPWR _437_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_368_ _463_/Q VGND VGND VPWR VPWR _368_/Y sky130_fd_sc_hd__clkinv_2
X_299_ _448_/Q _299_/B VGND VGND VPWR VPWR _299_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_222_ _347_/A _222_/B _222_/C VGND VGND VPWR VPWR _226_/A sky130_fd_sc_hd__nand3b_1
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _205_/A VGND VGND VPWR VPWR _469_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clkbuf_0_pll_clk90/X sky130_fd_sc_hd__clkbuf_16
XFILLER_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__456__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__461__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_470_ _413_/A1 _470_/D _343_/S VGND VGND VPWR VPWR _470_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _383_/X _436_/Q _467_/Q VGND VGND VPWR VPWR _384_/X sky130_fd_sc_hd__mux2_1
X_453_ _453_/CLK _453_/D _343_/S VGND VGND VPWR VPWR _453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_367_ _458_/Q _367_/B VGND VGND VPWR VPWR _367_/X sky130_fd_sc_hd__xor2_1
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_436_ _354_/Y _436_/D _343_/S VGND VGND VPWR VPWR _436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_221_ _466_/Q VGND VGND VPWR VPWR _222_/B sky130_fd_sc_hd__inv_2
X_419_ _464_/CLK _438_/Q VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfxtp_1
X_204_ _410_/X _469_/Q _436_/Q VGND VGND VPWR VPWR _205_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__421__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__425__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit4 _431_/Q VGND VGND VPWR VPWR _415_/D sky130_fd_sc_hd__clkbuf_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_383_ _262_/Y _436_/Q _408_/S VGND VGND VPWR VPWR _383_/X sky130_fd_sc_hd__mux2_1
X_452_ _453_/CLK _452_/D _343_/S VGND VGND VPWR VPWR _452_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__440__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_366_ _457_/Q _456_/Q VGND VGND VPWR VPWR _367_/B sky130_fd_sc_hd__nor2_1
X_435_ _354_/Y _435_/D _343_/S VGND VGND VPWR VPWR _438_/D sky130_fd_sc_hd__dfrtp_1
X_297_ _450_/Q _292_/Y _293_/Y _303_/B VGND VGND VPWR VPWR _450_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_220_ _220_/A _463_/Q VGND VGND VPWR VPWR _347_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input1_A ext_clk_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_418_ _464_/CLK _437_/Q VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfxtp_1
X_239__1 _464_/CLK VGND VGND VPWR VPWR _461_/CLK sky130_fd_sc_hd__inv_4
X_349_ _454_/Q _447_/Q VGND VGND VPWR VPWR _349_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__444__SET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__465__RESET_B _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__343__S _343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_382_ _381_/X _431_/Q _443_/Q VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__mux2_1
X_451_ _453_/CLK _451_/D _343_/S VGND VGND VPWR VPWR _451_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _457_/Q _456_/Q VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__xnor2_1
X_434_ _354_/Y _434_/D _343_/S VGND VGND VPWR VPWR _437_/D sky130_fd_sc_hd__dfstp_1
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_296_ _296_/A _296_/B VGND VGND VPWR VPWR _303_/B sky130_fd_sc_hd__nand2_1
X_244__2 _464_/CLK VGND VGND VPWR VPWR _459_/CLK sky130_fd_sc_hd__inv_4
Xrebuffer5 _397_/S VGND VGND VPWR VPWR _306_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_417_ _413_/A1 _436_/Q VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfxtp_1
X_279_ _303_/A VGND VGND VPWR VPWR _288_/A sky130_fd_sc_hd__clkbuf_2
X_348_ _432_/Q _415_/D VGND VGND VPWR VPWR _411_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ _355_/Y _431_/Q _406_/S VGND VGND VPWR VPWR _381_/X sky130_fd_sc_hd__mux2_1
X_450_ _453_/CLK _450_/D _343_/S VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__350__A_N _430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _354_/Y _433_/D _343_/S VGND VGND VPWR VPWR _436_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_295_ _449_/Q VGND VGND VPWR VPWR _296_/B sky130_fd_sc_hd__clkinv_4
Xrebuffer6 _397_/X VGND VGND VPWR VPWR _299_/B sky130_fd_sc_hd__buf_2
X_364_ _364_/A _444_/Q VGND VGND VPWR VPWR _403_/S sky130_fd_sc_hd__nand2_1
X_347_ _347_/A VGND VGND VPWR VPWR _391_/S sky130_fd_sc_hd__clkinv_4
X_278_ _432_/Q _431_/Q _430_/Q VGND VGND VPWR VPWR _303_/A sky130_fd_sc_hd__o21ai_2
X_416_ _411_/A1 _432_/Q VGND VGND VPWR VPWR _416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_380_ _379_/X _436_/Q _467_/Q VGND VGND VPWR VPWR _380_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

